// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Wed Jul 29 15:53:56 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, 
        INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(46[12:14])
    
    wire reset;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(49[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, GHB, GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(95[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(96[21:25])
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(131[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(132[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(141[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(238[21:45])
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(240[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(241[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(242[22:30])
    
    wire n66949;
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(243[22:24])
    
    wire n50102;
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(244[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(246[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(247[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(248[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(249[22:30])
    wire [15:0]current;   // verilog/TinyFPGA_B.v(250[22:29])
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(251[22:35])
    wire [31:0]baudrate;   // verilog/TinyFPGA_B.v(253[15:23])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(282[22:33])
    
    wire data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(351[11:24])
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(359[15:20])
    
    wire pwm_setpoint_23__N_207, n12184, n12188, n6, n260, n12224, 
        n294, n298, n299, n300, n301, n302, n303, n304, n305, 
        n306, n307, n308, n309, n50101, n15, n4928, n4927, n4926, 
        n4925, n4924, n4923, n4922, n4921, n4920, n4919, n4918, 
        n4917, n4916, n50100, n61622;
    wire [23:0]pwm_setpoint_23__N_3;
    
    wire n50099;
    wire [7:0]commutation_state_7__N_208;
    
    wire commutation_state_7__N_216;
    wire [7:0]commutation_state_7__N_27;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(237[11:28])
    
    wire n36759, GHA_N_355, GLA_N_372, GHB_N_377, GLB_N_386, GHC_N_391, 
        GLC_N_400, dti_N_404, n29969, n29968, RX_N_2, n1744, n1742;
    wire [31:0]motor_state_23__N_91;
    
    wire n68073;
    wire [32:0]encoder0_position_scaled_23__N_43;
    wire [23:0]displacement_23__N_67;
    
    wire n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, 
        n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
        n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, 
        n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
        read_N_409, n67937, n50098, n1319, n36723, n61616, n49171, 
        n7, n6_adj_5659, n5, n4, n26, n67257, n19, n17, n16, 
        n15_adj_5660, n13, n11, n9, n8, n7_adj_5661, n6_adj_5662, 
        n5_adj_5663, n4_adj_5664, n1784, n1786, n1788, n1790, n1792, 
        n1794, n1796;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(239[11:28])
    
    wire n1822, n1824;
    wire [10:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [1:0]state;   // verilog/neopixel.v(16[11:16])
    wire [4:0]bit_ctr;   // verilog/neopixel.v(17[11:18])
    wire [10:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(27[14:16])
    
    wire n49724, n4915, n4914, n4913, n4912, n50097, n4911, n4910, 
        n49723, n49170, n625, n61610, n4940, n4937, n50096, n50095, 
        n29959, n50094, n36694, n69384, n50093, n49722, n50092, 
        n49721, n29956, n29953, n50091, n50090, n623;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n10, n9_adj_5665, n25, n24, n8_adj_5666, n23, n22, n21, 
        n20, n49720, n19_adj_5667, n17_adj_5668, n16_adj_5669, n50089, 
        n50088, n50087, n50086, n49719, n622, n621, n2, n14, 
        n15_adj_5670, n16_adj_5671, n17_adj_5672, n18, n19_adj_5673, 
        n20_adj_5674, n21_adj_5675, n22_adj_5676, n23_adj_5677, n24_adj_5678, 
        n25_adj_5679, n5774, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(94[13:20])
    
    wire n61606, n50085, n49169;
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[3] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[1] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(100[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(105[12:33])
    
    wire tx_active, n49718, n49495;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(115[11:16])
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire \FRAME_MATCHER.rx_data_ready_prev , n49168, n3470, n49167, 
        n2820, n49494, n50084, n50083, n29949, n49717, n50082, 
        n25398, n50081, n49166, n2873, n161, n68097, n49716, n50080, 
        n50079, n50078, n49715, n68099, n49154, n50077, n68101, 
        n67762, n61600, n50076, n49493, n50075, n50074, n50073, 
        n49165, n50072, n4909, n61598, n49714, n4908, n4907, n50071, 
        n50070, n50069, n50068, n61596, n50067, n50066, n50065, 
        n56912, n56911, n56910, n56909, n56908, n56907, n56906, 
        n56774, n56905, n56904, n56903, n56902, n56901, n56900, 
        n56899, n56898, n56897, n56896, n56895, n56894, n56893, 
        n56892, n56891, n56890, n56889, n56888, n56887, n56886, 
        n56885, n56884, n56883, n56882, n56881, n56880, n56879, 
        n56878, n56877, n56876, n56875, n29046, n56874, n56873, 
        n56872, n56871, n56870, n56869, n56868, n56867, n56866, 
        n56865, n56864, n56863, n56862, n56861, n56860, n29030, 
        n56859, n56858, n56857, n56856, n56855, n56854, n56853, 
        n56852, n56851, n56850, n56776, n56778, n56779, n56780, 
        n56781, n56782, n56784, n56785, n56786, n56787, n56788, 
        n56789, n56790, n56791, n56792, n56793, n56775, n56794, 
        n56795, n56796, n56797, n56798, n56799, n56800, n56801, 
        n56802, n56803, n56804, n56805, n56806, n28989, n56807, 
        n28987, n56808, n56809, n56810, n56811, n56812, n28981, 
        n56813, n56814, n56815, n56816, n56817, n56818, n56819, 
        n56820, n56821, n56822, n56823, n56824, n56825, n56826, 
        n56827, n56828, n56829, n56830, n56831, n56832, n56833, 
        n56834, n56835, n56836, n56837, n56838, n56839, n56840, 
        n56773, n56783, n56841, n56842, n56843, n56844, n56845, 
        n56847, n56848, n56849, n15_adj_5680, n49492, n49491, n50064, 
        n50063, n29946, n50062, n49713, n67728, n50061, n49490, 
        n50060, n50059, n50058, n49489, n49712, n50057, n49711, 
        n50056, n50055, n49488, n68808, n50054, n50621, n49487, 
        n49710, n50053, n50620, n50619, n50052, n49709, n50618, 
        n50617, n50616, n50051, n50050, n49153, n50615, n50614, 
        n50613, n50612, n50611, n50610, n50049, n50048, n50047, 
        n50609, n50608, n50607, n50046, n50045, n50606, n50605, 
        n61582, n50604, n50044, n50603, n50043, n50602, n50601, 
        n50600, n50599, n50598, n50597, n50596, n50595, n50594, 
        n50042, n50593, n50041, n50592, n50591, n50040, n50039, 
        n50038, n50037, n50036, n50035, n50034, n50033, n50032, 
        n50031, n50030, n50029, n50028, n50027, n50026, n50025, 
        n50024, n50023, n50022, n50021, n50020, n50019, n50018, 
        n50017, n50016, n50015, n50014, n61574, n50013, n50012, 
        n50011, n50010, n50009, n50008, n50007, n50006, n50005, 
        n50004, n50003, n61854, n50002, n50001, n50000, n49999, 
        n49998, n49474, n49997, n49996, n49681, n49995, n49994, 
        n49993, n49680, n49992, n49679, n49991, n49678, n49473, 
        n49990, n49989, n49472, n49988, n49987, n49986, n49677, 
        n49164, n49471, n49676, n49675, n49985, n49984, n49983, 
        n49674, n49673, n49672, n49982, n49671, n49981, n49980, 
        n42774, n42699, n49979, n49978, n61568, n49670, n49152, 
        n49669, n49668, n49977, n49470, n42804, n49976, n49975, 
        n42746, n42723, n68551, n25516, n61558, n25864, n59282, 
        n49974, n69378, n69372, n49973, n15_adj_5681, n11_adj_5682, 
        n49667, n10_adj_5683, n66068, n61552, n49469, n25810, n66995, 
        n61548, n4_adj_5684, n59675, n58659, n61540, n61538, n58000, 
        n12222, n59710, n32, n31, n49972, n49971, n49468, n67571, 
        n13_adj_5685, n67245, n67570, n14_adj_5686, n13_adj_5687, 
        n61524, Kp_23__N_1301, n61518, n61514, n61502, n61498, n25952, 
        n57948, n57935, n61492, n61488, n57921, n30, n29, n28, 
        n12186, n27, n26_adj_5688, n25_adj_5689, n24_adj_5690, n23_adj_5691, 
        n22_adj_5692, n21_adj_5693, n20_adj_5694, n19_adj_5695, n18_adj_5696, 
        n49467, n17_adj_5697, n16_adj_5698, n15_adj_5699, n14_adj_5700, 
        n13_adj_5701, n12, n11_adj_5702, n10_adj_5703, n9_adj_5704, 
        n8_adj_5705, n7_adj_5706, n6_adj_5707, \FRAME_MATCHER.i_31__N_2509 , 
        \FRAME_MATCHER.i_31__N_2513 , Kp_23__N_1748, n61478, n57917, 
        n5_adj_5708, n49970, n43474, n43530, n43462, n43349, n29889, 
        n29885, n29884, n29881, n29878, n29874, n29870, n29867, 
        n29866, n59879, n29853, n29849, n29848, n29847, n29846, 
        n29845, n29844, n29843, n29842, n29841, n29840, n29839, 
        n29837, n29836, n29835, n29834, n29833, n29832, n29831, 
        n29830, n29829, n29828, n29827, n29826, n29825, n29824, 
        n29823, n29822, n29821, n29820, n29819, n29818, n29817, 
        n29816, n29815, n29814, n29813, n29812, n29811, n29810, 
        n29809, n29808, n29807, n29806, n29805, n29804, n29803, 
        n29802, n29801, n29800, n29799, n29797, n29796, n29795, 
        n29794, n29793, n29792, n29791, n29790, n29789, n29788, 
        n29787, n29786, n29785, n29784, n29783, n29782, n29781, 
        n29780, n29779, n29778, n29777, n29775, n29774, n29773, 
        n29772, n56846, n43512, n43510, n29746, n43506, n43402, 
        n29736, n29735, n29734, n29733, n29732, n29731, n5_adj_5709, 
        n524, n523, n522, n521, n29727, n29726, n29725, n29724, 
        n29723, n29722, n29721, n29720, n29719, n29718, n29717, 
        n29716, n29712, n29711, n29708, n29707, n29706, n29705, 
        n29704, n29703, n29702, n29698, n29694, n29691, n29687, 
        n43398, n29684, n29677, n29674, n29673, n29672, n29669, 
        n43494, n29663, n29662, n29661, n43492, n29654, n29648, 
        n29647, n29646, n29644, n29643, n29641, n29639, n29638, 
        n29637, n29636, n29635, n43488, n43486, n29628, n29627, 
        n29626, n29625, n29624, n29617, n29613, n29612, n29608, 
        n29607, n29606, n29605, n29604, n29600, n29594, n29591, 
        n29588, n29579, n57398, n29546, n29543, n29540, n57295, 
        n56101, n56103, n68785, n30_adj_5710, n23_adj_5711, n21_adj_5712, 
        n19_adj_5713, n61472, n520, n4_adj_5714, n3, n2_adj_5715, 
        n17_adj_5716, n16_adj_5717, n15_adj_5718, n13_adj_5719, n11_adj_5720, 
        n10_adj_5721, n9_adj_5722, n8_adj_5723, n7_adj_5724, n6_adj_5725, 
        n4_adj_5726, n61466, n61464, n25424, n61458, n61456, n4_adj_5727, 
        n30741, n4_adj_5728, n30740, n30739, n30655, n30649, n30647, 
        n67639, n10_adj_5729, n61440, n30585, n6_adj_5730, n30569, 
        n30519, n30518, n30517, n30515, n30514, n30513, n30512, 
        n519, n518, n516, control_update;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(35[23:31])
    
    wire n61434, n30506, n30502, n30498, n155, n212, n213, n214, 
        n219;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3715 ;
    
    wire n361, n375, n376, n401, n69366, n455, n456, n12182, 
        n30492, n30488, n8_adj_5731, n6_adj_5732, n30470, n56199, 
        n30468, n30467, n30466, n30465, n15_adj_5733, n11_adj_5734, 
        n30464, n30463, n30462, n30461;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire b_prev, n30460, n30459, n61428, n30458, n30457, position_31__N_3827, 
        n1, n61426, n30456, n30455, n30454, n30453, n30452, n30451, 
        n30450, n30449, n30448, n30447, n30445, n30444, n30443, 
        n30442, n30441, n30440, n49969, n30439;
    wire [1:0]a_new_adj_5954;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire b_prev_adj_5736, position_31__N_3827_adj_5737, n69525, n61420, 
        n12_adj_5738;
    wire [7:0]data_adj_5966;   // verilog/eeprom.v(23[12:16])
    
    wire ready_prev, rw;
    wire [7:0]state_adj_5967;   // verilog/eeprom.v(27[11:16])
    wire [7:0]state_7__N_3916;
    
    wire n61412, n8_adj_5741, n57820, n57818, n57816, n69360, n30406, 
        n30405, n57814, n30404, n57811, n30403, n30402, n30401, 
        n30400, n30399, n30398, n30396, n6617, n30395, n30394, 
        n30393, n49968, n30392, n30391, n30390, n30389, n30388, 
        n30387, n30386, n30385, n30384, n30383, n30375, n25410, 
        n4906, n4905, n61408, clk_out;
    wire [15:0]data_adj_5974;   // verilog/tli4970.v(27[14:18])
    wire [7:0]state_adj_5976;   // verilog/tli4970.v(29[13:18])
    
    wire n19_adj_5752, n18_adj_5753, n17_adj_5754, n4_adj_5755, n3_adj_5756, 
        n2_adj_5757, n57805, n10_adj_5758, n66678, n30350, n30349, 
        n30348, n30347, n30343, n30339, n49967, n61406, n30323, 
        n30322, n30321, n30320, n30319, n30318, n30317, n12190, 
        n12192, n12194, n12196, state_7__N_4317, n30316, n30315, 
        n16_adj_5759, n30308, n43522, n30305, n30299, n8_adj_5760, 
        n25540, n49466, n49465, n29509, n52677, r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(33[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n22849, n12198, n12200, n12202, n12204, n12206, n12208, 
        n12210, n12212, n30282, n30281, n30280, n68450, n61402, 
        n69354, n69348, n69342;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n12214, n12216, n12218, n12220, n15_adj_5761, n14_adj_5762, 
        n13_adj_5763, n12_adj_5764;
    wire [2:0]r_SM_Main_adj_5986;   // verilog/uart_tx.v(32[16:25])
    wire [8:0]r_Clock_Count_adj_5987;   // verilog/uart_tx.v(33[16:29])
    
    wire n49966, n11_adj_5775, n10_adj_5776, n9_adj_5777, n30250, 
        n8_adj_5778, n7_adj_5779, n6_adj_5780, n52657, n30232, n27_adj_5781;
    wire [7:0]state_adj_5997;   // verilog/i2c_controller.v(33[12:17])
    
    wire n4_adj_5783;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire enable_slow_N_4211, n5_adj_5784, n5_adj_5785;
    wire [7:0]state_7__N_4108;
    
    wire n49965, n49964, n6428;
    wire [7:0]state_7__N_4124;
    
    wire n69396, n30221, n30216, n30215, n30214, n30213, n30212, 
        n8_adj_5786, n30211, n30210, n30207, n29499, n30201, n48856, 
        n30200, n29496, n29493, n29490, n56201, n56203, n30196, 
        n49963, n49962, n49464, n18_adj_5787, n30192, n17_adj_5788, 
        n16_adj_5789, n14_adj_5790, n12_adj_5791, n30189, n43524, 
        n49463, n7455, n7454, n7453, n7452, n7451, n7450, n828, 
        n829, n830, n831, n832, n833, n861, n49961, n49960, 
        n896, n897, n898, n899, n900, n901, n49959, n927, n928, 
        n929, n930, n931, n932, n933, n939, n940, n941, n942, 
        n943, n944, n945, n946, n947, n948, n949, n950, n951, 
        n952, n953, n954, n955, n956, n957, n960, n49958, n995, 
        n996, n997, n998, n999, n1000, n1001, n1026, n1027, 
        n1028, n1029, n1030, n1031, n1032, n1033, n1059, n1093, 
        n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, 
        n49957, n1125, n1126, n1127, n1128, n1129, n1130, n1131, 
        n1132, n1133, n42235, n42234, n1158, n61382, n1193, n1194, 
        n1195, n1196, n1197, n1198, n1199, n1200, n1201, n61376, 
        n1224_adj_5792, n1225_adj_5793, n1226_adj_5794, n1227_adj_5795, 
        n1228_adj_5796, n1229_adj_5797, n1230_adj_5798, n1231_adj_5799, 
        n1232_adj_5800, n1233_adj_5801, n1257, n49462, n1292, n1293, 
        n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, 
        n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, 
        n1331, n1332, n1333, n61370, n1356, n49956, n49955, n49954, 
        n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, 
        n1399, n1400, n1401, n49953, n4_adj_5802, n1422, n1423, 
        n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, 
        n1432, n1433, n49952, n1455, n49951, n49461, n1489, n1490, 
        n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, 
        n1499, n1500, n1501, n49950, n49949, n1521, n1522, n1523, 
        n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, 
        n1532, n1533, n67638, n49948, n1554, n25_adj_5803, n1589, 
        n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, 
        n1598, n1599, n1600, n1601, n49460, n1620, n1621, n1622, 
        n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, 
        n1631, n1632, n1633, n1653, n49459, n1688, n1689, n1690, 
        n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, 
        n1699, n1700, n1701, n1719, n1720, n1721, n1722, n1723, 
        n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, 
        n1732, n1733, n41621, n41622, n1752, n1787, n1788_adj_5804, 
        n1789, n1790_adj_5805, n1791, n1792_adj_5806, n1793, n1794_adj_5807, 
        n1795, n1796_adj_5808, n1797, n1798, n1799, n1800, n1801, 
        n61356, n1818, n1819, n1820, n1821, n1822_adj_5809, n1823, 
        n1824_adj_5810, n1825, n1826, n1827, n1828, n1829, n1830, 
        n1831, n1832, n1833, n1851, n490, n61354, n1885, n1886, 
        n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, 
        n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1917, 
        n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, 
        n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, 
        n1950, n49947, n1984, n1985, n1986, n1987, n1988, n1989, 
        n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, 
        n1998, n1999, n2000, n2001, n2016, n2017, n2018, n2019, 
        n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, 
        n2028, n2029, n2030, n2031, n2032, n2033, n68812, n2049, 
        n19_adj_5811, n61348, n20_adj_5812, n2084, n2085, n2086, 
        n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, 
        n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2115, 
        n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, 
        n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, 
        n2132, n2133, n2148, n61344, n2183, n2184, n2185, n2186, 
        n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, 
        n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2214, 
        n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
        n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, 
        n2231, n2232, n2233, n2247, n49648, n49946, n2282, n2283, 
        n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, 
        n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, 
        n2300, n2301, n2313, n2314, n2315, n2316, n2317, n2318, 
        n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, 
        n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2346, 
        n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, 
        n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
        n2397, n2398, n2399, n2400, n2401, n49458, n2412, n2413, 
        n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, 
        n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, 
        n2430, n2431, n2432, n2433, n2445, n40973, n41003, n130, 
        n41018, n61336, n92, n2480, n2481, n2482, n2483, n2484, 
        n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, 
        n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, 
        n2501, n2511, n2512, n2513, n2514, n2515, n2516, n2517, 
        n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, 
        n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, 
        n2544, n49945, n67642, n2579, n2580, n2581, n2582, n2583, 
        n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, 
        n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, 
        n2600, n2601, n2610, n2611, n2612, n2613, n2614, n2615, 
        n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, 
        n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, 
        n2632, n2633, n2643, n61332, n49944, n61330, n2677, n2678, 
        n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, 
        n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, 
        n2695, n2696, n2697, n2698, n2699, n2700, n2701, n61328, 
        n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, 
        n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, 
        n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, 
        n2733, n2742, n172, n49943, n42632, n2777, n2778, n2779, 
        n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, 
        n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, 
        n2796, n2797, n2798, n2799, n2800, n2801, n2808, n2809, 
        n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, 
        n2818, n2819, n2820_adj_5813, n2821, n2822, n2823, n2824, 
        n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, 
        n2833, n2841, n2876, n2877, n2878, n2879, n2880, n2881, 
        n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, 
        n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, 
        n2898, n2899, n2900, n2901, n2907, n2908, n2909, n2910, 
        n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, 
        n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, 
        n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2940, 
        n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, 
        n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, 
        n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, 
        n2998, n2999, n3000, n3001, n49647, n3006, n3007, n3008, 
        n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, 
        n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, 
        n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, 
        n3033, n3039, n111, n134, n417, n142, n3074, n3075, 
        n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, 
        n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, 
        n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, 
        n3100, n3101, n49457, n3105, n3106, n3107, n3108, n3109, 
        n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, 
        n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, 
        n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, 
        n3138, n111_adj_5814, n61314, n3173, n3174, n3175, n3176, 
        n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, 
        n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, 
        n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, 
        n3201, n3204, n3205, n3206, n3207, n3208, n3209, n3210, 
        n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, 
        n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, 
        n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3237, 
        n69489, n3272, n3273, n3274, n3275, n3276, n3277, n3278, 
        n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, 
        n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, 
        n3295, n3296, n69309, n3298, n3301, n61308, n4_adj_5815, 
        n61300, n20194, n24_adj_5816, n61292, n62, n49456, n61286, 
        n49646, n49942, n61282, n61276, n49941, n61274, n27997, 
        n30186, n61262, n27966, n65997, n68763, n43, n45, n49940, 
        n61256, n49455, n49645, n49454, n49453, n49939, n61250, 
        n57701, n49644, n49938, n49643, n49937, n49452, n52803, 
        n30182, n61248, n49936, n49935, n30179, n60010, n27920, 
        n61242, n30176, n49934, n49933, n49642, n30172, n30169, 
        n30166, n49641, n49640, n49451, n49639, n49450, n49932, 
        n49638, n49931, n49930, n61238, n49449, n49929, n49928, 
        n61236, n49637, n25404, n30156, n30155, n49927, n49636, 
        n30152, n49926, n49925, n30149, n49635, n27780, n49924, 
        n49923, n49922, n49921, n27724, n61224, n65995, n61222, 
        n4_adj_5817, n4_adj_5818, n30_adj_5819, n32_adj_5820, n4_adj_5821, 
        n69078, n68734, n56425, n27706, n61220, n61218, n27698, 
        n27696, n27692, n61216, n58789, n61214, n49920, n49919, 
        n49918, n49917, n61212, n61210, n344, n61208, n61206, 
        n61204, n49916, n61202, n61200, n271, n61196, n49915, 
        n49914, n49913, n49912, n49911, n61188, n49910, n61186, 
        n61184, n27646, n61182, n61180, n65985, n14_adj_5822, n49909, 
        n49908, n10_adj_5823, n61176, n65983, n49907, n198, n204, 
        n61170, n49906, n42779, n69065, n49905, n27622, n61162, 
        n61160, n69306, n49904, n49903, n66513, n66511, n131, 
        n61154, n125, n61148, n110, n66503, n68512, n49902, n49901, 
        n49163, n61138, n6_adj_5824, n49900, n49899, n56, n53, 
        n38, n61132, n57125, n49898, n50393, n49897, n69051, n43_adj_5825, 
        n37189, n61126, n50392, n49896, n6_adj_5826, n49895, n50391, 
        n50390, n50389, n61120, n61118, n50388, n49894, n49893, 
        n50387, n49892, n26482, n49891, n61104, n59230, n49890, 
        n61098, n61096, n61090, n6_adj_5827, n61086, n49889, n61078, 
        n57473, n49888, n49887, n61074, n25571, n61068, n61060, 
        n61054, n61048, n49886, n4_adj_5828, n6_adj_5829, n8_adj_5830, 
        n9_adj_5831, n4_adj_5832, n6_adj_5833, n8_adj_5834, n9_adj_5835, 
        n11_adj_5836, n13_adj_5837, n15_adj_5838, n49885, n49884, 
        n49883, n49882, n61042, n25535, n38_adj_5839, n39, n40, 
        n41, n42, n43_adj_5840, n44, n45_adj_5841, n29480, n29478, 
        n49881, n11610, n11579, n11577, n49880, n49879, n57012, 
        n49878, n61036, n67761, n4_adj_5842, n61032, n60042, n61030, 
        n5_adj_5843, n53307, n29162, n57467, n56952, n56951, n56950, 
        n56949, n56948, n56947, n56946, n56945, n56944, n56943, 
        n56942, n56941, n56772, n56940, n29117, n29116, n29115, 
        n56939, n56938, n56937, n56936, n56935, n56934, n56933, 
        n56932, n56931, n56930, n56929, n56928, n56927, n56926, 
        n56925, n56924, n56923, n56922, n56921, n56920, n57044, 
        n57039, n28438, n28436, n28434, n28428, n59575, n28417, 
        n28885, n28878, n28387, n28383, n28381, n28379, n28375, 
        n61018, n69005, n49877, n61012, n10_adj_5844, n49876, n69456, 
        n49875, n49610, n3_adj_5845, n49874, n49873, n49872, n49162, 
        n49871, n49609, n49608, n49870, n49607, n49869, n49606, 
        n49868, n24_adj_5846, n22_adj_5847, n22726, n49605, n20_adj_5848, 
        n56057, n20195, n56919, n16_adj_5849, n58643, n25527, n49604, 
        n49603, n49867, n25532, n20196, n61002, n69032, n49602, 
        n49161, n62508, n49866, n25519, n49601, n49865, n49864, 
        n30095, n30092, n30089, n30085, n30082, n30079, n49160, 
        n49600, n49863, n49599, n20149, n30075, n30072, n30069, 
        n43588, n30066, n43586, n30063, n43584, n30057, n30054, 
        n30050, n43578, n30047, n21_adj_5850, n66254, n68442, n58718, 
        n58714, n49862, n43576, n43572, n43570, n43566, n49598, 
        n49861, n43560, n49860, n52851, n49859, n43552, n43550, 
        n29995, n29992, n43546, n29989, n29986, n43542, n29982, 
        n29979, n29976, n29973, n49151, n49858, n49857, n49856, 
        n49159, n49855, n49854, n49853, n49852, n49851, n49850, 
        n49849, n49848, n49847, n49846, n49845, n68703, n49844, 
        n66233, n49843, n2_adj_5851, n3_adj_5852, n4_adj_5853, n5_adj_5854, 
        n6_adj_5855, n7_adj_5856, n8_adj_5857, n9_adj_5858, n10_adj_5859, 
        n11_adj_5860, n12_adj_5861, n13_adj_5862, n14_adj_5863, n15_adj_5864, 
        n16_adj_5865, n17_adj_5866, n18_adj_5867, n19_adj_5868, n20_adj_5869, 
        n21_adj_5870, n22_adj_5871, n23_adj_5872, n24_adj_5873, n25_adj_5874, 
        n26_adj_5875, n27_adj_5876, n28_adj_5877, n29_adj_5878, n30_adj_5879, 
        n31_adj_5880, n32_adj_5881, n66231, n49842, n49841, n49840, 
        n49839, n49838, n49837, n49415, n49414, n49836, n49581, 
        n49835, n49413, n49580, n49579, n49834, n49833, n49832, 
        n49412, n49150, n49578, n49577, n49576, n49575, n49574, 
        n49573, n49411, n49410, n49409, n49572, n49408, n49571, 
        n49407, n49570, n49406, n49405, n69450, n49404, n49286, 
        n49403, n49285, n49402, n49809, n49284, n49401, n49400, 
        n49808, n49807, n49806, n49283, n49805, n49399, n57812, 
        n49158, n49282, n49398, n49281, n49397, n49804, n49280, 
        n6_adj_5882, n49803, n49396, n49395, n49548, n49547, n49279, 
        n49546, n49278, n49802, n49801, n4_adj_5883, n49394, n49393, 
        n49392, n49545, n49800, n49391, n49390, n49544, n49157, 
        n49277, n49389, n49799, n49798, n62712, n49543, n49276, 
        n49797, n49542, n49388, n49541, n49275, n49796, n49387, 
        n49795, n49540, n49539, n49794, n49793, n49274, n49538, 
        n49273, n49792, n49386, n49272, n49385, n49271, n49384, 
        n49383, n49270, n49382, n49269, n49149, n66181, n49381, 
        n49380, n49268, n49267, n49266, n66171, n49265, n49156, 
        n50149, n50148, n50147, n49264, n50146, n50145, n50144, 
        n50143, n12_adj_5884, n50142, n50141, n50140, n50139, n50138, 
        n50137, n50136, n50135, n50134, n49523, n50133, n66144, 
        n49761, n50132, n50131, n49760, n50130, n50129, n49522, 
        n49759, n49758, n49521, n49520, n49757, n17_adj_5885, n19_adj_5886, 
        n50128, n21_adj_5887, n27_adj_5888, n29_adj_5889, n33, n59, 
        n61, n49756, n50127, n69444, n49755, n50126, n49754, n50125, 
        n50124, n49155, n50123, n50122, n49177, n49753, n49148, 
        n50121, n50120, n49752, n49751, n50119, n49519, n49750, 
        n50118, n49176, n49518, n49517, n49516, n50117, n49175, 
        n49515, n49749, n50116, n50115, n56918, n49514, n49748, 
        n49747, n20894, n20890, n49746, n50114, n20222, n33761, 
        n49745, n49174, n62711, n69682, n61740, n56917, n57717, 
        n61732, n56777, n56916, n56915, n56914, n33769, n61726, 
        n61720, n61714, n56913, n11642, n25422, n25507, n51730, 
        n68676, n26524, n62627, n61708, n50113, n59574, n50112, 
        n49173, n62858, n50111, n49147, n50110, n25523, n50109, 
        n65487, n49172, n20151, n25530, n12_adj_5890, n20150, n50108, 
        n50107, n50106, n51676, n50105, n51654, n68255, n50104, 
        n61702, n51640, n69438, n65486, n61700, n67727, n6_adj_5891, 
        n61696, n69432, n68312, n60804, n68943, n68643, n51598, 
        n67757, n59242, n50103, n65481, n60788, n68923, n60772, 
        n56959, n67787, n68025, n65447, n60756, n65444, n6_adj_5892, 
        n4_adj_5893, n60740, n65441, n55331, n5_adj_5894, n24_adj_5895, 
        n60724, n17_adj_5896, n25_adj_5897, n7_adj_5898, n69426, n65437, 
        n60708, n65436, n65433, n65432, n55417, n60692, n10_adj_5899, 
        n61684, n6_adj_5900, n68902, n67051, n58681, n14_adj_5901, 
        n10_adj_5902, n67477, n65412, n67471, n56771, n57131, n65411, 
        n10_adj_5903, n67475, n57629, n59193, n65401, n57720, n60070, 
        n57377, n57350, n5_adj_5904, n67017, n69420, n68319, n57768, 
        n59466, n5_adj_5905, n59858, n57741, n57516, n25_adj_5906, 
        n57780, n57361, n68609, n58765, n68881, n4_adj_5907, n62365, 
        n15_adj_5908, n14_adj_5909, n57232, n58640, n55999, n56027, 
        n56031, n56037, n56041, n56045, n56049, n69414, n56053, 
        n62859, n56061, n56065, n56071, n57503, n56075, n56079, 
        n56083, n56087, n56091, n56095, n57680, n56099, n56107, 
        n9_adj_5910, n65309, n59636, n8_adj_5911, n68857, n12_adj_5912, 
        n65285, n69408, n56249, n68339, n68335, n67043, n56303, 
        n56343, n62633, n62631, n58740, n62630, n56988, n58638, 
        n60174, n57456, n68263, n68262, n68256, n23_adj_5913, n8_adj_5914, 
        n7_adj_5915, n68583, n67067, n58743, n68182, n68257, n68074, 
        n68174, n69402, n7_adj_5916, n69390;
    
    VCC i2 (.Y(VCC_net));
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(clk16MHz), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF dir_183 (.Q(dir), .C(clk16MHz), .D(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_add_1503_20_lut (.I0(GND_net), .I1(n2216), 
            .I2(VCC_net), .I3(n49868), .O(n2283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_20_lut.LUT_INIT = 16'hC33C;
    SB_DFFE dti_185 (.Q(dti), .C(clk16MHz), .E(n27622), .D(dti_N_404));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[0]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_add_1034_4_lut (.I0(GND_net), .I1(n1532), 
            .I2(GND_net), .I3(n49599), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[0]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(clk16MHz), 
           .D(encoder1_position[2]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk16MHz), .D(displacement_23__N_67[0]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4124[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_30__I_0_add_1503_20 (.CI(n49868), .I0(n2216), 
            .I1(VCC_net), .CO(n49869));
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.timer({timer}), .GND_net(GND_net), 
            .clk16MHz(clk16MHz), .state({state}), .n25(n25_adj_5906), 
            .VCC_net(VCC_net), .bit_ctr({Open_0, Open_1, Open_2, bit_ctr[1:0]}), 
            .neopxl_color({neopxl_color}), .n111(n111), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .n29677(n29677), .n27920(n27920), .n30323(n30323), .n30322(n30322), 
            .n30321(n30321), .n30320(n30320), .n30319(n30319), .n30318(n30318), 
            .n30317(n30317), .n30316(n30316), .n30315(n30315), .n30308(n30308), 
            .n30221(n30221), .n5(n5_adj_5904), .NEOPXL_c(NEOPXL_c), .LED_c(LED_c), 
            .n43462(n43462), .n23(n23_adj_5913)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(51[24] 57[2])
    SB_CARRY encoder0_position_30__I_0_add_1034_4 (.CI(n49599), .I0(n1532), 
            .I1(GND_net), .CO(n49600));
    SB_LUT4 encoder0_position_30__I_0_add_1034_3_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n49598), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_3 (.CI(n49598), .I0(n1533), 
            .I1(VCC_net), .CO(n49599));
    SB_LUT4 encoder0_position_30__I_0_add_1503_19_lut (.I0(GND_net), .I1(n2217), 
            .I2(VCC_net), .I3(n49867), .O(n2284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_19_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i22 (.Q(delay_counter[22]), .C(clk16MHz), .E(n27698), 
            .D(n1217), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i6_4_lut (.I0(n57768), .I1(n57232), .I2(n57629), .I3(\data_out_frame[23] [2]), 
            .O(n14_adj_5822));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(n52677), .I1(n14_adj_5822), .I2(n10_adj_5823), 
            .I3(n57295), .O(n51598));
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\data_out_frame[18] [3]), .I1(n59193), .I2(n52803), 
            .I3(n51654), .O(n57768));
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[22] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n57629));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_2_lut (.I0(n51730), .I1(\data_out_frame[22] [6]), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_5849));
    defparam i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut (.I0(n68335), .I1(n57377), .I2(n57741), .I3(\data_out_frame[14] [4]), 
            .O(n22_adj_5847));
    defparam i9_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i11_4_lut (.I0(n51640), .I1(n22_adj_5847), .I2(n16_adj_5849), 
            .I3(n57768), .O(n24_adj_5846));
    defparam i11_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut (.I0(\data_out_frame[19] [3]), .I1(n24_adj_5846), 
            .I2(n20_adj_5848), .I3(\data_out_frame[18] [7]), .O(n52657));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut (.I0(\data_out_frame[16] [4]), .I1(n57398), .I2(n25_adj_5803), 
            .I3(\data_out_frame[16] [5]), .O(n12_adj_5884));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1818 (.I0(n59466), .I1(n12_adj_5884), .I2(\data_out_frame[21] [0]), 
            .I3(\data_out_frame[18] [6]), .O(n57350));
    defparam i6_4_lut_adj_1818.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut (.I0(state_adj_5967[2]), .I1(state_adj_5967[1]), .I2(state_adj_5967[0]), 
            .I3(n42699), .O(n55999));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_4_lut.LUT_INIT = 16'ha8e8;
    SB_LUT4 i15596_4_lut (.I0(CS_MISO_c), .I1(data_adj_5974[1]), .I2(n6), 
            .I3(n25519), .O(n29604));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15596_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15597_4_lut (.I0(CS_MISO_c), .I1(data_adj_5974[2]), .I2(n5_adj_5784), 
            .I3(n25527), .O(n29605));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15597_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15598_4_lut (.I0(CS_MISO_c), .I1(data_adj_5974[3]), .I2(n42774), 
            .I3(n25527), .O(n29606));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15598_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15599_4_lut (.I0(CS_MISO_c), .I1(data_adj_5974[4]), .I2(n6_adj_5732), 
            .I3(n25571), .O(n29607));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15599_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15600_4_lut (.I0(CS_MISO_c), .I1(data_adj_5974[5]), .I2(n6_adj_5732), 
            .I3(n25519), .O(n29608));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15600_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15604_4_lut (.I0(CS_MISO_c), .I1(data_adj_5974[6]), .I2(n5_adj_5784), 
            .I3(n4_adj_5783), .O(n29612));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15604_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15609_4_lut (.I0(CS_MISO_c), .I1(data_adj_5974[7]), .I2(n6_adj_5732), 
            .I3(n25532), .O(n29617));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15609_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15616_4_lut (.I0(CS_MISO_c), .I1(data_adj_5974[8]), .I2(n5_adj_5708), 
            .I3(n25523), .O(n29624));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15616_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15617_4_lut (.I0(CS_MISO_c), .I1(data_adj_5974[9]), .I2(n6_adj_5730), 
            .I3(n25519), .O(n29625));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15617_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15618_4_lut (.I0(CS_MISO_c), .I1(data_adj_5974[10]), .I2(n5_adj_5784), 
            .I3(n25523), .O(n29626));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15618_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15876_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n60724), 
            .I3(n27_adj_5781), .O(n29884));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15876_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15619_4_lut (.I0(CS_MISO_c), .I1(data_adj_5974[11]), .I2(n42774), 
            .I3(n25523), .O(n29627));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15619_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15620_4_lut (.I0(CS_MISO_c), .I1(data_adj_5974[12]), .I2(n42779), 
            .I3(n25571), .O(n29628));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15620_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15629_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n22726), .I3(GND_net), .O(n29637));   // verilog/coms.v(130[12] 305[6])
    defparam i15629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15633_3_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .I2(control_update), .I3(GND_net), .O(n29641));   // verilog/motorControl.v(41[14] 62[8])
    defparam i15633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15635_4_lut (.I0(CS_MISO_c), .I1(data_adj_5974[15]), .I2(n42779), 
            .I3(n25532), .O(n29643));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15635_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i11_2_lut (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[18] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n25810));   // verilog/coms.v(100[12:26])
    defparam i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(\data_out_frame[19] [4]), .I1(n68339), .I2(n57456), 
            .I3(n6_adj_5824), .O(n57741));
    defparam i4_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1819 (.I0(state_adj_5967[2]), .I1(data_ready), 
            .I2(n3_adj_5845), .I3(n25516), .O(n56425));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_4_lut_adj_1819.LUT_INIT = 16'hcca8;
    SB_LUT4 i15638_3_lut (.I0(current[0]), .I1(data_adj_5974[0]), .I2(n27706), 
            .I3(GND_net), .O(n29646));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15639_4_lut (.I0(rw), .I1(state_adj_5967[1]), .I2(state_adj_5967[2]), 
            .I3(n5774), .O(n29647));   // verilog/eeprom.v(35[8] 81[4])
    defparam i15639_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i15640_3_lut (.I0(CS_c), .I1(state_adj_5976[0]), .I2(state_adj_5976[1]), 
            .I3(GND_net), .O(n29648));   // verilog/tli4970.v(35[10] 68[6])
    defparam i15640_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 i53466_4_lut (.I0(n15_adj_5733), .I1(clk_out), .I2(state_adj_5976[0]), 
            .I3(state_adj_5976[1]), .O(n9_adj_5910));   // verilog/tli4970.v(35[10] 68[6])
    defparam i53466_4_lut.LUT_INIT = 16'hc8fc;
    SB_DFFESR delay_counter__i23 (.Q(delay_counter[23]), .C(clk16MHz), .E(n27698), 
            .D(n1216), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i24 (.Q(delay_counter[24]), .C(clk16MHz), .E(n27698), 
            .D(n1215), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i25 (.Q(delay_counter[25]), .C(clk16MHz), .E(n27698), 
            .D(n1214), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i26 (.Q(delay_counter[26]), .C(clk16MHz), .E(n27698), 
            .D(n1213), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i27 (.Q(delay_counter[27]), .C(clk16MHz), .E(n27698), 
            .D(n1212), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i28 (.Q(delay_counter[28]), .C(clk16MHz), .E(n27698), 
            .D(n1211), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i29 (.Q(delay_counter[29]), .C(clk16MHz), .E(n27698), 
            .D(n1210), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i30 (.Q(delay_counter[30]), .C(clk16MHz), .E(n27698), 
            .D(n1209), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i31 (.Q(delay_counter[31]), .C(clk16MHz), .E(n27698), 
            .D(n1208), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i15646_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(n57012), .I3(state_7__N_4108[0]), 
            .O(n29654));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15646_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i1_2_lut_adj_1820 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5803));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1820.LUT_INIT = 16'h6666;
    SB_LUT4 i15664_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n22726), .I3(GND_net), .O(n29672));   // verilog/coms.v(130[12] 305[6])
    defparam i15664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15665_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n22726), .I3(GND_net), .O(n29673));   // verilog/coms.v(130[12] 305[6])
    defparam i15665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1171_3_lut (.I0(n1720), .I1(n1787), 
            .I2(n1752), .I3(GND_net), .O(n1819));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15669_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n29677));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15669_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i46947_3_lut (.I0(n4908), .I1(duty[20]), .I2(n11579), .I3(GND_net), 
            .O(n62633));
    defparam i46947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1238_3_lut (.I0(n1819), .I1(n1886), 
            .I2(n1851), .I3(GND_net), .O(n1918));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1305_3_lut (.I0(n1918), .I1(n1985), 
            .I2(n1950), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i46949_3_lut (.I0(n62633), .I1(n62631), .I2(n11577), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[20]));
    defparam i46949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46944_3_lut (.I0(n4907), .I1(duty[21]), .I2(n11579), .I3(GND_net), 
            .O(n62630));
    defparam i46944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46946_3_lut (.I0(n62630), .I1(n62631), .I2(n11577), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[21]));
    defparam i46946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46945_3_lut (.I0(current[15]), .I1(duty[23]), .I2(n11579), 
            .I3(GND_net), .O(n62631));
    defparam i46945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46941_3_lut (.I0(n4906), .I1(duty[22]), .I2(n11579), .I3(GND_net), 
            .O(n62627));
    defparam i46941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46943_3_lut (.I0(n62627), .I1(n62631), .I2(n11577), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[22]));
    defparam i46943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7213_3_lut (.I0(n4905), .I1(current[15]), .I2(n11577), .I3(GND_net), 
            .O(n20894));
    defparam i7213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7214_3_lut (.I0(n20894), .I1(duty[23]), .I2(n11579), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[23]));
    defparam i7214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1372_3_lut (.I0(n2017), .I1(n2084), 
            .I2(n2049), .I3(GND_net), .O(n2116));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7468_2_lut (.I0(hall3), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(n20890));   // verilog/TinyFPGA_B.v(160[4] 162[7])
    defparam i7468_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i8783_2_lut (.I0(hall3), .I1(hall1), .I2(GND_net), .I3(GND_net), 
            .O(commutation_state_7__N_27[2]));   // verilog/TinyFPGA_B.v(166[4] 168[7])
    defparam i8783_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i42177_3_lut (.I0(n4_adj_5907), .I1(commutation_state_7__N_27[2]), 
            .I2(commutation_state[2]), .I3(GND_net), .O(n57805));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i42177_3_lut.LUT_INIT = 16'hdcdc;
    SB_LUT4 i15683_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n22726), .I3(GND_net), .O(n29691));   // verilog/coms.v(130[12] 305[6])
    defparam i15683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15686_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n22726), .I3(GND_net), .O(n29694));   // verilog/coms.v(130[12] 305[6])
    defparam i15686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29643_4_lut (.I0(n519), .I1(n831), .I2(n832), .I3(n833), 
            .O(n43552));
    defparam i29643_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i15690_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n22726), .I3(GND_net), .O(n29698));   // verilog/coms.v(130[12] 305[6])
    defparam i15690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23859_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n22726), .I3(GND_net), .O(n29702));
    defparam i23859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1821 (.I0(n36759), .I1(Ki[3]), .I2(GND_net), 
            .I3(GND_net), .O(n271));
    defparam i1_2_lut_adj_1821.LUT_INIT = 16'h8888;
    SB_LUT4 i15695_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n22726), .I3(GND_net), .O(n29703));   // verilog/coms.v(130[12] 305[6])
    defparam i15695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15877_3_lut (.I0(\data_in_frame[1] [6]), .I1(rx_data[6]), .I2(n57044), 
            .I3(GND_net), .O(n29885));   // verilog/coms.v(130[12] 305[6])
    defparam i15877_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1584_i10_3_lut (.I0(duty[12]), .I1(duty[9]), .I2(n260), 
            .I3(GND_net), .O(n12208));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(current[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5677));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1822 (.I0(n36759), .I1(Ki[4]), .I2(GND_net), 
            .I3(GND_net), .O(n344));
    defparam i1_2_lut_adj_1822.LUT_INIT = 16'h8888;
    SB_LUT4 i28718_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(90[16:31])
    defparam i28718_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i28835_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(88[16:31])
    defparam i28835_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_add_1034_2_lut (.I0(GND_net), .I1(n940), 
            .I2(GND_net), .I3(VCC_net), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(current[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_5676));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1823 (.I0(n36759), .I1(Ki[5]), .I2(GND_net), 
            .I3(GND_net), .O(n417));
    defparam i1_2_lut_adj_1823.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_1824 (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), 
            .I2(delay_counter[31]), .I3(\ID_READOUT_FSM.state [0]), .O(n60174));
    defparam i3_4_lut_adj_1824.LUT_INIT = 16'h0004;
    SB_LUT4 i15679_3_lut (.I0(\data_in_frame[22] [6]), .I1(rx_data[6]), 
            .I2(n28428), .I3(GND_net), .O(n29687));   // verilog/coms.v(130[12] 305[6])
    defparam i15679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15703_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n22726), .I3(GND_net), .O(n29711));   // verilog/coms.v(130[12] 305[6])
    defparam i15703_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15881_3_lut (.I0(\data_in_frame[1] [7]), .I1(rx_data[7]), .I2(n57044), 
            .I3(GND_net), .O(n29889));   // verilog/coms.v(130[12] 305[6])
    defparam i15881_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15710_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n22726), .I3(GND_net), .O(n29718));   // verilog/coms.v(130[12] 305[6])
    defparam i15710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15711_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n22726), .I3(GND_net), .O(n29719));   // verilog/coms.v(130[12] 305[6])
    defparam i15711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29757_4_lut (.I0(n829), .I1(n828), .I2(n43552), .I3(n830), 
            .O(n861));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i29757_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i15712_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n22726), .I3(GND_net), .O(n29720));   // verilog/coms.v(130[12] 305[6])
    defparam i15712_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15713_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n22726), .I3(GND_net), .O(n29721));   // verilog/coms.v(130[12] 305[6])
    defparam i15713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1825 (.I0(n36694), .I1(Ki[2]), .I2(GND_net), 
            .I3(GND_net), .O(n204));
    defparam i1_2_lut_adj_1825.LUT_INIT = 16'h8888;
    SB_CARRY encoder0_position_30__I_0_add_1034_2 (.CI(VCC_net), .I0(n940), 
            .I1(GND_net), .CO(n49598));
    SB_LUT4 i1_2_lut_adj_1826 (.I0(n36694), .I1(Ki[1]), .I2(GND_net), 
            .I3(GND_net), .O(n131));
    defparam i1_2_lut_adj_1826.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(current[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5675));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15676_3_lut (.I0(\data_in_frame[22] [5]), .I1(rx_data[5]), 
            .I2(n28428), .I3(GND_net), .O(n29684));   // verilog/coms.v(130[12] 305[6])
    defparam i15676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22725_3_lut (.I0(n212), .I1(IntegralLimit[19]), .I2(n155), 
            .I3(GND_net), .O(n36694));
    defparam i22725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22755_3_lut (.I0(n213), .I1(IntegralLimit[18]), .I2(n155), 
            .I3(GND_net), .O(n36723));
    defparam i22755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1827 (.I0(n36759), .I1(Ki[6]), .I2(GND_net), 
            .I3(GND_net), .O(n490));
    defparam i1_2_lut_adj_1827.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(current[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5674));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i42182_3_lut (.I0(n3), .I1(n7451), .I2(n57811), .I3(GND_net), 
            .O(n57812));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42182_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1503_19 (.CI(n49867), .I0(n2217), 
            .I1(VCC_net), .CO(n49868));
    SB_LUT4 encoder0_position_30__I_0_add_1503_18_lut (.I0(GND_net), .I1(n2218), 
            .I2(VCC_net), .I3(n49866), .O(n2285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i42183_3_lut (.I0(encoder0_position[29]), .I1(n57812), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n829));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_5881));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29641_4_lut (.I0(n520), .I1(n931), .I2(n932), .I3(n933), 
            .O(n43550));
    defparam i29641_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i15714_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n22726), .I3(GND_net), .O(n29722));   // verilog/coms.v(130[12] 305[6])
    defparam i15714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15715_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n22726), .I3(GND_net), .O(n29723));   // verilog/coms.v(130[12] 305[6])
    defparam i15715_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1503_18 (.CI(n49866), .I0(n2218), 
            .I1(VCC_net), .CO(n49867));
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[1]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i15717_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n22726), .I3(GND_net), .O(n29725));   // verilog/coms.v(130[12] 305[6])
    defparam i15717_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[3]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_5880));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1584_i11_3_lut (.I0(duty[13]), .I1(duty[10]), .I2(n260), 
            .I3(GND_net), .O(n12206));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_5879));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1828 (.I0(\data_out_frame[7] [3]), .I1(n57516), 
            .I2(GND_net), .I3(GND_net), .O(n26524));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1828.LUT_INIT = 16'h6666;
    SB_LUT4 i15718_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n22726), .I3(GND_net), .O(n29726));   // verilog/coms.v(130[12] 305[6])
    defparam i15718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_5878));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15719_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n22726), .I3(GND_net), .O(n29727));   // verilog/coms.v(130[12] 305[6])
    defparam i15719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_add_1503_17_lut (.I0(GND_net), .I1(n2219), 
            .I2(VCC_net), .I3(n49865), .O(n2286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_17 (.CI(n49865), .I0(n2219), 
            .I1(VCC_net), .CO(n49866));
    SB_LUT4 encoder0_position_30__I_0_add_1503_16_lut (.I0(GND_net), .I1(n2220), 
            .I2(VCC_net), .I3(n49864), .O(n2287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_5877));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 n11579_bdd_4_lut (.I0(n11579), .I1(current[15]), .I2(duty[22]), 
            .I3(n11577), .O(n69456));
    defparam n11579_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_CARRY encoder0_position_30__I_0_add_1503_16 (.CI(n49864), .I0(n2220), 
            .I1(VCC_net), .CO(n49865));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_5876));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[19]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 n69456_bdd_4_lut (.I0(n69456), .I1(duty[19]), .I2(n4909), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[19]));
    defparam n69456_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_5875));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5874));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1503_15_lut (.I0(GND_net), .I1(n2221), 
            .I2(VCC_net), .I3(n49863), .O(n2288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_15_lut.LUT_INIT = 16'hC33C;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(clk16MHz));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[2]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_in_frame[8] [6]), .I1(n57680), .I2(n25952), 
            .I3(GND_net), .O(Kp_23__N_1301));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[8] [6]), .I1(n57680), .I2(\data_in_frame[13] [5]), 
            .I3(n10_adj_5899), .O(n59636));   // verilog/coms.v(99[12:25])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY encoder0_position_30__I_0_add_1503_15 (.CI(n49863), .I0(n2221), 
            .I1(VCC_net), .CO(n49864));
    SB_LUT4 encoder0_position_30__I_0_add_1503_14_lut (.I0(GND_net), .I1(n2222), 
            .I2(VCC_net), .I3(n49862), .O(n2289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5873));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_151_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n49149), .O(n1236)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[5] [1]), .I3(GND_net), .O(n57516));   // verilog/coms.v(100[12:26])
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_CARRY encoder0_position_30__I_0_add_1503_14 (.CI(n49862), .I0(n2222), 
            .I1(VCC_net), .CO(n49863));
    SB_LUT4 encoder0_position_30__I_0_add_1503_13_lut (.I0(GND_net), .I1(n2223), 
            .I2(VCC_net), .I3(n49861), .O(n2290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_14 (.CI(n49158), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n49159));
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[23]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_CARRY encoder0_position_30__I_0_add_1503_13 (.CI(n49861), .I0(n2223), 
            .I1(VCC_net), .CO(n49862));
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(current[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5673));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[22]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_add_1503_12_lut (.I0(GND_net), .I1(n2224), 
            .I2(VCC_net), .I3(n49860), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[21]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[20]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5872));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1503_12 (.CI(n49860), .I0(n2224), 
            .I1(VCC_net), .CO(n49861));
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[19]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_add_1503_11_lut (.I0(GND_net), .I1(n2225), 
            .I2(VCC_net), .I3(n49859), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_11_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[18]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_CARRY encoder0_position_30__I_0_add_1503_11 (.CI(n49859), .I0(n2225), 
            .I1(VCC_net), .CO(n49860));
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(current[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n49415), .O(n294)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[17]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[16]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 add_151_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n49157), .O(n1228)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[15]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[14]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[13]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_add_1503_10_lut (.I0(GND_net), .I1(n2226), 
            .I2(VCC_net), .I3(n49858), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_10 (.CI(n49858), .I0(n2226), 
            .I1(VCC_net), .CO(n49859));
    SB_LUT4 encoder0_position_30__I_0_add_1503_9_lut (.I0(GND_net), .I1(n2227), 
            .I2(VCC_net), .I3(n49857), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_9 (.CI(n49857), .I0(n2227), 
            .I1(VCC_net), .CO(n49858));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5871));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_967_14_lut (.I0(GND_net), .I1(n1422), 
            .I2(VCC_net), .I3(n49581), .O(n1489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_14_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[12]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_add_967_13_lut (.I0(GND_net), .I1(n1423), 
            .I2(VCC_net), .I3(n49580), .O(n1490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[11]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_add_1503_8_lut (.I0(GND_net), .I1(n2228), 
            .I2(VCC_net), .I3(n49856), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(clk16MHz), .D(encoder0_position_scaled_23__N_43[10]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[9]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[8]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_CARRY encoder0_position_30__I_0_add_1503_8 (.CI(n49856), .I0(n2228), 
            .I1(VCC_net), .CO(n49857));
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[7]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 encoder0_position_30__I_0_add_1503_7_lut (.I0(GND_net), .I1(n2229), 
            .I2(GND_net), .I3(n49855), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[6]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[5]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[4]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[3]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[2]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 n11579_bdd_4_lut_53716 (.I0(n11579), .I1(current[15]), .I2(duty[21]), 
            .I3(n11577), .O(n69450));
    defparam n11579_bdd_4_lut_53716.LUT_INIT = 16'he4aa;
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(clk16MHz), 
           .D(encoder0_position_scaled_23__N_43[1]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n49414), .O(n298)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_13 (.CI(n49580), .I0(n1423), 
            .I1(VCC_net), .CO(n49581));
    SB_CARRY encoder0_position_30__I_0_add_1503_7 (.CI(n49855), .I0(n2229), 
            .I1(GND_net), .CO(n49856));
    SB_LUT4 encoder0_position_30__I_0_add_1503_6_lut (.I0(GND_net), .I1(n2230), 
            .I2(GND_net), .I3(n49854), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n49414), .I0(GND_net), .I1(n2), 
            .CO(n49415));
    SB_LUT4 encoder0_position_30__I_0_add_967_12_lut (.I0(GND_net), .I1(n1424), 
            .I2(VCC_net), .I3(n49579), .O(n1491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n69450_bdd_4_lut (.I0(n69450), .I1(duty[18]), .I2(n4910), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[18]));
    defparam n69450_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY encoder0_position_30__I_0_add_1503_6 (.CI(n49854), .I0(n2230), 
            .I1(GND_net), .CO(n49855));
    SB_CARRY encoder0_position_30__I_0_add_967_12 (.CI(n49579), .I0(n1424), 
            .I1(VCC_net), .CO(n49580));
    SB_LUT4 encoder0_position_30__I_0_add_967_11_lut (.I0(GND_net), .I1(n1425), 
            .I2(VCC_net), .I3(n49578), .O(n1492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_5_lut (.I0(GND_net), .I1(n2231), 
            .I2(VCC_net), .I3(n49853), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5870));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5869));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1584_i12_3_lut (.I0(duty[14]), .I1(duty[11]), .I2(n260), 
            .I3(GND_net), .O(n12204));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5868));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5867));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5866));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15728_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n22726), .I3(GND_net), .O(n29736));   // verilog/coms.v(130[12] 305[6])
    defparam i15728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5865));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5864));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5863));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5862));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5861));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1503_5 (.CI(n49853), .I0(n2231), 
            .I1(VCC_net), .CO(n49854));
    SB_CARRY encoder0_position_30__I_0_add_967_11 (.CI(n49578), .I0(n1425), 
            .I1(VCC_net), .CO(n49579));
    SB_LUT4 encoder0_position_30__I_0_add_1503_4_lut (.I0(GND_net), .I1(n2232), 
            .I2(GND_net), .I3(n49852), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_5 (.CI(n49149), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n49150));
    SB_CARRY encoder0_position_30__I_0_add_1503_4 (.CI(n49852), .I0(n2232), 
            .I1(GND_net), .CO(n49853));
    SB_LUT4 encoder0_position_30__I_0_add_967_10_lut (.I0(GND_net), .I1(n1426), 
            .I2(VCC_net), .I3(n49577), .O(n1493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1503_3_lut (.I0(GND_net), .I1(n2233), 
            .I2(VCC_net), .I3(n49851), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_3 (.CI(n49851), .I0(n2233), 
            .I1(VCC_net), .CO(n49852));
    SB_LUT4 encoder0_position_30__I_0_add_1503_2_lut (.I0(GND_net), .I1(n947), 
            .I2(GND_net), .I3(VCC_net), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1503_2 (.CI(VCC_net), .I0(n947), 
            .I1(GND_net), .CO(n49851));
    SB_CARRY encoder0_position_30__I_0_add_967_10 (.CI(n49577), .I0(n1426), 
            .I1(VCC_net), .CO(n49578));
    SB_CARRY add_151_13 (.CI(n49157), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n49158));
    SB_LUT4 encoder0_position_30__I_0_add_1436_21_lut (.I0(n68812), .I1(n2115), 
            .I2(VCC_net), .I3(n49850), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_967_9_lut (.I0(GND_net), .I1(n1427), 
            .I2(VCC_net), .I3(n49576), .O(n1494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5860));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5859));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_1436_20_lut (.I0(GND_net), .I1(n2116), 
            .I2(VCC_net), .I3(n49849), .O(n2183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_20 (.CI(n49849), .I0(n2116), 
            .I1(VCC_net), .CO(n49850));
    SB_CARRY encoder0_position_30__I_0_add_967_9 (.CI(n49576), .I0(n1427), 
            .I1(VCC_net), .CO(n49577));
    SB_LUT4 encoder0_position_30__I_0_add_1436_19_lut (.I0(GND_net), .I1(n2117), 
            .I2(VCC_net), .I3(n49848), .O(n2184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_19 (.CI(n49848), .I0(n2117), 
            .I1(VCC_net), .CO(n49849));
    SB_LUT4 encoder0_position_30__I_0_add_1436_18_lut (.I0(GND_net), .I1(n2118), 
            .I2(VCC_net), .I3(n49847), .O(n2185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_18 (.CI(n49847), .I0(n2118), 
            .I1(VCC_net), .CO(n49848));
    SB_LUT4 encoder0_position_30__I_0_add_1436_17_lut (.I0(GND_net), .I1(n2119), 
            .I2(VCC_net), .I3(n49846), .O(n2186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_17 (.CI(n49846), .I0(n2119), 
            .I1(VCC_net), .CO(n49847));
    SB_LUT4 encoder0_position_30__I_0_add_1436_16_lut (.I0(GND_net), .I1(n2120), 
            .I2(VCC_net), .I3(n49845), .O(n2187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_16 (.CI(n49845), .I0(n2120), 
            .I1(VCC_net), .CO(n49846));
    SB_LUT4 encoder0_position_30__I_0_add_1436_15_lut (.I0(GND_net), .I1(n2121), 
            .I2(VCC_net), .I3(n49844), .O(n2188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_15 (.CI(n49844), .I0(n2121), 
            .I1(VCC_net), .CO(n49845));
    SB_LUT4 encoder0_position_30__I_0_add_1436_14_lut (.I0(GND_net), .I1(n2122), 
            .I2(VCC_net), .I3(n49843), .O(n2189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_14 (.CI(n49843), .I0(n2122), 
            .I1(VCC_net), .CO(n49844));
    SB_LUT4 encoder0_position_30__I_0_add_967_8_lut (.I0(GND_net), .I1(n1428), 
            .I2(VCC_net), .I3(n49575), .O(n1495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14), 
            .I3(n49413), .O(n299)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_8 (.CI(n49575), .I0(n1428), 
            .I1(VCC_net), .CO(n49576));
    SB_LUT4 encoder0_position_30__I_0_add_1436_13_lut (.I0(GND_net), .I1(n2123), 
            .I2(VCC_net), .I3(n49842), .O(n2190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5858));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i26_1_lut (.I0(encoder0_position[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5857));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i27_1_lut (.I0(encoder0_position[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5856));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1584_i13_3_lut (.I0(duty[15]), .I1(duty[12]), .I2(n260), 
            .I3(GND_net), .O(n12202));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i13_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY encoder0_position_30__I_0_add_1436_13 (.CI(n49842), .I0(n2123), 
            .I1(VCC_net), .CO(n49843));
    SB_LUT4 encoder0_position_30__I_0_add_1436_12_lut (.I0(GND_net), .I1(n2124), 
            .I2(VCC_net), .I3(n49841), .O(n2191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_12 (.CI(n49841), .I0(n2124), 
            .I1(VCC_net), .CO(n49842));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i28_1_lut (.I0(encoder0_position[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5855));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_967_7_lut (.I0(GND_net), .I1(n1429), 
            .I2(GND_net), .I3(n49574), .O(n1496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i29_1_lut (.I0(encoder0_position[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5854));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_967_7 (.CI(n49574), .I0(n1429), 
            .I1(GND_net), .CO(n49575));
    SB_CARRY unary_minus_16_add_3_13 (.CI(n49413), .I0(GND_net), .I1(n14), 
            .CO(n49414));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5670), 
            .I3(n49412), .O(n300)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_6_lut (.I0(GND_net), .I1(n1430), 
            .I2(GND_net), .I3(n49573), .O(n1497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n49412), .I0(GND_net), .I1(n15_adj_5670), 
            .CO(n49413));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i30_1_lut (.I0(encoder0_position[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5853));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_1584_i14_3_lut (.I0(duty[16]), .I1(duty[13]), .I2(n260), 
            .I3(GND_net), .O(n12200));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_add_1436_11_lut (.I0(GND_net), .I1(n2125), 
            .I2(VCC_net), .I3(n49840), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5671), 
            .I3(n49411), .O(n301)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i31_1_lut (.I0(encoder0_position[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5852));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n49411), .I0(GND_net), .I1(n16_adj_5671), 
            .CO(n49412));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_inv_0_i32_1_lut (.I0(encoder0_position[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5851));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[20]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_30__I_0_add_967_6 (.CI(n49573), .I0(n1430), 
            .I1(GND_net), .CO(n49574));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5672), 
            .I3(n49410), .O(n302)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_967_5_lut (.I0(GND_net), .I1(n1431), 
            .I2(VCC_net), .I3(n49572), .O(n1498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_967_5 (.CI(n49572), .I0(n1431), 
            .I1(VCC_net), .CO(n49573));
    SB_CARRY unary_minus_16_add_3_10 (.CI(n49410), .I0(GND_net), .I1(n17_adj_5672), 
            .CO(n49411));
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(current[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5672));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_967_4_lut (.I0(GND_net), .I1(n1432), 
            .I2(GND_net), .I3(n49571), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18), 
            .I3(n49409), .O(n303)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(current[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5671));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_967_4 (.CI(n49571), .I0(n1432), 
            .I1(GND_net), .CO(n49572));
    SB_LUT4 encoder0_position_30__I_0_add_967_3_lut (.I0(GND_net), .I1(n1433), 
            .I2(VCC_net), .I3(n49570), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n49409), .I0(GND_net), .I1(n18), 
            .CO(n49410));
    SB_CARRY encoder0_position_30__I_0_add_967_3 (.CI(n49570), .I0(n1433), 
            .I1(VCC_net), .CO(n49571));
    SB_LUT4 encoder0_position_30__I_0_add_967_2_lut (.I0(GND_net), .I1(n939), 
            .I2(GND_net), .I3(VCC_net), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_967_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_4310_i23_3_lut (.I0(encoder0_position[22]), .I1(n10_adj_5703), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n521));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i709_3_lut (.I0(n521), .I1(n1101), 
            .I2(n1059), .I3(GND_net), .O(n1133));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i776_3_lut (.I0(n1133), .I1(n1200), 
            .I2(n1158), .I3(GND_net), .O(n1232_adj_5800));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i843_3_lut (.I0(n1232_adj_5800), .I1(n1299), 
            .I2(n1257), .I3(GND_net), .O(n1331));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5673), 
            .I3(n49408), .O(n304)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i910_3_lut (.I0(n1331), .I1(n1398), 
            .I2(n1356), .I3(GND_net), .O(n1430));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i910_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_967_2 (.CI(VCC_net), .I0(n939), 
            .I1(GND_net), .CO(n49570));
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(current[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5670));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_4310_i24_3_lut (.I0(encoder0_position[23]), .I1(n9_adj_5704), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n520));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1436_11 (.CI(n49840), .I0(n2125), 
            .I1(VCC_net), .CO(n49841));
    SB_LUT4 encoder0_position_30__I_0_i641_3_lut (.I0(n520), .I1(n1001), 
            .I2(n960), .I3(GND_net), .O(n1033));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i708_3_lut (.I0(n1033), .I1(n1100), 
            .I2(n1059), .I3(GND_net), .O(n1132));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i775_3_lut (.I0(n1132), .I1(n1199), 
            .I2(n1158), .I3(GND_net), .O(n1231_adj_5799));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i775_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n49408), .I0(GND_net), .I1(n19_adj_5673), 
            .CO(n49409));
    SB_LUT4 encoder0_position_30__I_0_i842_3_lut (.I0(n1231_adj_5799), .I1(n1298), 
            .I2(n1257), .I3(GND_net), .O(n1330));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1436_10_lut (.I0(GND_net), .I1(n2126), 
            .I2(VCC_net), .I3(n49839), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i909_3_lut (.I0(n1330), .I1(n1397), 
            .I2(n1356), .I3(GND_net), .O(n1429));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i909_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1436_10 (.CI(n49839), .I0(n2126), 
            .I1(VCC_net), .CO(n49840));
    SB_LUT4 encoder0_position_30__I_0_add_1436_9_lut (.I0(GND_net), .I1(n2127), 
            .I2(VCC_net), .I3(n49838), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20_adj_5674), 
            .I3(n49407), .O(n305)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11579_bdd_4_lut_53711 (.I0(n11579), .I1(current[15]), .I2(duty[20]), 
            .I3(n11577), .O(n69444));
    defparam n11579_bdd_4_lut_53711.LUT_INIT = 16'he4aa;
    SB_CARRY encoder0_position_30__I_0_add_1436_9 (.CI(n49838), .I0(n2127), 
            .I1(VCC_net), .CO(n49839));
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n8_adj_5760), .I1(n3470), .I2(n161), 
            .I3(n10_adj_5683), .O(n28417));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n49407), .I0(GND_net), .I1(n20_adj_5674), 
            .CO(n49408));
    SB_LUT4 i1_2_lut_adj_1829 (.I0(n929), .I1(n930), .I2(GND_net), .I3(GND_net), 
            .O(n61300));
    defparam i1_2_lut_adj_1829.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21_adj_5675), 
            .I3(n49406), .O(n306)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n49156), .O(n1229)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1584_i15_3_lut (.I0(duty[17]), .I1(duty[14]), .I2(n260), 
            .I3(GND_net), .O(n12198));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i52764_1_lut (.I0(n3237), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68450));
    defparam i52764_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52756_1_lut (.I0(n43530), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68442));
    defparam i52756_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i2193_3_lut (.I0(n3222), .I1(n3289), 
            .I2(n3237), .I3(GND_net), .O(n27_adj_5888));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2193_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1830 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n56959));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i1_2_lut_adj_1830.LUT_INIT = 16'h2222;
    SB_LUT4 encoder0_position_30__I_0_i2198_3_lut (.I0(n3227), .I1(n3294), 
            .I2(n3237), .I3(GND_net), .O(n17_adj_5885));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2196_3_lut (.I0(n3225), .I1(n3292), 
            .I2(n3237), .I3(GND_net), .O(n21_adj_5887));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2197_3_lut (.I0(n3226), .I1(n3293), 
            .I2(n3237), .I3(GND_net), .O(n19_adj_5886));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1831 (.I0(n3224), .I1(n27_adj_5888), .I2(n3291), 
            .I3(n3237), .O(n61182));
    defparam i1_4_lut_adj_1831.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_i2190_3_lut (.I0(n3219), .I1(n3286), 
            .I2(n3237), .I3(GND_net), .O(n33));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2190_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1832 (.I0(n3229), .I1(n19_adj_5886), .I2(n3296), 
            .I3(n3237), .O(n61188));
    defparam i1_4_lut_adj_1832.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1833 (.I0(n3220), .I1(n21_adj_5887), .I2(n3287), 
            .I3(n3237), .O(n61180));
    defparam i1_4_lut_adj_1833.LUT_INIT = 16'heefc;
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY unary_minus_16_add_3_6 (.CI(n49406), .I0(GND_net), .I1(n21_adj_5675), 
            .CO(n49407));
    SB_LUT4 encoder0_position_30__I_0_add_1436_8_lut (.I0(GND_net), .I1(n2128), 
            .I2(VCC_net), .I3(n49837), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1834 (.I0(n61180), .I1(n61188), .I2(n33), .I3(n61182), 
            .O(n61196));
    defparam i1_4_lut_adj_1834.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n3231), .I1(n65401), .I2(n3237), .I3(n3230), 
            .O(n5_adj_5843));
    defparam i16_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 i50209_3_lut (.I0(n957), .I1(n3232), .I2(n3233), .I3(GND_net), 
            .O(n65411));
    defparam i50209_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22_adj_5676), 
            .I3(n49405), .O(n307)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_8 (.CI(n49837), .I0(n2128), 
            .I1(VCC_net), .CO(n49838));
    SB_CARRY unary_minus_16_add_3_5 (.CI(n49405), .I0(GND_net), .I1(n22_adj_5676), 
            .CO(n49406));
    SB_LUT4 i15764_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n60740), 
            .I3(n27_adj_5781), .O(n29772));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15764_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_add_1436_7_lut (.I0(GND_net), .I1(n2129), 
            .I2(GND_net), .I3(n49836), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5677), 
            .I3(n49404), .O(n308)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i2192_3_lut (.I0(n3221), .I1(n3288), 
            .I2(n3237), .I3(GND_net), .O(n29_adj_5889));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2192_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i52687_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n42632), .I3(GND_net), .O(n27698));
    defparam i52687_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_CARRY encoder0_position_30__I_0_add_1436_7 (.CI(n49836), .I0(n2129), 
            .I1(GND_net), .CO(n49837));
    SB_LUT4 encoder0_position_30__I_0_add_1436_6_lut (.I0(GND_net), .I1(n2130), 
            .I2(GND_net), .I3(n49835), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1835 (.I0(n3223), .I1(n17_adj_5885), .I2(n3290), 
            .I3(n3237), .O(n61186));
    defparam i1_4_lut_adj_1835.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1836 (.I0(n3228), .I1(n29_adj_5889), .I2(n3295), 
            .I3(n3237), .O(n61184));
    defparam i1_4_lut_adj_1836.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1837 (.I0(n65411), .I1(n5_adj_5843), .I2(n65412), 
            .I3(n3237), .O(n53307));
    defparam i1_4_lut_adj_1837.LUT_INIT = 16'h88c0;
    SB_LUT4 i1_4_lut_adj_1838 (.I0(n3218), .I1(n61196), .I2(n3285), .I3(n3237), 
            .O(n61200));
    defparam i1_4_lut_adj_1838.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1839 (.I0(n61200), .I1(n53307), .I2(n61184), 
            .I3(n61186), .O(n61202));
    defparam i1_4_lut_adj_1839.LUT_INIT = 16'hfffe;
    SB_LUT4 n69444_bdd_4_lut (.I0(n69444), .I1(duty[17]), .I2(n4911), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[17]));
    defparam n69444_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1840 (.I0(n3217), .I1(n61202), .I2(n3284), .I3(n3237), 
            .O(n61204));
    defparam i1_4_lut_adj_1840.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1841 (.I0(n3216), .I1(n61204), .I2(n3283), .I3(n3237), 
            .O(n61206));
    defparam i1_4_lut_adj_1841.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_30__I_0_add_1436_6 (.CI(n49835), .I0(n2130), 
            .I1(GND_net), .CO(n49836));
    SB_LUT4 i1_4_lut_adj_1842 (.I0(n3215), .I1(n61206), .I2(n3282), .I3(n3237), 
            .O(n61208));
    defparam i1_4_lut_adj_1842.LUT_INIT = 16'heefc;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n49404), .I0(GND_net), .I1(n23_adj_5677), 
            .CO(n49405));
    SB_LUT4 i1_4_lut_adj_1843 (.I0(n3214), .I1(n61208), .I2(n3281), .I3(n3237), 
            .O(n61210));
    defparam i1_4_lut_adj_1843.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_30__I_0_add_1436_5_lut (.I0(GND_net), .I1(n2131), 
            .I2(VCC_net), .I3(n49834), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_5 (.CI(n49834), .I0(n2131), 
            .I1(VCC_net), .CO(n49835));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5678), 
            .I3(n49403), .O(n309)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n49403), .I0(GND_net), .I1(n24_adj_5678), 
            .CO(n49404));
    SB_LUT4 encoder0_position_30__I_0_add_1436_4_lut (.I0(GND_net), .I1(n2132), 
            .I2(GND_net), .I3(n49833), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50087_2_lut_3_lut (.I0(n62), .I1(delay_counter[31]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n65309));
    defparam i50087_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_4_lut_adj_1844 (.I0(n3213), .I1(n61210), .I2(n3280), .I3(n3237), 
            .O(n61212));
    defparam i1_4_lut_adj_1844.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1845 (.I0(n3212), .I1(n61212), .I2(n3279), .I3(n3237), 
            .O(n61214));
    defparam i1_4_lut_adj_1845.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1846 (.I0(n3211), .I1(n61214), .I2(n3278), .I3(n3237), 
            .O(n61216));
    defparam i1_4_lut_adj_1846.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_30__I_0_add_1436_4 (.CI(n49833), .I0(n2132), 
            .I1(GND_net), .CO(n49834));
    SB_LUT4 encoder0_position_30__I_0_add_1436_3_lut (.I0(GND_net), .I1(n2133), 
            .I2(VCC_net), .I3(n49832), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16511_3_lut_4_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30519));   // verilog/coms.v(130[12] 305[6])
    defparam i16511_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_4_lut_adj_1847 (.I0(n3210), .I1(n61216), .I2(n3277), .I3(n3237), 
            .O(n61218));
    defparam i1_4_lut_adj_1847.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1848 (.I0(n3209), .I1(n61218), .I2(n3276), .I3(n3237), 
            .O(n61220));
    defparam i1_4_lut_adj_1848.LUT_INIT = 16'heefc;
    SB_LUT4 n11579_bdd_4_lut_53706 (.I0(n11579), .I1(current[15]), .I2(duty[19]), 
            .I3(n11577), .O(n69438));
    defparam n11579_bdd_4_lut_53706.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_4_lut_adj_1849 (.I0(n3208), .I1(n61220), .I2(n3275), .I3(n3237), 
            .O(n61222));
    defparam i1_4_lut_adj_1849.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1850 (.I0(n3207), .I1(n61222), .I2(n3274), .I3(n3237), 
            .O(n61224));
    defparam i1_4_lut_adj_1850.LUT_INIT = 16'heefc;
    SB_LUT4 i16510_3_lut_4_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30518));   // verilog/coms.v(130[12] 305[6])
    defparam i16510_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i2177_3_lut (.I0(n3206), .I1(n3273), 
            .I2(n3237), .I3(GND_net), .O(n59));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2176_3_lut (.I0(n3205), .I1(n3272), 
            .I2(n3237), .I3(GND_net), .O(n61));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15765_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n60788), 
            .I3(n27_adj_5781), .O(n29773));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15765_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_adj_1851 (.I0(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I1(Ki[1]), .I2(GND_net), .I3(GND_net), .O(n110));
    defparam i1_2_lut_adj_1851.LUT_INIT = 16'h8888;
    SB_LUT4 i28844_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n42632), .I3(GND_net), .O(n42746));
    defparam i28844_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i52759_4_lut (.I0(n61), .I1(n62365), .I2(n59), .I3(n61224), 
            .O(n43530));
    defparam i52759_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i16509_3_lut_4_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30517));   // verilog/coms.v(130[12] 305[6])
    defparam i16509_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mux_1584_i8_3_lut (.I0(duty[10]), .I1(duty[7]), .I2(n260), 
            .I3(GND_net), .O(n12212));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_i2110_3_lut (.I0(n3107), .I1(n3174), 
            .I2(n3138), .I3(GND_net), .O(n3206));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2109_3_lut (.I0(n3106), .I1(n3173), 
            .I2(n3138), .I3(GND_net), .O(n3205));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2113_3_lut (.I0(n3110), .I1(n3177), 
            .I2(n3138), .I3(GND_net), .O(n3209));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut_4_lut_4_lut (.I0(reset), .I1(n130), .I2(n8_adj_5731), 
            .I3(\FRAME_MATCHER.i [5]), .O(n28434));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 encoder0_position_30__I_0_i2112_3_lut (.I0(n3109), .I1(n3176), 
            .I2(n3138), .I3(GND_net), .O(n3208));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2111_3_lut (.I0(n3108), .I1(n3175), 
            .I2(n3138), .I3(GND_net), .O(n3207));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2116_3_lut (.I0(n3113), .I1(n3180), 
            .I2(n3138), .I3(GND_net), .O(n3212));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2115_3_lut (.I0(n3112), .I1(n3179), 
            .I2(n3138), .I3(GND_net), .O(n3211));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2114_3_lut (.I0(n3111), .I1(n3178), 
            .I2(n3138), .I3(GND_net), .O(n3210));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2120_3_lut (.I0(n3117), .I1(n3184), 
            .I2(n3138), .I3(GND_net), .O(n3216));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2119_3_lut (.I0(n3116), .I1(n3183), 
            .I2(n3138), .I3(GND_net), .O(n3215));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15766_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n60756), 
            .I3(n27_adj_5781), .O(n29774));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15766_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i2124_3_lut (.I0(n3121), .I1(n3188), 
            .I2(n3138), .I3(GND_net), .O(n3220));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n43349), .I1(GND_net), .I2(n25_adj_5679), 
            .I3(VCC_net), .O(n65285)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_i2122_3_lut (.I0(n3119), .I1(n3186), 
            .I2(n3138), .I3(GND_net), .O(n3218));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2118_3_lut (.I0(n3115), .I1(n3182), 
            .I2(n3138), .I3(GND_net), .O(n3214));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2117_3_lut (.I0(n3114), .I1(n3181), 
            .I2(n3138), .I3(GND_net), .O(n3213));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2129_3_lut (.I0(n3126), .I1(n3193), 
            .I2(n3138), .I3(GND_net), .O(n3225));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2123_3_lut (.I0(n3120), .I1(n3187), 
            .I2(n3138), .I3(GND_net), .O(n3219));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16507_3_lut_4_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30515));   // verilog/coms.v(130[12] 305[6])
    defparam i16507_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i2126_3_lut (.I0(n3123), .I1(n3190), 
            .I2(n3138), .I3(GND_net), .O(n3222));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2130_3_lut (.I0(n3127), .I1(n3194), 
            .I2(n3138), .I3(GND_net), .O(n3226));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2131_3_lut (.I0(n3128), .I1(n3195), 
            .I2(n3138), .I3(GND_net), .O(n3227));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2127_3_lut (.I0(n3124), .I1(n3191), 
            .I2(n3138), .I3(GND_net), .O(n3223));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2135_3_lut (.I0(n3132), .I1(n3199), 
            .I2(n3138), .I3(GND_net), .O(n3231));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2134_3_lut (.I0(n3131), .I1(n3198), 
            .I2(n3138), .I3(GND_net), .O(n3230));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2133_3_lut (.I0(n3130), .I1(n3197), 
            .I2(n3138), .I3(GND_net), .O(n3229));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16506_3_lut_4_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30514));   // verilog/coms.v(130[12] 305[6])
    defparam i16506_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i22434_3_lut (.I0(n219), .I1(IntegralLimit[12]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 [12]));
    defparam i22434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i2137_3_lut (.I0(n956), .I1(n3201), 
            .I2(n3138), .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2137_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1436_3 (.CI(n49832), .I0(n2133), 
            .I1(VCC_net), .CO(n49833));
    SB_LUT4 encoder0_position_30__I_0_add_1436_2_lut (.I0(GND_net), .I1(n946), 
            .I2(GND_net), .I3(VCC_net), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1436_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1436_2 (.CI(VCC_net), .I0(n946), 
            .I1(GND_net), .CO(n49832));
    SB_LUT4 i16505_3_lut_4_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30513));   // verilog/coms.v(130[12] 305[6])
    defparam i16505_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_5679), 
            .CO(n49403));
    SB_LUT4 i1_2_lut_adj_1852 (.I0(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I1(Ki[0]), .I2(GND_net), .I3(GND_net), .O(n38));
    defparam i1_2_lut_adj_1852.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_i2136_3_lut (.I0(n3133), .I1(n3200), 
            .I2(n3138), .I3(GND_net), .O(n3232));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(current[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53126_1_lut (.I0(n2148), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68812));
    defparam i53126_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_4310_i11_3_lut (.I0(encoder0_position[10]), .I1(n22_adj_5692), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n947));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_4310_i1_3_lut (.I0(encoder0_position[0]), .I1(n32), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n957));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i2128_3_lut (.I0(n3125), .I1(n3192), 
            .I2(n3138), .I3(GND_net), .O(n3224));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2132_3_lut (.I0(n3129), .I1(n3196), 
            .I2(n3138), .I3(GND_net), .O(n3228));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2_adj_5757), .I3(n49402), .O(displacement_23__N_67[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1853 (.I0(n927), .I1(n61300), .I2(n928), .I3(n43550), 
            .O(n960));
    defparam i1_4_lut_adj_1853.LUT_INIT = 16'hfefa;
    SB_LUT4 i16504_3_lut_4_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30512));   // verilog/coms.v(130[12] 305[6])
    defparam i16504_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i2125_3_lut (.I0(n3122), .I1(n3189), 
            .I2(n3138), .I3(GND_net), .O(n3221));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2121_3_lut (.I0(n3118), .I1(n3185), 
            .I2(n3138), .I3(GND_net), .O(n3217));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1854 (.I0(n3223), .I1(n3227), .I2(GND_net), .I3(GND_net), 
            .O(n61684));
    defparam i1_2_lut_adj_1854.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1855 (.I0(n3226), .I1(n3222), .I2(n3219), .I3(n3225), 
            .O(n61696));
    defparam i1_4_lut_adj_1855.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1584_i16_3_lut (.I0(duty[18]), .I1(duty[15]), .I2(n260), 
            .I3(GND_net), .O(n12196));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_5756), .I3(n49401), .O(displacement_23__N_67[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1856 (.I0(n3217), .I1(n3221), .I2(n3228), .I3(n3224), 
            .O(n61700));
    defparam i1_4_lut_adj_1856.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1857 (.I0(n3218), .I1(n61696), .I2(n61684), .I3(n3220), 
            .O(n61702));
    defparam i1_4_lut_adj_1857.LUT_INIT = 16'hfffe;
    SB_LUT4 i29615_3_lut (.I0(n957), .I1(n3232), .I2(n3233), .I3(GND_net), 
            .O(n43524));
    defparam i29615_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1858 (.I0(n3215), .I1(n61702), .I2(n3216), .I3(n61700), 
            .O(n61708));
    defparam i1_4_lut_adj_1858.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n49401), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_5756), .CO(n49402));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5755), .I3(n49400), .O(displacement_23__N_67[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1859 (.I0(n3229), .I1(n43524), .I2(n3230), .I3(n3231), 
            .O(n58789));
    defparam i1_4_lut_adj_1859.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1860 (.I0(n3213), .I1(n3214), .I2(n58789), .I3(n61708), 
            .O(n61714));
    defparam i1_4_lut_adj_1860.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1861 (.I0(n3210), .I1(n3211), .I2(n3212), .I3(n61714), 
            .O(n61720));
    defparam i1_4_lut_adj_1861.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1862 (.I0(n3207), .I1(n3208), .I2(n3209), .I3(n61720), 
            .O(n61726));
    defparam i1_4_lut_adj_1862.LUT_INIT = 16'hfffe;
    SB_LUT4 i52795_4_lut (.I0(n3205), .I1(n3204), .I2(n3206), .I3(n61726), 
            .O(n3237));
    defparam i52795_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i2043_3_lut (.I0(n3008), .I1(n3075), 
            .I2(n3039), .I3(GND_net), .O(n3107));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_4_lut (.I0(n62), .I1(delay_counter[31]), .I2(data_ready), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n6_adj_5900));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h2022;
    SB_LUT4 encoder0_position_30__I_0_i2042_3_lut (.I0(n3007), .I1(n3074), 
            .I2(n3039), .I3(GND_net), .O(n3106));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2042_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n49400), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5755), .CO(n49401));
    SB_LUT4 encoder0_position_30__I_0_i2046_3_lut (.I0(n3011), .I1(n3078), 
            .I2(n3039), .I3(GND_net), .O(n3110));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2045_3_lut (.I0(n3010), .I1(n3077), 
            .I2(n3039), .I3(GND_net), .O(n3109));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2044_3_lut (.I0(n3009), .I1(n3076), 
            .I2(n3039), .I3(GND_net), .O(n3108));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2051_3_lut (.I0(n3016), .I1(n3083), 
            .I2(n3039), .I3(GND_net), .O(n3115));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5785), .I3(n49399), .O(displacement_23__N_67[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i2050_3_lut (.I0(n3015), .I1(n3082), 
            .I2(n3039), .I3(GND_net), .O(n3114));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2049_3_lut (.I0(n3014), .I1(n3081), 
            .I2(n3039), .I3(GND_net), .O(n3113));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2049_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n49399), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5785), .CO(n49400));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5780), .I3(n49398), .O(displacement_23__N_67[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i2048_3_lut (.I0(n3013), .I1(n3080), 
            .I2(n3039), .I3(GND_net), .O(n3112));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2048_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n49398), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5780), .CO(n49399));
    SB_LUT4 encoder0_position_30__I_0_i2047_3_lut (.I0(n3012), .I1(n3079), 
            .I2(n3039), .I3(GND_net), .O(n3111));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2054_3_lut (.I0(n3019), .I1(n3086), 
            .I2(n3039), .I3(GND_net), .O(n3118));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2053_3_lut (.I0(n3018), .I1(n3085), 
            .I2(n3039), .I3(GND_net), .O(n3117));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2052_3_lut (.I0(n3017), .I1(n3084), 
            .I2(n3039), .I3(GND_net), .O(n3116));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2063_3_lut (.I0(n3028), .I1(n3095), 
            .I2(n3039), .I3(GND_net), .O(n3127));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2056_3_lut (.I0(n3021), .I1(n3088), 
            .I2(n3039), .I3(GND_net), .O(n3120));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2059_3_lut (.I0(n3024), .I1(n3091), 
            .I2(n3039), .I3(GND_net), .O(n3123));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2064_3_lut (.I0(n3029), .I1(n3096), 
            .I2(n3039), .I3(GND_net), .O(n3128));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2069_3_lut (.I0(n955), .I1(n3101), 
            .I2(n3039), .I3(GND_net), .O(n3133));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2069_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2068_3_lut (.I0(n3033), .I1(n3100), 
            .I2(n3039), .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2068_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[21]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_4310_i2_3_lut (.I0(encoder0_position[1]), .I1(n31), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n956));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i2067_3_lut (.I0(n3032), .I1(n3099), 
            .I2(n3039), .I3(GND_net), .O(n3131));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2067_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1855_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1319), .I3(n42632), .O(n6617));   // verilog/TinyFPGA_B.v(361[5] 387[12])
    defparam i1855_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5779), .I3(n49397), .O(displacement_23__N_67[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i2066_3_lut (.I0(n3031), .I1(n3098), 
            .I2(n3039), .I3(GND_net), .O(n3130));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2066_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2065_3_lut (.I0(n3030), .I1(n3097), 
            .I2(n3039), .I3(GND_net), .O(n3129));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1319), .I3(n42632), .O(n24_adj_5895));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 encoder0_position_30__I_0_add_900_13_lut (.I0(n69032), .I1(n1323), 
            .I2(VCC_net), .I3(n49548), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_i2062_3_lut (.I0(n3027), .I1(n3094), 
            .I2(n3039), .I3(GND_net), .O(n3126));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2055_3_lut (.I0(n3020), .I1(n3087), 
            .I2(n3039), .I3(GND_net), .O(n3119));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2061_3_lut (.I0(n3026), .I1(n3093), 
            .I2(n3039), .I3(GND_net), .O(n3125));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2061_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n49397), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5779), .CO(n49398));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5778), .I3(n49396), .O(displacement_23__N_67[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i2057_3_lut (.I0(n3022), .I1(n3089), 
            .I2(n3039), .I3(GND_net), .O(n3121));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i2058_3_lut (.I0(n3023), .I1(n3090), 
            .I2(n3039), .I3(GND_net), .O(n3122));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n69438_bdd_4_lut (.I0(n69438), .I1(duty[16]), .I2(n4912), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[16]));
    defparam n69438_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i2060_3_lut (.I0(n3025), .I1(n3092), 
            .I2(n3039), .I3(GND_net), .O(n3124));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i52826_1_lut (.I0(n3138), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68512));
    defparam i52826_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n49396), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5778), .CO(n49397));
    SB_LUT4 i29613_3_lut (.I0(n956), .I1(n3132), .I2(n3133), .I3(GND_net), 
            .O(n43522));
    defparam i29613_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1863 (.I0(n3128), .I1(n3123), .I2(n3120), .I3(n3127), 
            .O(n61030));
    defparam i1_4_lut_adj_1863.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5777), .I3(n49395), .O(displacement_23__N_67[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1864 (.I0(n3124), .I1(n3122), .I2(n3121), .I3(n3125), 
            .O(n61032));
    defparam i1_4_lut_adj_1864.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1865 (.I0(n61032), .I1(n61030), .I2(n3119), .I3(n3126), 
            .O(n61036));
    defparam i1_4_lut_adj_1865.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1866 (.I0(n3129), .I1(n43522), .I2(n3130), .I3(n3131), 
            .O(n58743));
    defparam i1_4_lut_adj_1866.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1867 (.I0(n3116), .I1(n3117), .I2(n61036), .I3(n3118), 
            .O(n61042));
    defparam i1_4_lut_adj_1867.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n49395), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5777), .CO(n49396));
    SB_LUT4 i1_4_lut_adj_1868 (.I0(n3114), .I1(n3115), .I2(n61042), .I3(n58743), 
            .O(n61048));
    defparam i1_4_lut_adj_1868.LUT_INIT = 16'hfffe;
    SB_LUT4 i50642_2_lut_3_lut (.I0(enable_slow_N_4211), .I1(ready_prev), 
            .I2(state_adj_5967[1]), .I3(GND_net), .O(n65486));   // verilog/eeprom.v(35[8] 81[4])
    defparam i50642_2_lut_3_lut.LUT_INIT = 16'hd0d0;
    SB_LUT4 i1_4_lut_adj_1869 (.I0(n3111), .I1(n3112), .I2(n3113), .I3(n61048), 
            .O(n61054));
    defparam i1_4_lut_adj_1869.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_900_12_lut (.I0(GND_net), .I1(n1324), 
            .I2(VCC_net), .I3(n49547), .O(n1391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1870 (.I0(n3108), .I1(n3109), .I2(n3110), .I3(n61054), 
            .O(n61060));
    defparam i1_4_lut_adj_1870.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_245_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[22]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(reset), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [2]), 
            .O(n56908));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_900_12 (.CI(n49547), .I0(n1324), 
            .I1(VCC_net), .CO(n49548));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1871 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [3]), 
            .O(n56907));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1871.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5776), .I3(n49394), .O(displacement_23__N_67[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52829_4_lut (.I0(n3106), .I1(n3105), .I2(n3107), .I3(n61060), 
            .O(n3138));
    defparam i52829_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1872 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [4]), 
            .O(n56906));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1872.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1976_3_lut (.I0(n2909), .I1(n2976), 
            .I2(n2940), .I3(GND_net), .O(n3008));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1974_3_lut (.I0(n2907), .I1(n2974), 
            .I2(n2940), .I3(GND_net), .O(n3006));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1975_3_lut (.I0(n2908), .I1(n2975), 
            .I2(n2940), .I3(GND_net), .O(n3007));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11579_bdd_4_lut_53701 (.I0(n11579), .I1(current[15]), .I2(duty[18]), 
            .I3(n11577), .O(n69432));
    defparam n11579_bdd_4_lut_53701.LUT_INIT = 16'he4aa;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n49394), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5776), .CO(n49395));
    SB_LUT4 encoder0_position_30__I_0_i1457_3_lut (.I0(n946), .I1(n2201), 
            .I2(n2148), .I3(GND_net), .O(n2233));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1457_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1456_3_lut (.I0(n2133), .I1(n2200), 
            .I2(n2148), .I3(GND_net), .O(n2232));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1873 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [5]), 
            .O(n56905));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1873.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1874 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [6]), 
            .O(n56952));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1874.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5775), .I3(n49393), .O(displacement_23__N_67[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1979_3_lut (.I0(n2912), .I1(n2979), 
            .I2(n2940), .I3(GND_net), .O(n3011));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1875 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [7]), 
            .O(n56904));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1875.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1876 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [0]), 
            .O(n56773));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1876.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1978_3_lut (.I0(n2911), .I1(n2978), 
            .I2(n2940), .I3(GND_net), .O(n3010));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1877 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [1]), 
            .O(n56903));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1877.LUT_INIT = 16'h2300;
    SB_LUT4 i12_3_lut_4_lut (.I0(rx_data_ready), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n27724), .O(n52851));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 encoder0_position_30__I_0_i1977_3_lut (.I0(n2910), .I1(n2977), 
            .I2(n2940), .I3(GND_net), .O(n3009));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_900_11_lut (.I0(GND_net), .I1(n1325), 
            .I2(VCC_net), .I3(n49546), .O(n1392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_11 (.CI(n49546), .I0(n1325), 
            .I1(VCC_net), .CO(n49547));
    SB_LUT4 encoder0_position_30__I_0_add_900_10_lut (.I0(GND_net), .I1(n1326), 
            .I2(VCC_net), .I3(n49545), .O(n1393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1878 (.I0(control_mode[3]), .I1(control_mode[4]), 
            .I2(control_mode[6]), .I3(control_mode[2]), .O(n61854));   // verilog/TinyFPGA_B.v(287[5:22])
    defparam i1_4_lut_adj_1878.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_add_900_10 (.CI(n49545), .I0(n1326), 
            .I1(VCC_net), .CO(n49546));
    SB_LUT4 encoder0_position_30__I_0_add_900_9_lut (.I0(GND_net), .I1(n1327), 
            .I2(VCC_net), .I3(n49544), .O(n1394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_9 (.CI(n49544), .I0(n1327), 
            .I1(VCC_net), .CO(n49545));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n49393), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5775), .CO(n49394));
    SB_LUT4 add_151_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n49177), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1879 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [2]), 
            .O(n56902));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1879.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_900_8_lut (.I0(GND_net), .I1(n1328), 
            .I2(VCC_net), .I3(n49543), .O(n1395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5764), .I3(n49392), .O(displacement_23__N_67[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n49176), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_8 (.CI(n49543), .I0(n1328), 
            .I1(VCC_net), .CO(n49544));
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_151_32 (.CI(n49176), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n49177));
    SB_LUT4 encoder0_position_30__I_0_add_900_7_lut (.I0(GND_net), .I1(n1329), 
            .I2(GND_net), .I3(n49542), .O(n1396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1369_20_lut (.I0(n68808), .I1(n2016), 
            .I2(VCC_net), .I3(n49809), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 n69432_bdd_4_lut (.I0(n69432), .I1(duty[15]), .I2(n4913), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[15]));
    defparam n69432_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11579_bdd_4_lut_53696 (.I0(n11579), .I1(current[15]), .I2(duty[17]), 
            .I3(n11577), .O(n69426));
    defparam n11579_bdd_4_lut_53696.LUT_INIT = 16'he4aa;
    SB_LUT4 n69426_bdd_4_lut (.I0(n69426), .I1(duty[14]), .I2(n4914), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[14]));
    defparam n69426_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11579_bdd_4_lut_53691 (.I0(n11579), .I1(current[15]), .I2(duty[16]), 
            .I3(n11577), .O(n69420));
    defparam n11579_bdd_4_lut_53691.LUT_INIT = 16'he4aa;
    SB_LUT4 n69420_bdd_4_lut (.I0(n69420), .I1(duty[13]), .I2(n4915), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[13]));
    defparam n69420_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11579_bdd_4_lut_53686 (.I0(n11579), .I1(current[15]), .I2(duty[15]), 
            .I3(n11577), .O(n69414));
    defparam n11579_bdd_4_lut_53686.LUT_INIT = 16'he4aa;
    SB_LUT4 n69414_bdd_4_lut (.I0(n69414), .I1(duty[12]), .I2(n4916), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[12]));
    defparam n69414_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11579_bdd_4_lut_53681 (.I0(n11579), .I1(current[11]), .I2(duty[14]), 
            .I3(n11577), .O(n69408));
    defparam n11579_bdd_4_lut_53681.LUT_INIT = 16'he4aa;
    SB_LUT4 n69408_bdd_4_lut (.I0(n69408), .I1(duty[11]), .I2(n4917), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[11]));
    defparam n69408_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11579_bdd_4_lut_53676 (.I0(n11579), .I1(current[10]), .I2(duty[13]), 
            .I3(n11577), .O(n69402));
    defparam n11579_bdd_4_lut_53676.LUT_INIT = 16'he4aa;
    SB_LUT4 n69402_bdd_4_lut (.I0(n69402), .I1(duty[10]), .I2(n4918), 
            .I3(n11577), .O(pwm_setpoint_23__N_3[10]));
    defparam n69402_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11579_bdd_4_lut_53671 (.I0(n11579), .I1(current[9]), .I2(duty[12]), 
            .I3(n11577), .O(n69396));
    defparam n11579_bdd_4_lut_53671.LUT_INIT = 16'he4aa;
    SB_LUT4 n69396_bdd_4_lut (.I0(n69396), .I1(duty[9]), .I2(n4919), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[9]));
    defparam n69396_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n11579_bdd_4_lut_53666 (.I0(n11579), .I1(current[8]), .I2(duty[11]), 
            .I3(n11577), .O(n69390));
    defparam n11579_bdd_4_lut_53666.LUT_INIT = 16'he4aa;
    SB_LUT4 n69390_bdd_4_lut (.I0(n69390), .I1(duty[8]), .I2(n4920), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[8]));
    defparam n69390_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1880 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [3]), 
            .O(n56901));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1880.LUT_INIT = 16'h2300;
    SB_LUT4 n11579_bdd_4_lut_53661 (.I0(n11579), .I1(current[7]), .I2(duty[10]), 
            .I3(n11577), .O(n69384));
    defparam n11579_bdd_4_lut_53661.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_3_lut_adj_1881 (.I0(n61854), .I1(control_mode[5]), .I2(control_mode[7]), 
            .I3(GND_net), .O(n25507));   // verilog/TinyFPGA_B.v(287[5:22])
    defparam i1_3_lut_adj_1881.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_30__I_0_add_900_7 (.CI(n49542), .I0(n1329), 
            .I1(GND_net), .CO(n49543));
    SB_LUT4 encoder0_position_30__I_0_add_1369_19_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n49808), .O(n2084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_19 (.CI(n49808), .I0(n2017), 
            .I1(VCC_net), .CO(n49809));
    SB_LUT4 encoder0_position_30__I_0_i1983_3_lut (.I0(n2916), .I1(n2983), 
            .I2(n2940), .I3(GND_net), .O(n3015));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1369_18_lut (.I0(GND_net), .I1(n2018), 
            .I2(VCC_net), .I3(n49807), .O(n2085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_18 (.CI(n49807), .I0(n2018), 
            .I1(VCC_net), .CO(n49808));
    SB_LUT4 encoder0_position_30__I_0_add_900_6_lut (.I0(GND_net), .I1(n1330), 
            .I2(GND_net), .I3(n49541), .O(n1397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1369_17_lut (.I0(GND_net), .I1(n2019), 
            .I2(VCC_net), .I3(n49806), .O(n2086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_6 (.CI(n49541), .I0(n1330), 
            .I1(GND_net), .CO(n49542));
    SB_LUT4 encoder0_position_30__I_0_i1982_3_lut (.I0(n2915), .I1(n2982), 
            .I2(n2940), .I3(GND_net), .O(n3014));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_900_5_lut (.I0(GND_net), .I1(n1331), 
            .I2(VCC_net), .I3(n49540), .O(n1398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1882 (.I0(n25398), .I1(control_mode[1]), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(287[5:22])
    defparam i1_2_lut_adj_1882.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_3_lut_adj_1883 (.I0(control_mode[0]), .I1(n25507), .I2(control_mode[1]), 
            .I3(GND_net), .O(n15_adj_5681));   // verilog/TinyFPGA_B.v(286[5:22])
    defparam i1_3_lut_adj_1883.LUT_INIT = 16'hfdfd;
    SB_LUT4 mux_245_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[23]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_30__I_0_add_1369_17 (.CI(n49806), .I0(n2019), 
            .I1(VCC_net), .CO(n49807));
    SB_LUT4 encoder0_position_30__I_0_i1981_3_lut (.I0(n2914), .I1(n2981), 
            .I2(n2940), .I3(GND_net), .O(n3013));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1981_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_900_5 (.CI(n49540), .I0(n1331), 
            .I1(VCC_net), .CO(n49541));
    SB_LUT4 encoder0_position_30__I_0_i1980_3_lut (.I0(n2913), .I1(n2980), 
            .I2(n2940), .I3(GND_net), .O(n3012));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1369_16_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n49805), .O(n2087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1884 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [4]), 
            .O(n56900));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1884.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_900_4_lut (.I0(GND_net), .I1(n1332), 
            .I2(GND_net), .I3(n49539), .O(n1399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_16 (.CI(n49805), .I0(n2020), 
            .I1(VCC_net), .CO(n49806));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n49392), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5764), .CO(n49393));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5763), .I3(n49391), .O(displacement_23__N_67[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_4 (.CI(n49539), .I0(n1332), 
            .I1(GND_net), .CO(n49540));
    SB_LUT4 encoder0_position_30__I_0_add_1369_15_lut (.I0(GND_net), .I1(n2021), 
            .I2(VCC_net), .I3(n49804), .O(n2088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n49391), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5763), .CO(n49392));
    SB_LUT4 encoder0_position_30__I_0_i1998_3_lut (.I0(n2931), .I1(n2998), 
            .I2(n2940), .I3(GND_net), .O(n3030));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1998_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1369_15 (.CI(n49804), .I0(n2021), 
            .I1(VCC_net), .CO(n49805));
    SB_LUT4 encoder0_position_30__I_0_add_900_3_lut (.I0(GND_net), .I1(n1333), 
            .I2(VCC_net), .I3(n49538), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1997_3_lut (.I0(n2930), .I1(n2997), 
            .I2(n2940), .I3(GND_net), .O(n3029));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1369_14_lut (.I0(GND_net), .I1(n2022), 
            .I2(VCC_net), .I3(n49803), .O(n2089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i2001_3_lut (.I0(n954), .I1(n3001), 
            .I2(n2940), .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2001_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_900_3 (.CI(n49538), .I0(n1333), 
            .I1(VCC_net), .CO(n49539));
    SB_LUT4 encoder0_position_30__I_0_add_900_2_lut (.I0(GND_net), .I1(n524), 
            .I2(GND_net), .I3(VCC_net), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_900_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_14 (.CI(n49803), .I0(n2022), 
            .I1(VCC_net), .CO(n49804));
    SB_LUT4 encoder0_position_30__I_0_add_1369_13_lut (.I0(GND_net), .I1(n2023), 
            .I2(VCC_net), .I3(n49802), .O(n2090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_13 (.CI(n49802), .I0(n2023), 
            .I1(VCC_net), .CO(n49803));
    SB_LUT4 encoder0_position_30__I_0_add_1369_12_lut (.I0(GND_net), .I1(n2024), 
            .I2(VCC_net), .I3(n49801), .O(n2091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_12 (.CI(n49801), .I0(n2024), 
            .I1(VCC_net), .CO(n49802));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14_adj_5762), .I3(n49390), .O(displacement_23__N_67[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_900_2 (.CI(VCC_net), .I0(n524), 
            .I1(GND_net), .CO(n49538));
    SB_LUT4 encoder0_position_30__I_0_add_1369_11_lut (.I0(GND_net), .I1(n2025), 
            .I2(VCC_net), .I3(n49800), .O(n2092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_11 (.CI(n49800), .I0(n2025), 
            .I1(VCC_net), .CO(n49801));
    SB_LUT4 encoder0_position_30__I_0_add_1369_10_lut (.I0(GND_net), .I1(n2026), 
            .I2(VCC_net), .I3(n49799), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_10 (.CI(n49799), .I0(n2026), 
            .I1(VCC_net), .CO(n49800));
    SB_LUT4 encoder0_position_30__I_0_add_1369_9_lut (.I0(GND_net), .I1(n2027), 
            .I2(VCC_net), .I3(n49798), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_9 (.CI(n49798), .I0(n2027), 
            .I1(VCC_net), .CO(n49799));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n49390), .I0(encoder0_position_scaled[11]), 
            .I1(n14_adj_5762), .CO(n49391));
    SB_LUT4 encoder0_position_30__I_0_add_1369_8_lut (.I0(GND_net), .I1(n2028), 
            .I2(VCC_net), .I3(n49797), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1885 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [5]), 
            .O(n56899));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1885.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i2000_3_lut (.I0(n2933), .I1(n3000), 
            .I2(n2940), .I3(GND_net), .O(n3032));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i2000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5761), .I3(n49389), .O(displacement_23__N_67[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_8 (.CI(n49797), .I0(n2028), 
            .I1(VCC_net), .CO(n49798));
    SB_LUT4 encoder0_position_30__I_0_add_1369_7_lut (.I0(GND_net), .I1(n2029), 
            .I2(GND_net), .I3(n49796), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1999_3_lut (.I0(n2932), .I1(n2999), 
            .I2(n2940), .I3(GND_net), .O(n3031));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1886 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [6]), 
            .O(n56898));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1886.LUT_INIT = 16'h2300;
    SB_LUT4 mux_4310_i3_3_lut (.I0(encoder0_position[2]), .I1(n30), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n955));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_30__I_0_add_1369_7 (.CI(n49796), .I0(n2029), 
            .I1(GND_net), .CO(n49797));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n49389), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5761), .CO(n49390));
    SB_LUT4 encoder0_position_30__I_0_add_1369_6_lut (.I0(GND_net), .I1(n2030), 
            .I2(GND_net), .I3(n49795), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1989_3_lut (.I0(n2922), .I1(n2989), 
            .I2(n2940), .I3(GND_net), .O(n3021));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1989_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1369_6 (.CI(n49795), .I0(n2030), 
            .I1(GND_net), .CO(n49796));
    SB_LUT4 add_151_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n49175), .O(n1210)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1369_5_lut (.I0(GND_net), .I1(n2031), 
            .I2(VCC_net), .I3(n49794), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1995_3_lut (.I0(n2928), .I1(n2995), 
            .I2(n2940), .I3(GND_net), .O(n3027));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16_4_lut_4_lut (.I0(state_adj_5997[0]), .I1(n65481), .I2(n6428), 
            .I3(n10_adj_5729), .O(n8_adj_5911));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut_4_lut.LUT_INIT = 16'h3a7a;
    SB_LUT4 encoder0_position_30__I_0_i1991_3_lut (.I0(n2924), .I1(n2991), 
            .I2(n2940), .I3(GND_net), .O(n3023));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1991_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1369_5 (.CI(n49794), .I0(n2031), 
            .I1(VCC_net), .CO(n49795));
    SB_LUT4 encoder0_position_30__I_0_i1993_3_lut (.I0(n2926), .I1(n2993), 
            .I2(n2940), .I3(GND_net), .O(n3025));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1887 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [7]), 
            .O(n56897));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1887.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1985_3_lut (.I0(n2918), .I1(n2985), 
            .I2(n2940), .I3(GND_net), .O(n3017));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1985_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1888 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [0]), 
            .O(n56896));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1888.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1984_3_lut (.I0(n2917), .I1(n2984), 
            .I2(n2940), .I3(GND_net), .O(n3016));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1889 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [1]), 
            .O(n56895));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1889.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1890 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [2]), 
            .O(n56894));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1890.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1988_3_lut (.I0(n2921), .I1(n2988), 
            .I2(n2940), .I3(GND_net), .O(n3020));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1988_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1891 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [3]), 
            .O(n56893));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1891.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1369_4_lut (.I0(GND_net), .I1(n2032), 
            .I2(GND_net), .I3(n49793), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_4 (.CI(n49793), .I0(n2032), 
            .I1(GND_net), .CO(n49794));
    SB_LUT4 encoder0_position_30__I_0_add_1369_3_lut (.I0(GND_net), .I1(n2033), 
            .I2(VCC_net), .I3(n49792), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_3 (.CI(n49792), .I0(n2033), 
            .I1(VCC_net), .CO(n49793));
    SB_LUT4 encoder0_position_30__I_0_add_1369_2_lut (.I0(GND_net), .I1(n945), 
            .I2(GND_net), .I3(VCC_net), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1369_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5759), .I3(n49388), .O(displacement_23__N_67[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1369_2 (.CI(VCC_net), .I0(n945), 
            .I1(GND_net), .CO(n49792));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1892 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [4]), 
            .O(n56892));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1892.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1986_3_lut (.I0(n2919), .I1(n2986), 
            .I2(n2940), .I3(GND_net), .O(n3018));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1986_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_151_31 (.CI(n49175), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n49176));
    SB_LUT4 n69384_bdd_4_lut (.I0(n69384), .I1(duty[7]), .I2(n4921), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[7]));
    defparam n69384_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1893 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [5]), 
            .O(n56891));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1893.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1894 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [6]), 
            .O(n56890));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1894.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1895 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [7]), 
            .O(n56889));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1895.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1455_3_lut (.I0(n2132), .I1(n2199), 
            .I2(n2148), .I3(GND_net), .O(n2231));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1896 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [0]), 
            .O(n56888));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1896.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1990_3_lut (.I0(n2923), .I1(n2990), 
            .I2(n2940), .I3(GND_net), .O(n3022));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1990_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n49388), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5759), .CO(n49389));
    SB_CARRY add_151_12 (.CI(n49156), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n49157));
    SB_LUT4 add_151_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n49174), .O(n1211)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1996_3_lut (.I0(n2929), .I1(n2996), 
            .I2(n2940), .I3(GND_net), .O(n3028));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1897 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [1]), 
            .O(n56887));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1897.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5754), .I3(n49387), .O(displacement_23__N_67[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1987_3_lut (.I0(n2920), .I1(n2987), 
            .I2(n2940), .I3(GND_net), .O(n3019));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1992_3_lut (.I0(n2925), .I1(n2992), 
            .I2(n2940), .I3(GND_net), .O(n3024));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1994_3_lut (.I0(n2927), .I1(n2994), 
            .I2(n2940), .I3(GND_net), .O(n3026));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1994_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n49387), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5754), .CO(n49388));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18_adj_5753), .I3(n49386), .O(displacement_23__N_67[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n49386), .I0(encoder0_position_scaled[7]), 
            .I1(n18_adj_5753), .CO(n49387));
    SB_LUT4 add_151_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n49148), .O(n1237)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19_adj_5752), .I3(n49385), .O(displacement_23__N_67[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n49385), .I0(encoder0_position_scaled[6]), 
            .I1(n19_adj_5752), .CO(n49386));
    SB_CARRY add_151_30 (.CI(n49174), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n49175));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20), .I3(n49384), .O(displacement_23__N_67[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n49384), .I0(encoder0_position_scaled[5]), 
            .I1(n20), .CO(n49385));
    SB_LUT4 i52865_1_lut (.I0(n3039), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68551));
    defparam i52865_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1898 (.I0(n3025), .I1(n3023), .I2(n3027), .I3(n3021), 
            .O(n61598));
    defparam i1_4_lut_adj_1898.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1899 (.I0(n3026), .I1(n3024), .I2(n3019), .I3(n3028), 
            .O(n61596));
    defparam i1_4_lut_adj_1899.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1900 (.I0(n61598), .I1(n3022), .I2(n3018), .I3(n3020), 
            .O(n61600));
    defparam i1_4_lut_adj_1900.LUT_INIT = 16'hfffe;
    SB_LUT4 n11579_bdd_4_lut_53656 (.I0(n11579), .I1(current[6]), .I2(duty[9]), 
            .I3(n11577), .O(n69378));
    defparam n11579_bdd_4_lut_53656.LUT_INIT = 16'he4aa;
    SB_LUT4 i29661_4_lut (.I0(n955), .I1(n3031), .I2(n3032), .I3(n3033), 
            .O(n43570));
    defparam i29661_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21), .I3(n49383), .O(displacement_23__N_67[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n49155), .O(n1230)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1901 (.I0(n3016), .I1(n61600), .I2(n3017), .I3(n61596), 
            .O(n61606));
    defparam i1_4_lut_adj_1901.LUT_INIT = 16'hfffe;
    SB_LUT4 n69378_bdd_4_lut (.I0(n69378), .I1(duty[6]), .I2(n4922), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[6]));
    defparam n69378_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n49383), .I0(encoder0_position_scaled[4]), 
            .I1(n21), .CO(n49384));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22), .I3(n49382), .O(displacement_23__N_67[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1902 (.I0(n3029), .I1(n3030), .I2(GND_net), .I3(GND_net), 
            .O(n61740));
    defparam i1_2_lut_adj_1902.LUT_INIT = 16'h8888;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n49382), .I0(encoder0_position_scaled[3]), 
            .I1(n22), .CO(n49383));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23), .I3(n49381), .O(displacement_23__N_67[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n49381), .I0(encoder0_position_scaled[2]), 
            .I1(n23), .CO(n49382));
    SB_LUT4 i1_4_lut_adj_1903 (.I0(n3015), .I1(n61740), .I2(n61606), .I3(n43570), 
            .O(n61610));
    defparam i1_4_lut_adj_1903.LUT_INIT = 16'hfefa;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24), .I3(n49380), .O(displacement_23__N_67[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1904 (.I0(n3012), .I1(n3013), .I2(n3014), .I3(n61610), 
            .O(n61616));
    defparam i1_4_lut_adj_1904.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1905 (.I0(n3009), .I1(n3010), .I2(n3011), .I3(n61616), 
            .O(n61622));
    defparam i1_4_lut_adj_1905.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n49380), .I0(encoder0_position_scaled[1]), 
            .I1(n24), .CO(n49381));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder0_position_scaled[0]), 
            .I2(n25), .I3(VCC_net), .O(displacement_23__N_67[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52868_4_lut (.I0(n3007), .I1(n3006), .I2(n3008), .I3(n61622), 
            .O(n3039));
    defparam i52868_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 add_1097_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_207), 
            .I3(n49286), .O(n4905)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1097_24_lut (.I0(GND_net), .I1(GND_net), .I2(n12182), 
            .I3(n49285), .O(n4906)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1908_3_lut (.I0(n2809), .I1(n2876), 
            .I2(n2841), .I3(GND_net), .O(n2908));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1908_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1097_24 (.CI(n49285), .I0(GND_net), .I1(n12182), .CO(n49286));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1906 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [2]), 
            .O(n56886));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1906.LUT_INIT = 16'h2300;
    SB_LUT4 mux_1584_i17_3_lut (.I0(duty[19]), .I1(duty[16]), .I2(n260), 
            .I3(GND_net), .O(n12194));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_i1914_3_lut (.I0(n2815), .I1(n2882), 
            .I2(n2841), .I3(GND_net), .O(n2914));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1914_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder0_position_scaled[0]), 
            .I1(n25), .CO(n49380));
    SB_LUT4 encoder0_position_30__I_0_add_833_12_lut (.I0(n69005), .I1(n1224_adj_5792), 
            .I2(VCC_net), .I3(n49523), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_1097_23_lut (.I0(GND_net), .I1(GND_net), .I2(n12184), 
            .I3(n49284), .O(n4907)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1097_23 (.CI(n49284), .I0(GND_net), .I1(n12184), .CO(n49285));
    SB_LUT4 encoder0_position_30__I_0_add_833_11_lut (.I0(GND_net), .I1(n1225_adj_5793), 
            .I2(VCC_net), .I3(n49522), .O(n1292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_11 (.CI(n49522), .I0(n1225_adj_5793), 
            .I1(VCC_net), .CO(n49523));
    SB_LUT4 encoder0_position_30__I_0_i1910_3_lut (.I0(n2811), .I1(n2878), 
            .I2(n2841), .I3(GND_net), .O(n2910));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_833_10_lut (.I0(GND_net), .I1(n1226_adj_5794), 
            .I2(VCC_net), .I3(n49521), .O(n1293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1912_3_lut (.I0(n2813), .I1(n2880), 
            .I2(n2841), .I3(GND_net), .O(n2912));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1912_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_833_10 (.CI(n49521), .I0(n1226_adj_5794), 
            .I1(VCC_net), .CO(n49522));
    SB_LUT4 encoder0_position_30__I_0_add_833_9_lut (.I0(GND_net), .I1(n1227_adj_5795), 
            .I2(VCC_net), .I3(n49520), .O(n1294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_9 (.CI(n49520), .I0(n1227_adj_5795), 
            .I1(VCC_net), .CO(n49521));
    SB_LUT4 encoder0_position_30__I_0_add_833_8_lut (.I0(GND_net), .I1(n1228_adj_5796), 
            .I2(VCC_net), .I3(n49519), .O(n1295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_8 (.CI(n49519), .I0(n1228_adj_5796), 
            .I1(VCC_net), .CO(n49520));
    SB_LUT4 add_1097_22_lut (.I0(GND_net), .I1(GND_net), .I2(n12186), 
            .I3(n49283), .O(n4908)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1097_22 (.CI(n49283), .I0(GND_net), .I1(n12186), .CO(n49284));
    SB_LUT4 add_1097_21_lut (.I0(GND_net), .I1(GND_net), .I2(n12188), 
            .I3(n49282), .O(n4909)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_833_7_lut (.I0(GND_net), .I1(n1229_adj_5797), 
            .I2(GND_net), .I3(n49518), .O(n1296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n49173), .O(n1212)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_7 (.CI(n49518), .I0(n1229_adj_5797), 
            .I1(GND_net), .CO(n49519));
    SB_LUT4 encoder0_position_30__I_0_i1930_3_lut (.I0(n2831), .I1(n2898), 
            .I2(n2841), .I3(GND_net), .O(n2930));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1929_3_lut (.I0(n2830), .I1(n2897), 
            .I2(n2841), .I3(GND_net), .O(n2929));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i42184_3_lut (.I0(n4_adj_5714), .I1(n7452), .I2(n57811), .I3(GND_net), 
            .O(n57814));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42185_3_lut (.I0(encoder0_position[28]), .I1(n57814), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n830));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i569_3_lut (.I0(n830), .I1(n897), 
            .I2(n861), .I3(GND_net), .O(n929));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i636_3_lut (.I0(n929), .I1(n996), 
            .I2(n960), .I3(GND_net), .O(n1028));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i703_3_lut (.I0(n1028), .I1(n1095), 
            .I2(n1059), .I3(GND_net), .O(n1127));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i770_3_lut (.I0(n1127), .I1(n1194), 
            .I2(n1158), .I3(GND_net), .O(n1226_adj_5794));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i770_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i837_3_lut (.I0(n1226_adj_5794), .I1(n1293), 
            .I2(n1257), .I3(GND_net), .O(n1325));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i904_3_lut (.I0(n1325), .I1(n1392), 
            .I2(n1356), .I3(GND_net), .O(n1424));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i904_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1907 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [3]), 
            .O(n56885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1907.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1908 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [4]), 
            .O(n56884));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1908.LUT_INIT = 16'h2300;
    SB_LUT4 i16462_3_lut_4_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30470));   // verilog/coms.v(130[12] 305[6])
    defparam i16462_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1920_3_lut (.I0(n2821), .I1(n2888), 
            .I2(n2841), .I3(GND_net), .O(n2920));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1920_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1097_21 (.CI(n49282), .I0(GND_net), .I1(n12188), .CO(n49283));
    SB_LUT4 encoder0_position_30__I_0_add_833_6_lut (.I0(GND_net), .I1(n1230_adj_5798), 
            .I2(GND_net), .I3(n49517), .O(n1297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1926_3_lut (.I0(n2827), .I1(n2894), 
            .I2(n2841), .I3(GND_net), .O(n2926));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1097_20_lut (.I0(GND_net), .I1(GND_net), .I2(n12190), 
            .I3(n49281), .O(n4910)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_11 (.CI(n49155), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n49156));
    SB_LUT4 encoder0_position_30__I_0_i1919_3_lut (.I0(n2820_adj_5813), .I1(n2887), 
            .I2(n2841), .I3(GND_net), .O(n2919));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1922_3_lut (.I0(n2823), .I1(n2890), 
            .I2(n2841), .I3(GND_net), .O(n2922));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1922_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_833_6 (.CI(n49517), .I0(n1230_adj_5798), 
            .I1(GND_net), .CO(n49518));
    SB_LUT4 encoder0_position_30__I_0_add_833_5_lut (.I0(GND_net), .I1(n1231_adj_5799), 
            .I2(VCC_net), .I3(n49516), .O(n1298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1909 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [5]), 
            .O(n56883));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1909.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1454_3_lut (.I0(n2131), .I1(n2198), 
            .I2(n2148), .I3(GND_net), .O(n2230));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1928_3_lut (.I0(n2829), .I1(n2896), 
            .I2(n2841), .I3(GND_net), .O(n2928));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1928_3_lut.LUT_INIT = 16'hacac;
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i16460_3_lut_4_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30468));   // verilog/coms.v(130[12] 305[6])
    defparam i16460_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1924_3_lut (.I0(n2825), .I1(n2892), 
            .I2(n2841), .I3(GND_net), .O(n2924));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1921_3_lut (.I0(n2822), .I1(n2889), 
            .I2(n2841), .I3(GND_net), .O(n2921));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1584_i18_3_lut (.I0(duty[20]), .I1(duty[17]), .I2(n260), 
            .I3(GND_net), .O(n12192));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_i1925_3_lut (.I0(n2826), .I1(n2893), 
            .I2(n2841), .I3(GND_net), .O(n2925));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1453_3_lut (.I0(n2130), .I1(n2197), 
            .I2(n2148), .I3(GND_net), .O(n2229));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1453_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1097_20 (.CI(n49281), .I0(GND_net), .I1(n12190), .CO(n49282));
    SB_LUT4 encoder0_position_30__I_0_i1916_3_lut (.I0(n2817), .I1(n2884), 
            .I2(n2841), .I3(GND_net), .O(n2916));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1916_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_833_5 (.CI(n49516), .I0(n1231_adj_5799), 
            .I1(VCC_net), .CO(n49517));
    SB_LUT4 encoder0_position_30__I_0_add_833_4_lut (.I0(GND_net), .I1(n1232_adj_5800), 
            .I2(GND_net), .I3(n49515), .O(n1299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1452_3_lut (.I0(n2129), .I1(n2196), 
            .I2(n2148), .I3(GND_net), .O(n2228));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1915_3_lut (.I0(n2816), .I1(n2883), 
            .I2(n2841), .I3(GND_net), .O(n2915));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1097_19_lut (.I0(GND_net), .I1(GND_net), .I2(n12192), 
            .I3(n49280), .O(n4911)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_833_4 (.CI(n49515), .I0(n1232_adj_5800), 
            .I1(GND_net), .CO(n49516));
    SB_LUT4 encoder0_position_30__I_0_i1927_3_lut (.I0(n2828), .I1(n2895), 
            .I2(n2841), .I3(GND_net), .O(n2927));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_833_3_lut (.I0(GND_net), .I1(n1233_adj_5801), 
            .I2(VCC_net), .I3(n49514), .O(n1300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1923_3_lut (.I0(n2824), .I1(n2891), 
            .I2(n2841), .I3(GND_net), .O(n2923));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1923_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_833_3 (.CI(n49514), .I0(n1233_adj_5801), 
            .I1(VCC_net), .CO(n49515));
    SB_LUT4 encoder0_position_30__I_0_add_833_2_lut (.I0(GND_net), .I1(n523), 
            .I2(GND_net), .I3(VCC_net), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_833_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1049_3_lut (.I0(n940), .I1(n1601), 
            .I2(n1554), .I3(GND_net), .O(n1633));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i19_3_lut (.I0(encoder0_position[18]), .I1(n14_adj_5700), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1116_3_lut (.I0(n1633), .I1(n1700), 
            .I2(n1653), .I3(GND_net), .O(n1732));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1183_3_lut (.I0(n1732), .I1(n1799), 
            .I2(n1752), .I3(GND_net), .O(n1831));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1250_3_lut (.I0(n1831), .I1(n1898), 
            .I2(n1851), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1317_3_lut (.I0(n1930), .I1(n1997), 
            .I2(n1950), .I3(GND_net), .O(n2029));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1384_3_lut (.I0(n2029), .I1(n2096), 
            .I2(n2049), .I3(GND_net), .O(n2128));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i981_3_lut (.I0(n939), .I1(n1501), 
            .I2(n1455), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1451_3_lut (.I0(n2128), .I1(n2195), 
            .I2(n2148), .I3(GND_net), .O(n2227));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_243_i1_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), .I2(motor_state_23__N_91[0]), 
            .I3(encoder0_position_scaled[0]), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i1048_3_lut (.I0(n1533), .I1(n1600), 
            .I2(n1554), .I3(GND_net), .O(n1632));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1115_3_lut (.I0(n1632), .I1(n1699), 
            .I2(n1653), .I3(GND_net), .O(n1731));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_243_i2_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), .I2(motor_state_23__N_91[1]), 
            .I3(encoder0_position_scaled[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY encoder0_position_30__I_0_add_833_2 (.CI(VCC_net), .I0(n523), 
            .I1(GND_net), .CO(n49514));
    SB_CARRY add_1097_19 (.CI(n49280), .I0(GND_net), .I1(n12192), .CO(n49281));
    SB_LUT4 encoder0_position_30__I_0_i1182_3_lut (.I0(n1731), .I1(n1798), 
            .I2(n1752), .I3(GND_net), .O(n1830));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1097_18_lut (.I0(GND_net), .I1(GND_net), .I2(n12194), 
            .I3(n49279), .O(n4912)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1913_3_lut (.I0(n2814), .I1(n2881), 
            .I2(n2841), .I3(GND_net), .O(n2913));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1913_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1097_18 (.CI(n49279), .I0(GND_net), .I1(n12194), .CO(n49280));
    SB_LUT4 encoder0_position_30__I_0_i1911_3_lut (.I0(n2812), .I1(n2879), 
            .I2(n2841), .I3(GND_net), .O(n2911));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1909_3_lut (.I0(n2810), .I1(n2877), 
            .I2(n2841), .I3(GND_net), .O(n2909));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1918_3_lut (.I0(n2819), .I1(n2886), 
            .I2(n2841), .I3(GND_net), .O(n2918));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_243_i3_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), .I2(motor_state_23__N_91[2]), 
            .I3(encoder0_position_scaled[2]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i1917_3_lut (.I0(n2818), .I1(n2885), 
            .I2(n2841), .I3(GND_net), .O(n2917));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1933_3_lut (.I0(n953), .I1(n2901), 
            .I2(n2841), .I3(GND_net), .O(n2933));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1932_3_lut (.I0(n2833), .I1(n2900), 
            .I2(n2841), .I3(GND_net), .O(n2932));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1932_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_151_29 (.CI(n49173), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n49174));
    SB_LUT4 encoder0_position_30__I_0_add_1302_19_lut (.I0(GND_net), .I1(n1917), 
            .I2(VCC_net), .I3(n49761), .O(n1984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1302_18_lut (.I0(GND_net), .I1(n1918), 
            .I2(VCC_net), .I3(n49760), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_18 (.CI(n49760), .I0(n1918), 
            .I1(VCC_net), .CO(n49761));
    SB_LUT4 encoder0_position_30__I_0_add_1302_17_lut (.I0(GND_net), .I1(n1919), 
            .I2(VCC_net), .I3(n49759), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_17 (.CI(n49759), .I0(n1919), 
            .I1(VCC_net), .CO(n49760));
    SB_LUT4 encoder0_position_30__I_0_i1931_3_lut (.I0(n2832), .I1(n2899), 
            .I2(n2841), .I3(GND_net), .O(n2931));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28320_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), .I2(n42234), 
            .I3(encoder0_position_scaled[3]), .O(n42235));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam i28320_3_lut_4_lut.LUT_INIT = 16'he0f1;
    SB_LUT4 mux_4310_i4_3_lut (.I0(encoder0_position[3]), .I1(n29), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n954));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52897_1_lut (.I0(n2940), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68583));
    defparam i52897_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1910 (.I0(n2923), .I1(n2927), .I2(GND_net), .I3(GND_net), 
            .O(n61344));
    defparam i1_2_lut_adj_1910.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1911 (.I0(n2915), .I1(n2916), .I2(n2925), .I3(GND_net), 
            .O(n61170));
    defparam i1_3_lut_adj_1911.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_243_i5_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), .I2(motor_state_23__N_91[4]), 
            .I3(encoder0_position_scaled[4]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i6_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), .I2(motor_state_23__N_91[5]), 
            .I3(encoder0_position_scaled[5]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i1249_3_lut (.I0(n1830), .I1(n1897), 
            .I2(n1851), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n11579_bdd_4_lut_53651 (.I0(n11579), .I1(current[5]), .I2(duty[8]), 
            .I3(n11577), .O(n69372));
    defparam n11579_bdd_4_lut_53651.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_add_1302_16_lut (.I0(GND_net), .I1(n1920), 
            .I2(VCC_net), .I3(n49758), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1316_3_lut (.I0(n1929), .I1(n1996), 
            .I2(n1950), .I3(GND_net), .O(n2028));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i27698_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), .I2(n41621), 
            .I3(encoder0_position_scaled[6]), .O(n41622));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam i27698_3_lut_4_lut.LUT_INIT = 16'he0f1;
    SB_LUT4 encoder0_position_30__I_0_i1383_3_lut (.I0(n2028), .I1(n2095), 
            .I2(n2049), .I3(GND_net), .O(n2127));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1912 (.I0(n2921), .I1(n61344), .I2(n2924), .I3(n2928), 
            .O(n61348));
    defparam i1_4_lut_adj_1912.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1450_3_lut (.I0(n2127), .I1(n2194), 
            .I2(n2148), .I3(GND_net), .O(n2226));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1450_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1302_16 (.CI(n49758), .I0(n1920), 
            .I1(VCC_net), .CO(n49759));
    SB_LUT4 encoder0_position_30__I_0_add_1302_15_lut (.I0(GND_net), .I1(n1921), 
            .I2(VCC_net), .I3(n49757), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_15 (.CI(n49757), .I0(n1921), 
            .I1(VCC_net), .CO(n49758));
    SB_LUT4 encoder0_position_30__I_0_add_1302_14_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n49756), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_14 (.CI(n49756), .I0(n1922), 
            .I1(VCC_net), .CO(n49757));
    SB_LUT4 i1_4_lut_adj_1913 (.I0(n2922), .I1(n2919), .I2(n2926), .I3(n2920), 
            .O(n60042));
    defparam i1_4_lut_adj_1913.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_1302_13_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n49755), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_13 (.CI(n49755), .I0(n1923), 
            .I1(VCC_net), .CO(n49756));
    SB_LUT4 encoder0_position_30__I_0_i568_3_lut (.I0(n829), .I1(n896), 
            .I2(n861), .I3(GND_net), .O(n928));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_243_i8_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), .I2(motor_state_23__N_91[7]), 
            .I3(encoder0_position_scaled[7]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i29663_4_lut (.I0(n954), .I1(n2931), .I2(n2932), .I3(n2933), 
            .O(n43572));
    defparam i29663_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1914 (.I0(n2917), .I1(n60042), .I2(n2918), .I3(n61348), 
            .O(n61354));
    defparam i1_4_lut_adj_1914.LUT_INIT = 16'hfffe;
    SB_LUT4 i16458_3_lut_4_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30466));   // verilog/coms.v(130[12] 305[6])
    defparam i16458_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mux_1584_i19_3_lut (.I0(duty[21]), .I1(duty[18]), .I2(n260), 
            .I3(GND_net), .O(n12190));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_243_i9_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), .I2(motor_state_23__N_91[8]), 
            .I3(encoder0_position_scaled[8]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_4_lut_adj_1915 (.I0(n2929), .I1(n61354), .I2(n43572), .I3(n2930), 
            .O(n61356));
    defparam i1_4_lut_adj_1915.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1916 (.I0(n2909), .I1(n2911), .I2(n2913), .I3(n61170), 
            .O(n61176));
    defparam i1_4_lut_adj_1916.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_1302_12_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n49754), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_12 (.CI(n49754), .I0(n1924), 
            .I1(VCC_net), .CO(n49755));
    SB_LUT4 encoder0_position_30__I_0_add_1302_11_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n49753), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_11 (.CI(n49753), .I0(n1925), 
            .I1(VCC_net), .CO(n49754));
    SB_LUT4 encoder0_position_30__I_0_add_1302_10_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n49752), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_10 (.CI(n49752), .I0(n1926), 
            .I1(VCC_net), .CO(n49753));
    SB_LUT4 add_151_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n49172), .O(n1213)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1302_9_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n49751), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_9 (.CI(n49751), .I0(n1927), 
            .I1(VCC_net), .CO(n49752));
    SB_LUT4 i1_4_lut_adj_1917 (.I0(n2912), .I1(n2910), .I2(n2914), .I3(n61356), 
            .O(n60010));
    defparam i1_4_lut_adj_1917.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_1302_8_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n49750), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52900_4_lut (.I0(n2908), .I1(n60010), .I2(n2907), .I3(n61176), 
            .O(n2940));
    defparam i52900_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1841_3_lut (.I0(n2710), .I1(n2777), 
            .I2(n2742), .I3(GND_net), .O(n2809));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1844_3_lut (.I0(n2713), .I1(n2780), 
            .I2(n2742), .I3(GND_net), .O(n2812));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28719_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(92[16:31])
    defparam i28719_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY encoder0_position_30__I_0_add_1302_8 (.CI(n49750), .I0(n1928), 
            .I1(VCC_net), .CO(n49751));
    SB_LUT4 encoder0_position_30__I_0_add_1302_7_lut (.I0(GND_net), .I1(n1929), 
            .I2(GND_net), .I3(n49749), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_7 (.CI(n49749), .I0(n1929), 
            .I1(GND_net), .CO(n49750));
    SB_LUT4 encoder0_position_30__I_0_add_1302_6_lut (.I0(GND_net), .I1(n1930), 
            .I2(GND_net), .I3(n49748), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_6 (.CI(n49748), .I0(n1930), 
            .I1(GND_net), .CO(n49749));
    SB_LUT4 encoder0_position_30__I_0_add_1302_5_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n49747), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_5 (.CI(n49747), .I0(n1931), 
            .I1(VCC_net), .CO(n49748));
    SB_LUT4 encoder0_position_30__I_0_i1842_3_lut (.I0(n2711), .I1(n2778), 
            .I2(n2742), .I3(GND_net), .O(n2810));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1843_3_lut (.I0(n2712), .I1(n2779), 
            .I2(n2742), .I3(GND_net), .O(n2811));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1584_i20_3_lut (.I0(duty[22]), .I1(duty[19]), .I2(n260), 
            .I3(GND_net), .O(n12188));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1584_i21_3_lut (.I0(duty[23]), .I1(duty[20]), .I2(n260), 
            .I3(GND_net), .O(n12186));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_4310_i20_3_lut (.I0(encoder0_position[19]), .I1(n13_adj_5701), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n524));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16457_3_lut_4_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30465));   // verilog/coms.v(130[12] 305[6])
    defparam i16457_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i913_3_lut (.I0(n524), .I1(n1401), 
            .I2(n1356), .I3(GND_net), .O(n1433));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i913_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_151_28 (.CI(n49172), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n49173));
    SB_LUT4 encoder0_position_30__I_0_i1857_3_lut (.I0(n2726), .I1(n2793), 
            .I2(n2742), .I3(GND_net), .O(n2825));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1857_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1853_3_lut (.I0(n2722), .I1(n2789), 
            .I2(n2742), .I3(GND_net), .O(n2821));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1853_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1849_3_lut (.I0(n2718), .I1(n2785), 
            .I2(n2742), .I3(GND_net), .O(n2817));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1859_3_lut (.I0(n2728), .I1(n2795), 
            .I2(n2742), .I3(GND_net), .O(n2827));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1854_3_lut (.I0(n2723), .I1(n2790), 
            .I2(n2742), .I3(GND_net), .O(n2822));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1854_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1851_3_lut (.I0(n2720), .I1(n2787), 
            .I2(n2742), .I3(GND_net), .O(n2819));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1858_3_lut (.I0(n2727), .I1(n2794), 
            .I2(n2742), .I3(GND_net), .O(n2826));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1858_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16456_3_lut_4_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30464));   // verilog/coms.v(130[12] 305[6])
    defparam i16456_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1855_3_lut (.I0(n2724), .I1(n2791), 
            .I2(n2742), .I3(GND_net), .O(n2823));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1855_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1852_3_lut (.I0(n2721), .I1(n2788), 
            .I2(n2742), .I3(GND_net), .O(n2820_adj_5813));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i980_3_lut (.I0(n1433), .I1(n1500), 
            .I2(n1455), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1865_3_lut (.I0(n952), .I1(n2801), 
            .I2(n2742), .I3(GND_net), .O(n2833));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1302_4_lut (.I0(GND_net), .I1(n1932), 
            .I2(GND_net), .I3(n49746), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_4 (.CI(n49746), .I0(n1932), 
            .I1(GND_net), .CO(n49747));
    SB_CARRY add_151_4 (.CI(n49148), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n49149));
    SB_LUT4 mux_1584_i22_3_lut (.I0(duty[23]), .I1(duty[21]), .I2(n260), 
            .I3(GND_net), .O(n12184));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_30__I_0_i1864_3_lut (.I0(n2733), .I1(n2800), 
            .I2(n2742), .I3(GND_net), .O(n2832));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i5_3_lut (.I0(encoder0_position[4]), .I1(n28), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n953));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1850_3_lut (.I0(n2719), .I1(n2786), 
            .I2(n2742), .I3(GND_net), .O(n2818));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1848_3_lut (.I0(n2717), .I1(n2784), 
            .I2(n2742), .I3(GND_net), .O(n2816));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1847_3_lut (.I0(n2716), .I1(n2783), 
            .I2(n2742), .I3(GND_net), .O(n2815));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1846_3_lut (.I0(n2715), .I1(n2782), 
            .I2(n2742), .I3(GND_net), .O(n2814));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1302_3_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n49745), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n49154), .O(n1231)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1097_17_lut (.I0(GND_net), .I1(GND_net), .I2(n12196), 
            .I3(n49278), .O(n4913)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_3 (.CI(n49745), .I0(n1933), 
            .I1(VCC_net), .CO(n49746));
    SB_LUT4 encoder0_position_30__I_0_add_1302_2_lut (.I0(GND_net), .I1(n944), 
            .I2(GND_net), .I3(VCC_net), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1302_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1302_2 (.CI(VCC_net), .I0(n944), 
            .I1(GND_net), .CO(n49745));
    SB_LUT4 encoder0_position_30__I_0_i1845_3_lut (.I0(n2714), .I1(n2781), 
            .I2(n2742), .I3(GND_net), .O(n2813));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1860_3_lut (.I0(n2729), .I1(n2796), 
            .I2(n2742), .I3(GND_net), .O(n2828));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53319_1_lut (.I0(n1257), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69005));
    defparam i53319_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1856_3_lut (.I0(n2725), .I1(n2792), 
            .I2(n2742), .I3(GND_net), .O(n2824));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1856_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1863_3_lut (.I0(n2732), .I1(n2799), 
            .I2(n2742), .I3(GND_net), .O(n2831));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1862_3_lut (.I0(n2731), .I1(n2798), 
            .I2(n2742), .I3(GND_net), .O(n2830));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1861_3_lut (.I0(n2730), .I1(n2797), 
            .I2(n2742), .I3(GND_net), .O(n2829));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1861_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1097_17 (.CI(n49278), .I0(GND_net), .I1(n12196), .CO(n49279));
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(clk16MHz), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i52957_1_lut (.I0(n2841), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68643));
    defparam i52957_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_151_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n49171), .O(n1214)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29597_3_lut (.I0(n953), .I1(n2832), .I2(n2833), .I3(GND_net), 
            .O(n43506));
    defparam i29597_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1918 (.I0(n2829), .I1(n43506), .I2(n2830), .I3(n2831), 
            .O(n58765));
    defparam i1_4_lut_adj_1918.LUT_INIT = 16'ha080;
    SB_LUT4 i1_3_lut_adj_1919 (.I0(n2820_adj_5813), .I1(n2823), .I2(n2826), 
            .I3(GND_net), .O(n61548));
    defparam i1_3_lut_adj_1919.LUT_INIT = 16'hfefe;
    SB_LUT4 add_1097_16_lut (.I0(GND_net), .I1(GND_net), .I2(n12198), 
            .I3(n49277), .O(n4914)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_27 (.CI(n49171), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n49172));
    SB_LUT4 i1_4_lut_adj_1920 (.I0(n61548), .I1(n2819), .I2(n2822), .I3(n2827), 
            .O(n61552));
    defparam i1_4_lut_adj_1920.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1921 (.I0(n2817), .I1(n58765), .I2(n2821), .I3(n2825), 
            .O(n59858));
    defparam i1_4_lut_adj_1921.LUT_INIT = 16'hfffe;
    SB_CARRY add_1097_16 (.CI(n49277), .I0(GND_net), .I1(n12198), .CO(n49278));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_33_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_5851), .I3(n50621), .O(n2_adj_5715)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_32_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_5852), .I3(n50620), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1097_15_lut (.I0(GND_net), .I1(GND_net), .I2(n12200), 
            .I3(n49276), .O(n4915)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_32 (.CI(n50620), 
            .I0(GND_net), .I1(n3_adj_5852), .CO(n50621));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_31_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_5853), .I3(n50619), .O(n4_adj_5714)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_31 (.CI(n50619), 
            .I0(GND_net), .I1(n4_adj_5853), .CO(n50620));
    SB_LUT4 mux_1584_i23_3_lut (.I0(duty[23]), .I1(duty[22]), .I2(n260), 
            .I3(GND_net), .O(n12182));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1922 (.I0(n2824), .I1(n2828), .I2(GND_net), .I3(GND_net), 
            .O(n61568));
    defparam i1_2_lut_adj_1922.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1923 (.I0(n2813), .I1(n2814), .I2(n2815), .I3(n61568), 
            .O(n61574));
    defparam i1_4_lut_adj_1923.LUT_INIT = 16'hfffe;
    SB_LUT4 add_151_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n49170), .O(n1215)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_30_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_5854), .I3(n50618), .O(n5_adj_5709)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_30 (.CI(n50618), 
            .I0(GND_net), .I1(n5_adj_5854), .CO(n50619));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_29_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_5855), .I3(n50617), .O(n6_adj_5707)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_29 (.CI(n50617), 
            .I0(GND_net), .I1(n6_adj_5855), .CO(n50618));
    SB_CARRY add_1097_15 (.CI(n49276), .I0(GND_net), .I1(n12200), .CO(n49277));
    SB_LUT4 add_1097_14_lut (.I0(GND_net), .I1(GND_net), .I2(n12202), 
            .I3(n49275), .O(n4916)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_28_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_5856), .I3(n50616), .O(n7_adj_5706)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_28 (.CI(n50616), 
            .I0(GND_net), .I1(n7_adj_5856), .CO(n50617));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_27_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_5857), .I3(n50615), .O(n8_adj_5705)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_27 (.CI(n50615), 
            .I0(GND_net), .I1(n8_adj_5857), .CO(n50616));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_5858), .I3(n50614), .O(n9_adj_5704)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_243_i10_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[9]), .I3(encoder0_position_scaled[9]), 
            .O(motor_state[9]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_26 (.CI(n50614), 
            .I0(GND_net), .I1(n9_adj_5858), .CO(n50615));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_5859), .I3(n50613), .O(n10_adj_5703)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1924 (.I0(n59858), .I1(n2816), .I2(n2818), .I3(n61552), 
            .O(n61558));
    defparam i1_4_lut_adj_1924.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1925 (.I0(n2811), .I1(n2810), .I2(n2812), .I3(n61574), 
            .O(n59879));
    defparam i1_4_lut_adj_1925.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_25 (.CI(n50613), 
            .I0(GND_net), .I1(n10_adj_5859), .CO(n50614));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_5860), .I3(n50612), .O(n11_adj_5702)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52960_4_lut (.I0(n2809), .I1(n2808), .I2(n59879), .I3(n61558), 
            .O(n2841));
    defparam i52960_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_24 (.CI(n50612), 
            .I0(GND_net), .I1(n11_adj_5860), .CO(n50613));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_5861), .I3(n50611), .O(n12)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_23 (.CI(n50611), 
            .I0(GND_net), .I1(n12_adj_5861), .CO(n50612));
    SB_LUT4 encoder0_position_30__I_0_i1775_3_lut (.I0(n2612), .I1(n2679), 
            .I2(n2643), .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(current[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_243_i11_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[10]), .I3(encoder0_position_scaled[10]), 
            .O(motor_state[10]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i28700_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), .I2(motor_state_23__N_91[11]), 
            .I3(encoder0_position_scaled[11]), .O(n1));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam i28700_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i1773_3_lut (.I0(n2610), .I1(n2677), 
            .I2(n2643), .I3(GND_net), .O(n2709));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1774_3_lut (.I0(n2611), .I1(n2678), 
            .I2(n2643), .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1047_3_lut (.I0(n1532), .I1(n1599), 
            .I2(n1554), .I3(GND_net), .O(n1631));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1114_3_lut (.I0(n1631), .I1(n1698), 
            .I2(n1653), .I3(GND_net), .O(n1730));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_5862), .I3(n50610), .O(n13_adj_5701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_22 (.CI(n50610), 
            .I0(GND_net), .I1(n13_adj_5862), .CO(n50611));
    SB_CARRY add_1097_14 (.CI(n49275), .I0(GND_net), .I1(n12202), .CO(n49276));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_5863), .I3(n50609), .O(n14_adj_5700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_21 (.CI(n50609), 
            .I0(GND_net), .I1(n14_adj_5863), .CO(n50610));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_5864), .I3(n50608), .O(n15_adj_5699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_20 (.CI(n50608), 
            .I0(GND_net), .I1(n15_adj_5864), .CO(n50609));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_5865), .I3(n50607), .O(n16_adj_5698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_19 (.CI(n50607), 
            .I0(GND_net), .I1(n16_adj_5865), .CO(n50608));
    SB_LUT4 encoder0_position_30__I_0_i1181_3_lut (.I0(n1730), .I1(n1797), 
            .I2(n1752), .I3(GND_net), .O(n1829));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_5866), .I3(n50606), .O(n17_adj_5697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1778_3_lut (.I0(n2615), .I1(n2682), 
            .I2(n2643), .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1778_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1777_3_lut (.I0(n2614), .I1(n2681), 
            .I2(n2643), .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1776_3_lut (.I0(n2613), .I1(n2680), 
            .I2(n2643), .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1781_3_lut (.I0(n2618), .I1(n2685), 
            .I2(n2643), .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1780_3_lut (.I0(n2617), .I1(n2684), 
            .I2(n2643), .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1248_3_lut (.I0(n1829), .I1(n1896), 
            .I2(n1851), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1248_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1315_3_lut (.I0(n1928), .I1(n1995), 
            .I2(n1950), .I3(GND_net), .O(n2027));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_18 (.CI(n50606), 
            .I0(GND_net), .I1(n17_adj_5866), .CO(n50607));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_5867), .I3(n50605), .O(n18_adj_5696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_17 (.CI(n50605), 
            .I0(GND_net), .I1(n18_adj_5867), .CO(n50606));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_5868), .I3(n50604), .O(n19_adj_5695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1097_13_lut (.I0(GND_net), .I1(GND_net), .I2(n12204), 
            .I3(n49274), .O(n4917)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_16 (.CI(n50604), 
            .I0(GND_net), .I1(n19_adj_5868), .CO(n50605));
    SB_LUT4 encoder0_position_30__I_0_i1779_3_lut (.I0(n2616), .I1(n2683), 
            .I2(n2643), .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_5869), .I3(n50603), .O(n20_adj_5694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_15 (.CI(n50603), 
            .I0(GND_net), .I1(n20_adj_5869), .CO(n50604));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_5870), .I3(n50602), .O(n21_adj_5693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1797_3_lut (.I0(n951), .I1(n2701), 
            .I2(n2643), .I3(GND_net), .O(n2733));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1797_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_14 (.CI(n50602), 
            .I0(GND_net), .I1(n21_adj_5870), .CO(n50603));
    SB_LUT4 encoder0_position_30__I_0_i1796_3_lut (.I0(n2633), .I1(n2700), 
            .I2(n2643), .I3(GND_net), .O(n2732));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1795_3_lut (.I0(n2632), .I1(n2699), 
            .I2(n2643), .I3(GND_net), .O(n2731));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1795_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i6_3_lut (.I0(encoder0_position[5]), .I1(n27), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n952));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_5871), .I3(n50601), .O(n22_adj_5692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_13 (.CI(n50601), 
            .I0(GND_net), .I1(n22_adj_5871), .CO(n50602));
    SB_LUT4 n69372_bdd_4_lut (.I0(n69372), .I1(duty[5]), .I2(n4923), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[5]));
    defparam n69372_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_5872), .I3(n50600), .O(n23_adj_5691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_12 (.CI(n50600), 
            .I0(GND_net), .I1(n23_adj_5872), .CO(n50601));
    SB_LUT4 n11579_bdd_4_lut_53646 (.I0(n11579), .I1(current[4]), .I2(duty[7]), 
            .I3(n11577), .O(n69366));
    defparam n11579_bdd_4_lut_53646.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_i1786_3_lut (.I0(n2623), .I1(n2690), 
            .I2(n2643), .I3(GND_net), .O(n2722));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n69366_bdd_4_lut (.I0(n69366), .I1(duty[4]), .I2(n4924), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[4]));
    defparam n69366_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_5873), .I3(n50599), .O(n24_adj_5690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1784_3_lut (.I0(n2621), .I1(n2688), 
            .I2(n2643), .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_243_i13_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[12]), .I3(encoder0_position_scaled[12]), 
            .O(motor_state[12]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_243_i14_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[13]), .I3(encoder0_position_scaled[13]), 
            .O(motor_state[13]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i1788_3_lut (.I0(n2625), .I1(n2692), 
            .I2(n2643), .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1794_3_lut (.I0(n2631), .I1(n2698), 
            .I2(n2643), .I3(GND_net), .O(n2730));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1382_3_lut (.I0(n2027), .I1(n2094), 
            .I2(n2049), .I3(GND_net), .O(n2126));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1382_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_11 (.CI(n50599), 
            .I0(GND_net), .I1(n24_adj_5873), .CO(n50600));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_5874), .I3(n50598), .O(n25_adj_5689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n11579_bdd_4_lut_53641 (.I0(n11579), .I1(current[3]), .I2(duty[6]), 
            .I3(n11577), .O(n69360));
    defparam n11579_bdd_4_lut_53641.LUT_INIT = 16'he4aa;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_10 (.CI(n50598), 
            .I0(GND_net), .I1(n25_adj_5874), .CO(n50599));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n26_adj_5875), .I3(n50597), .O(n26_adj_5688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_9 (.CI(n50597), 
            .I0(GND_net), .I1(n26_adj_5875), .CO(n50598));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n27_adj_5876), .I3(n50596), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_8 (.CI(n50596), 
            .I0(GND_net), .I1(n27_adj_5876), .CO(n50597));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n28_adj_5877), .I3(n50595), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1793_3_lut (.I0(n2630), .I1(n2697), 
            .I2(n2643), .I3(GND_net), .O(n2729));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1791_3_lut (.I0(n2628), .I1(n2695), 
            .I2(n2643), .I3(GND_net), .O(n2727));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1791_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_7 (.CI(n50595), 
            .I0(GND_net), .I1(n28_adj_5877), .CO(n50596));
    SB_LUT4 encoder0_position_30__I_0_i1789_3_lut (.I0(n2626), .I1(n2693), 
            .I2(n2643), .I3(GND_net), .O(n2725));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1789_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1097_13 (.CI(n49274), .I0(GND_net), .I1(n12204), .CO(n49275));
    SB_LUT4 encoder0_position_30__I_0_i1783_3_lut (.I0(n2620), .I1(n2687), 
            .I2(n2643), .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n29_adj_5878), .I3(n50594), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1782_3_lut (.I0(n2619), .I1(n2686), 
            .I2(n2643), .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1792_3_lut (.I0(n2629), .I1(n2696), 
            .I2(n2643), .I3(GND_net), .O(n2728));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1792_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_6 (.CI(n50594), 
            .I0(GND_net), .I1(n29_adj_5878), .CO(n50595));
    SB_LUT4 encoder0_position_30__I_0_i1790_3_lut (.I0(n2627), .I1(n2694), 
            .I2(n2643), .I3(GND_net), .O(n2726));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1790_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n30_adj_5879), .I3(n50593), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_5 (.CI(n50593), 
            .I0(GND_net), .I1(n30_adj_5879), .CO(n50594));
    SB_LUT4 add_1097_12_lut (.I0(GND_net), .I1(GND_net), .I2(n12206), 
            .I3(n49273), .O(n4918)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n31_adj_5880), .I3(n50592), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1449_3_lut (.I0(n2126), .I1(n2193), 
            .I2(n2148), .I3(GND_net), .O(n2225));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1785_3_lut (.I0(n2622), .I1(n2689), 
            .I2(n2643), .I3(GND_net), .O(n2721));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1787_3_lut (.I0(n2624), .I1(n2691), 
            .I2(n2643), .I3(GND_net), .O(n2723));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_243_i15_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[14]), .I3(encoder0_position_scaled[14]), 
            .O(motor_state[14]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_4 (.CI(n50592), 
            .I0(GND_net), .I1(n31_adj_5880), .CO(n50593));
    SB_LUT4 encoder0_position_30__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n32_adj_5881), .I3(n50591), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_3 (.CI(n50591), 
            .I0(GND_net), .I1(n32_adj_5881), .CO(n50592));
    SB_CARRY encoder0_position_30__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(VCC_net), .CO(n50591));
    SB_CARRY add_1097_12 (.CI(n49273), .I0(GND_net), .I1(n12206), .CO(n49274));
    SB_LUT4 mux_4310_i21_3_lut (.I0(encoder0_position[20]), .I1(n12), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n523));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_243_i19_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[18]), .I3(encoder0_position_scaled[18]), 
            .O(motor_state[18]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i845_3_lut (.I0(n523), .I1(n1301), 
            .I2(n1257), .I3(GND_net), .O(n1333));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i912_3_lut (.I0(n1333), .I1(n1400), 
            .I2(n1356), .I3(GND_net), .O(n1432));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i979_3_lut (.I0(n1432), .I1(n1499), 
            .I2(n1455), .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1046_3_lut (.I0(n1531), .I1(n1598), 
            .I2(n1554), .I3(GND_net), .O(n1630));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_DFF read_197 (.Q(state_7__N_3916[0]), .C(clk16MHz), .D(n60174));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 encoder0_position_30__I_0_i1113_3_lut (.I0(n1630), .I1(n1697), 
            .I2(n1653), .I3(GND_net), .O(n1729));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1180_3_lut (.I0(n1729), .I1(n1796_adj_5808), 
            .I2(n1752), .I3(GND_net), .O(n1828));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1180_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_243_i23_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[22]), .I3(encoder0_position_scaled[22]), 
            .O(motor_state[22]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i1247_3_lut (.I0(n1828), .I1(n1895), 
            .I2(n1851), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1247_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i52990_1_lut (.I0(n2742), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68676));
    defparam i52990_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1314_3_lut (.I0(n1927), .I1(n1994), 
            .I2(n1950), .I3(GND_net), .O(n2026));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1381_3_lut (.I0(n2026), .I1(n2093), 
            .I2(n2049), .I3(GND_net), .O(n2125));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1448_3_lut (.I0(n2125), .I1(n2192), 
            .I2(n2148), .I3(GND_net), .O(n2224));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1448_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1926 (.I0(n2725), .I1(n2727), .I2(GND_net), .I3(GND_net), 
            .O(n61236));
    defparam i1_2_lut_adj_1926.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1927 (.I0(n2723), .I1(n2721), .I2(n2726), .I3(n2728), 
            .O(n61238));
    defparam i1_4_lut_adj_1927.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1928 (.I0(n2724), .I1(n2720), .I2(n61236), .I3(n2722), 
            .O(n61242));
    defparam i1_4_lut_adj_1928.LUT_INIT = 16'hfffe;
    SB_LUT4 i29667_4_lut (.I0(n952), .I1(n2731), .I2(n2732), .I3(n2733), 
            .O(n43576));
    defparam i29667_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 mux_243_i20_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[19]), .I3(encoder0_position_scaled[19]), 
            .O(motor_state[19]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_4_lut_adj_1929 (.I0(n2718), .I1(n2719), .I2(n61242), .I3(n61238), 
            .O(n61248));
    defparam i1_4_lut_adj_1929.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_4310_i22_3_lut (.I0(encoder0_position[21]), .I1(n11_adj_5702), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n522));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1930 (.I0(n2729), .I1(n61248), .I2(n43576), .I3(n2730), 
            .O(n61250));
    defparam i1_4_lut_adj_1930.LUT_INIT = 16'heccc;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_30__I_0_add_1235_18_lut (.I0(GND_net), .I1(n1818), 
            .I2(VCC_net), .I3(n49724), .O(n1885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i777_3_lut (.I0(n522), .I1(n1201), 
            .I2(n1158), .I3(GND_net), .O(n1233_adj_5801));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1931 (.I0(n2715), .I1(n2716), .I2(n61250), .I3(n2717), 
            .O(n61256));
    defparam i1_4_lut_adj_1931.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i844_3_lut (.I0(n1233_adj_5801), .I1(n1300), 
            .I2(n1257), .I3(GND_net), .O(n1332));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i911_3_lut (.I0(n1332), .I1(n1399), 
            .I2(n1356), .I3(GND_net), .O(n1431));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1932 (.I0(n2712), .I1(n2713), .I2(n2714), .I3(n61256), 
            .O(n61262));
    defparam i1_4_lut_adj_1932.LUT_INIT = 16'hfffe;
    SB_LUT4 add_1097_11_lut (.I0(GND_net), .I1(GND_net), .I2(n12208), 
            .I3(n49272), .O(n4919)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52993_4_lut (.I0(n2710), .I1(n2709), .I2(n2711), .I3(n61262), 
            .O(n2742));
    defparam i52993_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i978_3_lut (.I0(n1431), .I1(n1498), 
            .I2(n1455), .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1707_3_lut (.I0(n2512), .I1(n2579), 
            .I2(n2544), .I3(GND_net), .O(n2611));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1714_3_lut (.I0(n2519), .I1(n2586), 
            .I2(n2544), .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1235_17_lut (.I0(GND_net), .I1(n1819), 
            .I2(VCC_net), .I3(n49723), .O(n1886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_17 (.CI(n49723), .I0(n1819), 
            .I1(VCC_net), .CO(n49724));
    SB_LUT4 encoder0_position_30__I_0_i1709_3_lut (.I0(n2514), .I1(n2581), 
            .I2(n2544), .I3(GND_net), .O(n2613));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n69360_bdd_4_lut (.I0(n69360), .I1(duty[3]), .I2(n4925), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[3]));
    defparam n69360_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1708_3_lut (.I0(n2513), .I1(n2580), 
            .I2(n2544), .I3(GND_net), .O(n2612));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1045_3_lut (.I0(n1530), .I1(n1597), 
            .I2(n1554), .I3(GND_net), .O(n1629));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1713_3_lut (.I0(n2518), .I1(n2585), 
            .I2(n2544), .I3(GND_net), .O(n2617));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1720_3_lut (.I0(n2525), .I1(n2592), 
            .I2(n2544), .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1720_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1716_3_lut (.I0(n2521), .I1(n2588), 
            .I2(n2544), .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_243_i22_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[21]), .I3(encoder0_position_scaled[21]), 
            .O(motor_state[21]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i1112_3_lut (.I0(n1629), .I1(n1696), 
            .I2(n1653), .I3(GND_net), .O(n1728));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1719_3_lut (.I0(n2524), .I1(n2591), 
            .I2(n2544), .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1179_3_lut (.I0(n1728), .I1(n1795), 
            .I2(n1752), .I3(GND_net), .O(n1827));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1246_3_lut (.I0(n1827), .I1(n1894), 
            .I2(n1851), .I3(GND_net), .O(n1926));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1246_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1721_3_lut (.I0(n2526), .I1(n2593), 
            .I2(n2544), .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1313_3_lut (.I0(n1926), .I1(n1993), 
            .I2(n1950), .I3(GND_net), .O(n2025));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1933 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [6]), 
            .O(n56882));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1933.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1235_16_lut (.I0(GND_net), .I1(n1820), 
            .I2(VCC_net), .I3(n49722), .O(n1887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_243_i16_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[15]), .I3(encoder0_position_scaled[15]), 
            .O(motor_state[15]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_30__I_0_i1380_3_lut (.I0(n2025), .I1(n2092), 
            .I2(n2049), .I3(GND_net), .O(n2124));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1447_3_lut (.I0(n2124), .I1(n2191), 
            .I2(n2148), .I3(GND_net), .O(n2223));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1934 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [7]), 
            .O(n56881));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1934.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1935 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [0]), 
            .O(n56880));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1935.LUT_INIT = 16'h2300;
    SB_LUT4 n11579_bdd_4_lut_53636 (.I0(n11579), .I1(current[2]), .I2(duty[5]), 
            .I3(n11577), .O(n69354));
    defparam n11579_bdd_4_lut_53636.LUT_INIT = 16'he4aa;
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(clk16MHz), 
           .D(n57805));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 n69354_bdd_4_lut (.I0(n69354), .I1(duty[2]), .I2(n4926), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[2]));
    defparam n69354_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(clk16MHz), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1936 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [1]), 
            .O(n56879));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1936.LUT_INIT = 16'h2300;
    SB_LUT4 n11579_bdd_4_lut_53631 (.I0(n11579), .I1(current[1]), .I2(duty[4]), 
            .I3(n11577), .O(n69348));
    defparam n11579_bdd_4_lut_53631.LUT_INIT = 16'he4aa;
    SB_LUT4 i12_4_lut_adj_1937 (.I0(\data_in_frame[22] [4]), .I1(n28375), 
            .I2(n28428), .I3(rx_data[4]), .O(n56031));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_1937.LUT_INIT = 16'h3a0a;
    SB_LUT4 mux_243_i21_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[20]), .I3(encoder0_position_scaled[20]), 
            .O(motor_state[20]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 n69348_bdd_4_lut (.I0(n69348), .I1(duty[1]), .I2(n4927), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[1]));
    defparam n69348_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 encoder0_position_30__I_0_i1723_3_lut (.I0(n2528), .I1(n2595), 
            .I2(n2544), .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1715_3_lut (.I0(n2520), .I1(n2587), 
            .I2(n2544), .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1718_3_lut (.I0(n2523), .I1(n2590), 
            .I2(n2544), .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1718_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1724_3_lut (.I0(n2529), .I1(n2596), 
            .I2(n2544), .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1724_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1717_3_lut (.I0(n2522), .I1(n2589), 
            .I2(n2544), .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1717_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1722_3_lut (.I0(n2527), .I1(n2594), 
            .I2(n2544), .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1722_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1712_3_lut (.I0(n2517), .I1(n2584), 
            .I2(n2544), .I3(GND_net), .O(n2616));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1711_3_lut (.I0(n2516), .I1(n2583), 
            .I2(n2544), .I3(GND_net), .O(n2615));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1711_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29583_3_lut (.I0(n521), .I1(n1032), .I2(n1033), .I3(GND_net), 
            .O(n43492));
    defparam i29583_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1938 (.I0(n1029), .I1(n43492), .I2(n1030), .I3(n1031), 
            .O(n58643));
    defparam i1_4_lut_adj_1938.LUT_INIT = 16'ha080;
    SB_LUT4 n11579_bdd_4_lut_53626 (.I0(n11579), .I1(current[0]), .I2(duty[3]), 
            .I3(n11577), .O(n69342));
    defparam n11579_bdd_4_lut_53626.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_i1710_3_lut (.I0(n2515), .I1(n2582), 
            .I2(n2544), .I3(GND_net), .O(n2614));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1726_3_lut (.I0(n2531), .I1(n2598), 
            .I2(n2544), .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1726_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1725_3_lut (.I0(n2530), .I1(n2597), 
            .I2(n2544), .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1729_3_lut (.I0(n950), .I1(n2601), 
            .I2(n2544), .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1728_3_lut (.I0(n2533), .I1(n2600), 
            .I2(n2544), .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1727_3_lut (.I0(n2532), .I1(n2599), 
            .I2(n2544), .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_243_i24_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[23]), .I3(encoder0_position_scaled[23]), 
            .O(motor_state[23]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_4310_i7_3_lut (.I0(encoder0_position[6]), .I1(n26_adj_5688), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n951));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), .I2(n19_adj_5811), 
            .I3(encoder0_position_scaled[16]), .O(n20_adj_5812));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i53077_1_lut (.I0(n2643), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68763));
    defparam i53077_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1939 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [2]), 
            .O(n56878));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1939.LUT_INIT = 16'h2300;
    SB_DFF pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[23]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_CARRY encoder0_position_30__I_0_add_1235_16 (.CI(n49722), .I0(n1820), 
            .I1(VCC_net), .CO(n49723));
    SB_LUT4 i1_4_lut_adj_1940 (.I0(n2626), .I1(n2621), .I2(n2628), .I3(n2622), 
            .O(n61538));
    defparam i1_4_lut_adj_1940.LUT_INIT = 16'hfffe;
    SB_LUT4 i53395_4_lut (.I0(n1026), .I1(n58643), .I2(n1027), .I3(n1028), 
            .O(n1059));
    defparam i53395_4_lut.LUT_INIT = 16'h0001;
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[22]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i635_3_lut (.I0(n928), .I1(n995), 
            .I2(n960), .I3(GND_net), .O(n1027));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i635_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[21]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i29651_4_lut (.I0(n522), .I1(n1131), .I2(n1132), .I3(n1133), 
            .O(n43560));
    defparam i29651_4_lut.LUT_INIT = 16'hfcec;
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[20]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_3_lut_adj_1941 (.I0(n1126), .I1(n1127), .I2(n1128), .I3(GND_net), 
            .O(n61002));
    defparam i1_3_lut_adj_1941.LUT_INIT = 16'hfefe;
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[19]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i29669_4_lut (.I0(n951), .I1(n2631), .I2(n2632), .I3(n2633), 
            .O(n43578));
    defparam i29669_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_243_i18_3_lut_4_lut (.I0(n25398), .I1(control_mode[1]), 
            .I2(motor_state_23__N_91[17]), .I3(encoder0_position_scaled[17]), 
            .O(motor_state[17]));   // verilog/TinyFPGA_B.v(285[5:22])
    defparam mux_243_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_2_lut_adj_1942 (.I0(n1129), .I1(n1130), .I2(GND_net), .I3(GND_net), 
            .O(n61308));
    defparam i1_2_lut_adj_1942.LUT_INIT = 16'h8888;
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[18]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1943 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [3]), 
            .O(n56877));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1943.LUT_INIT = 16'h2300;
    SB_LUT4 i53382_4_lut (.I0(n61308), .I1(n1125), .I2(n61002), .I3(n43560), 
            .O(n1158));
    defparam i53382_4_lut.LUT_INIT = 16'h0103;
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[17]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i702_3_lut (.I0(n1027), .I1(n1094), 
            .I2(n1059), .I3(GND_net), .O(n1126));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i702_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[16]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i29579_3_lut (.I0(n523), .I1(n1232_adj_5800), .I2(n1233_adj_5801), 
            .I3(GND_net), .O(n43488));
    defparam i29579_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[15]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_3_lut_adj_1944 (.I0(n1226_adj_5794), .I1(n1227_adj_5795), 
            .I2(n1228_adj_5796), .I3(GND_net), .O(n61314));
    defparam i1_3_lut_adj_1944.LUT_INIT = 16'hfefe;
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[14]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1945 (.I0(n1229_adj_5797), .I1(n43488), .I2(n1230_adj_5798), 
            .I3(n1231_adj_5799), .O(n58640));
    defparam i1_4_lut_adj_1945.LUT_INIT = 16'ha080;
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[13]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i53333_4_lut (.I0(n1225_adj_5793), .I1(n1224_adj_5792), .I2(n58640), 
            .I3(n61314), .O(n1257));
    defparam i53333_4_lut.LUT_INIT = 16'h0001;
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[12]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i769_3_lut (.I0(n1126), .I1(n1193), 
            .I2(n1158), .I3(GND_net), .O(n1225_adj_5793));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i769_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[11]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i29577_3_lut (.I0(n524), .I1(n1332), .I2(n1333), .I3(GND_net), 
            .O(n43486));
    defparam i29577_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[10]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1946 (.I0(n1325), .I1(n1326), .I2(n1327), .I3(n1328), 
            .O(n61148));
    defparam i1_4_lut_adj_1946.LUT_INIT = 16'hfffe;
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[9]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1947 (.I0(n2619), .I1(n2627), .I2(n2625), .I3(n2623), 
            .O(n61514));
    defparam i1_4_lut_adj_1947.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1948 (.I0(n1329), .I1(n43486), .I2(n1330), .I3(n1331), 
            .O(n58638));
    defparam i1_4_lut_adj_1948.LUT_INIT = 16'ha080;
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[8]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i53349_4_lut (.I0(n58638), .I1(n1323), .I2(n1324), .I3(n61148), 
            .O(n1356));
    defparam i53349_4_lut.LUT_INIT = 16'h0001;
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[7]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 encoder0_position_30__I_0_i836_3_lut (.I0(n1225_adj_5793), .I1(n1292), 
            .I2(n1257), .I3(GND_net), .O(n1324));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[6]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i29637_4_lut (.I0(n939), .I1(n1431), .I2(n1432), .I3(n1433), 
            .O(n43546));
    defparam i29637_4_lut.LUT_INIT = 16'hfcec;
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[5]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_2_lut_adj_1949 (.I0(n2629), .I1(n2630), .I2(GND_net), .I3(GND_net), 
            .O(n61732));
    defparam i1_2_lut_adj_1949.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_i1446_3_lut (.I0(n2123), .I1(n2190), 
            .I2(n2148), .I3(GND_net), .O(n2222));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1950 (.I0(n2617), .I1(n61732), .I2(n61514), .I3(n43578), 
            .O(n61518));
    defparam i1_4_lut_adj_1950.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_2_lut_adj_1951 (.I0(n1427), .I1(n1428), .I2(GND_net), .I3(GND_net), 
            .O(n61330));
    defparam i1_2_lut_adj_1951.LUT_INIT = 16'heeee;
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[4]));   // verilog/TinyFPGA_B.v(104[9] 129[5])
    SB_LUT4 i1_4_lut_adj_1952 (.I0(n2614), .I1(n2615), .I2(n2616), .I3(n61518), 
            .O(n61524));
    defparam i1_4_lut_adj_1952.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1953 (.I0(n61538), .I1(n2620), .I2(n2624), .I3(GND_net), 
            .O(n61540));
    defparam i1_3_lut_adj_1953.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1954 (.I0(n2612), .I1(n2610), .I2(n2613), .I3(n61524), 
            .O(n60070));
    defparam i1_4_lut_adj_1954.LUT_INIT = 16'hfffe;
    SB_LUT4 i53080_4_lut (.I0(n2618), .I1(n60070), .I2(n2611), .I3(n61540), 
            .O(n2643));
    defparam i53080_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1955 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [4]), 
            .O(n56876));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1955.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1646_3_lut (.I0(n2419), .I1(n2486), 
            .I2(n2445), .I3(GND_net), .O(n2518));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1645_3_lut (.I0(n2418), .I1(n2485), 
            .I2(n2445), .I3(GND_net), .O(n2517));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1649_3_lut (.I0(n2422), .I1(n2489), 
            .I2(n2445), .I3(GND_net), .O(n2521));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1649_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n27698), 
            .D(n1238), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1956 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [5]), 
            .O(n56875));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1956.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1648_3_lut (.I0(n2421), .I1(n2488), 
            .I2(n2445), .I3(GND_net), .O(n2520));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1647_3_lut (.I0(n2420), .I1(n2487), 
            .I2(n2445), .I3(GND_net), .O(n2519));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1647_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1641_3_lut (.I0(n2414), .I1(n2481), 
            .I2(n2445), .I3(GND_net), .O(n2513));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1640_3_lut (.I0(n2413), .I1(n2480), 
            .I2(n2445), .I3(GND_net), .O(n2512));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1640_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1644_3_lut (.I0(n2417), .I1(n2484), 
            .I2(n2445), .I3(GND_net), .O(n2516));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1644_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1643_3_lut (.I0(n2416), .I1(n2483), 
            .I2(n2445), .I3(GND_net), .O(n2515));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1642_3_lut (.I0(n2415), .I1(n2482), 
            .I2(n2445), .I3(GND_net), .O(n2514));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1656_3_lut (.I0(n2429), .I1(n2496), 
            .I2(n2445), .I3(GND_net), .O(n2528));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1656_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1654_3_lut (.I0(n2427), .I1(n2494), 
            .I2(n2445), .I3(GND_net), .O(n2526));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1654_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1651_3_lut (.I0(n2424), .I1(n2491), 
            .I2(n2445), .I3(GND_net), .O(n2523));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1651_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1653_3_lut (.I0(n2426), .I1(n2493), 
            .I2(n2445), .I3(GND_net), .O(n2525));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1653_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1661_3_lut (.I0(n949), .I1(n2501), 
            .I2(n2445), .I3(GND_net), .O(n2533));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1661_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1660_3_lut (.I0(n2433), .I1(n2500), 
            .I2(n2445), .I3(GND_net), .O(n2532));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1660_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i8_3_lut (.I0(encoder0_position[7]), .I1(n25_adj_5689), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n950));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter__i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n27698), 
            .D(n1237), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n27698), 
            .D(n1236), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n27698), 
            .D(n1235), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n27698), 
            .D(n1234), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n27698), 
            .D(n1233), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n27698), 
            .D(n1232), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n27698), 
            .D(n1231), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n27698), 
            .D(n1230), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i10 (.Q(delay_counter[10]), .C(clk16MHz), .E(n27698), 
            .D(n1229), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i11 (.Q(delay_counter[11]), .C(clk16MHz), .E(n27698), 
            .D(n1228), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i12 (.Q(delay_counter[12]), .C(clk16MHz), .E(n27698), 
            .D(n1227), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i13 (.Q(delay_counter[13]), .C(clk16MHz), .E(n27698), 
            .D(n1226), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i14 (.Q(delay_counter[14]), .C(clk16MHz), .E(n27698), 
            .D(n1225), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i15 (.Q(delay_counter[15]), .C(clk16MHz), .E(n27698), 
            .D(n1224), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i16 (.Q(delay_counter[16]), .C(clk16MHz), .E(n27698), 
            .D(n1223), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i17 (.Q(delay_counter[17]), .C(clk16MHz), .E(n27698), 
            .D(n1222), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i18 (.Q(delay_counter[18]), .C(clk16MHz), .E(n27698), 
            .D(n1221), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i19 (.Q(delay_counter[19]), .C(clk16MHz), .E(n27698), 
            .D(n1220), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i20 (.Q(delay_counter[20]), .C(clk16MHz), .E(n27698), 
            .D(n1219), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_DFFESR delay_counter__i21 (.Q(delay_counter[21]), .C(clk16MHz), .E(n27698), 
            .D(n1218), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 encoder0_position_30__I_0_i1659_3_lut (.I0(n2432), .I1(n2499), 
            .I2(n2445), .I3(GND_net), .O(n2531));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1659_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1658_3_lut (.I0(n2431), .I1(n2498), 
            .I2(n2445), .I3(GND_net), .O(n2530));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1658_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1657_3_lut (.I0(n2430), .I1(n2497), 
            .I2(n2445), .I3(GND_net), .O(n2529));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1657_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1652_3_lut (.I0(n2425), .I1(n2492), 
            .I2(n2445), .I3(GND_net), .O(n2524));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1652_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1957 (.I0(n1424), .I1(n1425), .I2(n1426), .I3(GND_net), 
            .O(n61336));
    defparam i1_3_lut_adj_1957.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_i1650_3_lut (.I0(n2423), .I1(n2490), 
            .I2(n2445), .I3(GND_net), .O(n2522));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1650_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1235_15_lut (.I0(GND_net), .I1(n1821), 
            .I2(VCC_net), .I3(n49721), .O(n1888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1655_3_lut (.I0(n2428), .I1(n2495), 
            .I2(n2445), .I3(GND_net), .O(n2527));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1655_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53048_1_lut (.I0(n2544), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68734));
    defparam i53048_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1235_15 (.CI(n49721), .I0(n1821), 
            .I1(VCC_net), .CO(n49722));
    SB_LUT4 encoder0_position_30__I_0_add_1235_14_lut (.I0(GND_net), .I1(n1822_adj_5809), 
            .I2(VCC_net), .I3(n49720), .O(n1889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_14 (.CI(n49720), .I0(n1822_adj_5809), 
            .I1(VCC_net), .CO(n49721));
    SB_LUT4 i29601_3_lut (.I0(n950), .I1(n2532), .I2(n2533), .I3(GND_net), 
            .O(n43510));
    defparam i29601_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1958 (.I0(n2525), .I1(n2523), .I2(n2526), .I3(n2528), 
            .O(n61118));
    defparam i1_4_lut_adj_1958.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1959 (.I0(n2527), .I1(n61118), .I2(n2522), .I3(n2524), 
            .O(n61120));
    defparam i1_4_lut_adj_1959.LUT_INIT = 16'hfffe;
    SB_LUT4 i16436_3_lut_4_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30444));   // verilog/coms.v(130[12] 305[6])
    defparam i16436_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_4_lut_adj_1960 (.I0(n2529), .I1(n43510), .I2(n2530), .I3(n2531), 
            .O(n58714));
    defparam i1_4_lut_adj_1960.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1961 (.I0(n2519), .I1(n2520), .I2(n2521), .I3(n61120), 
            .O(n61126));
    defparam i1_4_lut_adj_1961.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1962 (.I0(n2517), .I1(n2518), .I2(n61126), .I3(n58714), 
            .O(n61132));
    defparam i1_4_lut_adj_1962.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1963 (.I0(n2514), .I1(n2515), .I2(n2516), .I3(n61132), 
            .O(n61138));
    defparam i1_4_lut_adj_1963.LUT_INIT = 16'hfffe;
    SB_LUT4 i53051_4_lut (.I0(n2512), .I1(n2511), .I2(n2513), .I3(n61138), 
            .O(n2544));
    defparam i53051_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1964 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [6]), 
            .O(n56874));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1964.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1965 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [7]), 
            .O(n56873));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1965.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1966 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [0]), 
            .O(n29046));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1966.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1967 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [1]), 
            .O(n56872));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1967.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1968 (.I0(n1429), .I1(n61330), .I2(n43546), .I3(n1430), 
            .O(n61332));
    defparam i1_4_lut_adj_1968.LUT_INIT = 16'heccc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1969 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [2]), 
            .O(n56871));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1969.LUT_INIT = 16'h2300;
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFFESR dti_counter_1937__i1 (.Q(dti_counter[1]), .C(clk16MHz), .E(n27780), 
            .D(n44), .R(n29162));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1937__i2 (.Q(dti_counter[2]), .C(clk16MHz), .E(n27780), 
            .D(n43_adj_5840), .R(n29162));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1937__i3 (.Q(dti_counter[3]), .C(clk16MHz), .E(n27780), 
            .D(n42), .R(n29162));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1937__i4 (.Q(dti_counter[4]), .C(clk16MHz), .E(n27780), 
            .D(n41), .R(n29162));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1937__i5 (.Q(dti_counter[5]), .C(clk16MHz), .E(n27780), 
            .D(n40), .R(n29162));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1937__i6 (.Q(dti_counter[6]), .C(clk16MHz), .E(n27780), 
            .D(n39), .R(n29162));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_DFFESR dti_counter_1937__i7 (.Q(dti_counter[7]), .C(clk16MHz), .E(n27780), 
            .D(n38_adj_5839), .R(n29162));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 i53368_4_lut (.I0(n1422), .I1(n61332), .I2(n61336), .I3(n1423), 
            .O(n1455));
    defparam i53368_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1970 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [3]), 
            .O(n56870));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1970.LUT_INIT = 16'h2300;
    SB_DFFESR dti_counter_1937__i0 (.Q(dti_counter[0]), .C(clk16MHz), .E(n27780), 
            .D(n45_adj_5841), .R(n29162));   // verilog/TinyFPGA_B.v(174[23:37])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1971 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [4]), 
            .O(n56869));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1971.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1235_13_lut (.I0(GND_net), .I1(n1823), 
            .I2(VCC_net), .I3(n49719), .O(n1890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1972 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [5]), 
            .O(n56868));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1972.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1574_3_lut (.I0(n2315), .I1(n2382), 
            .I2(n2346), .I3(GND_net), .O(n2414));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1973 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [6]), 
            .O(n56867));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1973.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1573_3_lut (.I0(n2314), .I1(n2381), 
            .I2(n2346), .I3(GND_net), .O(n2413));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1580_3_lut (.I0(n2321), .I1(n2388), 
            .I2(n2346), .I3(GND_net), .O(n2420));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i903_3_lut (.I0(n1324), .I1(n1391), 
            .I2(n1356), .I3(GND_net), .O(n1423));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i903_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1577_3_lut (.I0(n2318), .I1(n2385), 
            .I2(n2346), .I3(GND_net), .O(n2417));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1577_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1591_3_lut (.I0(n2332), .I1(n2399), 
            .I2(n2346), .I3(GND_net), .O(n2431));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1591_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1590_3_lut (.I0(n2331), .I1(n2398), 
            .I2(n2346), .I3(GND_net), .O(n2430));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1590_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1235_13 (.CI(n49719), .I0(n1823), 
            .I1(VCC_net), .CO(n49720));
    SB_CARRY add_151_26 (.CI(n49170), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n49171));
    SB_LUT4 encoder0_position_30__I_0_add_1235_12_lut (.I0(GND_net), .I1(n1824_adj_5810), 
            .I2(VCC_net), .I3(n49718), .O(n1891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1589_3_lut (.I0(n2330), .I1(n2397), 
            .I2(n2346), .I3(GND_net), .O(n2429));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1576_3_lut (.I0(n2317), .I1(n2384), 
            .I2(n2346), .I3(GND_net), .O(n2416));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1575_3_lut (.I0(n2316), .I1(n2383), 
            .I2(n2346), .I3(GND_net), .O(n2415));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1585_3_lut (.I0(n2326), .I1(n2393), 
            .I2(n2346), .I3(GND_net), .O(n2425));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1585_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1235_12 (.CI(n49718), .I0(n1824_adj_5810), 
            .I1(VCC_net), .CO(n49719));
    SB_LUT4 encoder0_position_30__I_0_i1583_3_lut (.I0(n2324), .I1(n2391), 
            .I2(n2346), .I3(GND_net), .O(n2423));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1974 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [7]), 
            .O(n56866));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1974.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1581_3_lut (.I0(n2322), .I1(n2389), 
            .I2(n2346), .I3(GND_net), .O(n2421));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1588_3_lut (.I0(n2329), .I1(n2396), 
            .I2(n2346), .I3(GND_net), .O(n2428));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1588_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1586_3_lut (.I0(n2327), .I1(n2394), 
            .I2(n2346), .I3(GND_net), .O(n2426));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_1235_11_lut (.I0(GND_net), .I1(n1825), 
            .I2(VCC_net), .I3(n49717), .O(n1892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1975 (.I0(n1528), .I1(n1527), .I2(GND_net), .I3(GND_net), 
            .O(n61154));
    defparam i1_2_lut_adj_1975.LUT_INIT = 16'heeee;
    SB_LUT4 i29633_4_lut (.I0(n940), .I1(n1531), .I2(n1532), .I3(n1533), 
            .O(n43542));
    defparam i29633_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1976 (.I0(n1524), .I1(n1525), .I2(n1526), .I3(n61154), 
            .O(n61160));
    defparam i1_4_lut_adj_1976.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1977 (.I0(n1529), .I1(n61160), .I2(n43542), .I3(n1530), 
            .O(n61162));
    defparam i1_4_lut_adj_1977.LUT_INIT = 16'heccc;
    SB_LUT4 i53219_4_lut (.I0(n1522), .I1(n1521), .I2(n61162), .I3(n1523), 
            .O(n1554));
    defparam i53219_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i970_3_lut (.I0(n1423), .I1(n1490), 
            .I2(n1455), .I3(GND_net), .O(n1522));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1584_3_lut (.I0(n2325), .I1(n2392), 
            .I2(n2346), .I3(GND_net), .O(n2424));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1038_3_lut (.I0(n1523), .I1(n1590), 
            .I2(n1554), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1037_3_lut (.I0(n1522), .I1(n1589), 
            .I2(n1554), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29565_3_lut (.I0(n941), .I1(n1632), .I2(n1633), .I3(GND_net), 
            .O(n43474));
    defparam i29565_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1978 (.I0(n1625), .I1(n1627), .I2(n1626), .I3(n1628), 
            .O(n61370));
    defparam i1_4_lut_adj_1978.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1979 (.I0(n1629), .I1(n43474), .I2(n1630), .I3(n1631), 
            .O(n58659));
    defparam i1_4_lut_adj_1979.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1980 (.I0(n1623), .I1(n58659), .I2(n1624), .I3(n61370), 
            .O(n61376));
    defparam i1_4_lut_adj_1980.LUT_INIT = 16'hfffe;
    SB_LUT4 i53240_4_lut (.I0(n1621), .I1(n1620), .I2(n1622), .I3(n61376), 
            .O(n1653));
    defparam i53240_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_4310_i17_3_lut (.I0(encoder0_position[16]), .I1(n16_adj_5698), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n941));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1587_3_lut (.I0(n2328), .I1(n2395), 
            .I2(n2346), .I3(GND_net), .O(n2427));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1981 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [0]), 
            .O(n56865));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1981.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1117_3_lut (.I0(n941), .I1(n1701), 
            .I2(n1653), .I3(GND_net), .O(n1733));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1184_3_lut (.I0(n1733), .I1(n1800), 
            .I2(n1752), .I3(GND_net), .O(n1832));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1251_3_lut (.I0(n1832), .I1(n1899), 
            .I2(n1851), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1251_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1982 (.I0(n1728), .I1(n1727), .I2(n1726), .I3(GND_net), 
            .O(n61068));
    defparam i1_3_lut_adj_1982.LUT_INIT = 16'hfefe;
    SB_LUT4 i29585_4_lut (.I0(n942), .I1(n1731), .I2(n1732), .I3(n1733), 
            .O(n43494));
    defparam i29585_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1983 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [1]), 
            .O(n56864));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1983.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1984 (.I0(n1723), .I1(n1724), .I2(n61068), .I3(n1725), 
            .O(n61074));
    defparam i1_4_lut_adj_1984.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1582_3_lut (.I0(n2323), .I1(n2390), 
            .I2(n2346), .I3(GND_net), .O(n2422));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1582_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1985 (.I0(n1729), .I1(n1730), .I2(GND_net), .I3(GND_net), 
            .O(n61382));
    defparam i1_2_lut_adj_1985.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1986 (.I0(n61382), .I1(n1722), .I2(n61074), .I3(n43494), 
            .O(n61078));
    defparam i1_4_lut_adj_1986.LUT_INIT = 16'hfefc;
    SB_CARRY encoder0_position_30__I_0_add_1235_11 (.CI(n49717), .I0(n1825), 
            .I1(VCC_net), .CO(n49718));
    SB_LUT4 i53260_4_lut (.I0(n1720), .I1(n1719), .I2(n1721), .I3(n61078), 
            .O(n1752));
    defparam i53260_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_4310_i16_3_lut (.I0(encoder0_position[15]), .I1(n17_adj_5697), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n942));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1987 (.I0(n1825), .I1(n1826), .I2(n1827), .I3(n1828), 
            .O(n61402));
    defparam i1_4_lut_adj_1987.LUT_INIT = 16'hfffe;
    SB_LUT4 i29657_4_lut (.I0(n943), .I1(n1831), .I2(n1832), .I3(n1833), 
            .O(n43566));
    defparam i29657_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 dti_counter_1937_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[7]), 
            .I3(n50393), .O(n38_adj_5839)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1937_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_1937_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[6]), 
            .I3(n50392), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1937_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1937_add_4_8 (.CI(n50392), .I0(VCC_net), .I1(dti_counter[6]), 
            .CO(n50393));
    SB_LUT4 dti_counter_1937_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[5]), 
            .I3(n50391), .O(n40)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1937_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1937_add_4_7 (.CI(n50391), .I0(VCC_net), .I1(dti_counter[5]), 
            .CO(n50392));
    SB_LUT4 dti_counter_1937_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[4]), 
            .I3(n50390), .O(n41)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1937_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1937_add_4_6 (.CI(n50390), .I0(VCC_net), .I1(dti_counter[4]), 
            .CO(n50391));
    SB_LUT4 dti_counter_1937_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[3]), 
            .I3(n50389), .O(n42)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1937_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1937_add_4_5 (.CI(n50389), .I0(VCC_net), .I1(dti_counter[3]), 
            .CO(n50390));
    SB_LUT4 dti_counter_1937_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[2]), 
            .I3(n50388), .O(n43_adj_5840)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1937_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1937_add_4_4 (.CI(n50388), .I0(VCC_net), .I1(dti_counter[2]), 
            .CO(n50389));
    SB_LUT4 dti_counter_1937_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[1]), 
            .I3(n50387), .O(n44)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1937_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1937_add_4_3 (.CI(n50387), .I0(VCC_net), .I1(dti_counter[1]), 
            .CO(n50388));
    SB_LUT4 dti_counter_1937_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n45_adj_5841)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_1937_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_1937_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(dti_counter[0]), 
            .CO(n50387));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1988 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [2]), 
            .O(n56863));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1988.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1989 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [3]), 
            .O(n56862));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1989.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1990 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [4]), 
            .O(n56861));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1990.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1579_3_lut (.I0(n2320), .I1(n2387), 
            .I2(n2346), .I3(GND_net), .O(n2419));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1578_3_lut (.I0(n2319), .I1(n2386), 
            .I2(n2346), .I3(GND_net), .O(n2418));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1593_3_lut (.I0(n948), .I1(n2401), 
            .I2(n2346), .I3(GND_net), .O(n2433));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1592_3_lut (.I0(n2333), .I1(n2400), 
            .I2(n2346), .I3(GND_net), .O(n2432));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i9_3_lut (.I0(encoder0_position[8]), .I1(n24_adj_5690), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n949));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1991 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [5]), 
            .O(n56860));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1991.LUT_INIT = 16'h2300;
    SB_LUT4 i53017_1_lut (.I0(n2445), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68703));
    defparam i53017_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n55331));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1992 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [6]), 
            .O(n56859));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1992.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1993 (.I0(n2427), .I1(n2424), .I2(n2426), .I3(n2428), 
            .O(n61488));
    defparam i1_4_lut_adj_1993.LUT_INIT = 16'hfffe;
    SB_DFFE commutation_state_i1 (.Q(commutation_state[1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30488));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i29603_3_lut (.I0(n949), .I1(n2432), .I2(n2433), .I3(GND_net), 
            .O(n43512));
    defparam i29603_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1994 (.I0(n2421), .I1(n61488), .I2(n2423), .I3(n2425), 
            .O(n61492));
    defparam i1_4_lut_adj_1994.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1995 (.I0(n2429), .I1(n43512), .I2(n2430), .I3(n2431), 
            .O(n58740));
    defparam i1_4_lut_adj_1995.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1996 (.I0(n2417), .I1(n58740), .I2(n2420), .I3(n61492), 
            .O(n61498));
    defparam i1_4_lut_adj_1996.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1997 (.I0(n2418), .I1(n2419), .I2(n2422), .I3(GND_net), 
            .O(n61582));
    defparam i1_3_lut_adj_1997.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_add_1235_10_lut (.I0(GND_net), .I1(n1826), 
            .I2(VCC_net), .I3(n49716), .O(n1893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_766_11_lut (.I0(n69065), .I1(n1125), 
            .I2(VCC_net), .I3(n49495), .O(n1224_adj_5792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_1235_10 (.CI(n49716), .I0(n1826), 
            .I1(VCC_net), .CO(n49717));
    SB_LUT4 encoder0_position_30__I_0_add_1235_9_lut (.I0(GND_net), .I1(n1827), 
            .I2(VCC_net), .I3(n49715), .O(n1894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_9 (.CI(n49715), .I0(n1827), 
            .I1(VCC_net), .CO(n49716));
    SB_LUT4 encoder0_position_30__I_0_add_1235_8_lut (.I0(GND_net), .I1(n1828), 
            .I2(VCC_net), .I3(n49714), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_766_10_lut (.I0(GND_net), .I1(n1126), 
            .I2(VCC_net), .I3(n49494), .O(n1193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1998 (.I0(n61582), .I1(n2415), .I2(n61498), .I3(n2416), 
            .O(n61502));
    defparam i1_4_lut_adj_1998.LUT_INIT = 16'hfffe;
    SB_LUT4 i53020_4_lut (.I0(n2413), .I1(n2412), .I2(n2414), .I3(n61502), 
            .O(n2445));
    defparam i53020_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_30__I_0_add_766_10 (.CI(n49494), .I0(n1126), 
            .I1(VCC_net), .CO(n49495));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1999 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [7]), 
            .O(n56858));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1999.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2000 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [0]), 
            .O(n29030));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2000.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1511_3_lut (.I0(n2220), .I1(n2287), 
            .I2(n2247), .I3(GND_net), .O(n2319));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2001 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [1]), 
            .O(n56857));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2001.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1522_3_lut (.I0(n2231), .I1(n2298), 
            .I2(n2247), .I3(GND_net), .O(n2330));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2002 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [2]), 
            .O(n56856));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2002.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1521_3_lut (.I0(n2230), .I1(n2297), 
            .I2(n2247), .I3(GND_net), .O(n2329));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1514_3_lut (.I0(n2223), .I1(n2290), 
            .I2(n2247), .I3(GND_net), .O(n2322));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1514_3_lut.LUT_INIT = 16'hacac;
    SB_DFF \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(clk16MHz), 
           .D(n17_adj_5896));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 encoder0_position_30__I_0_i1513_3_lut (.I0(n2222), .I1(n2289), 
            .I2(n2247), .I3(GND_net), .O(n2321));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1512_3_lut (.I0(n2221), .I1(n2288), 
            .I2(n2247), .I3(GND_net), .O(n2320));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1507_3_lut (.I0(n2216), .I1(n2283), 
            .I2(n2247), .I3(GND_net), .O(n2315));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1506_3_lut (.I0(n2215), .I1(n2282), 
            .I2(n2247), .I3(GND_net), .O(n2314));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1506_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1515_3_lut (.I0(n2224), .I1(n2291), 
            .I2(n2247), .I3(GND_net), .O(n2323));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1515_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_2003 (.I0(n1823), .I1(n1824_adj_5810), .I2(n61402), 
            .I3(GND_net), .O(n61406));
    defparam i1_3_lut_adj_2003.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_i1517_3_lut (.I0(n2226), .I1(n2293), 
            .I2(n2247), .I3(GND_net), .O(n2325));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1510_3_lut (.I0(n2219), .I1(n2286), 
            .I2(n2247), .I3(GND_net), .O(n2318));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2004 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [3]), 
            .O(n56855));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2004.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1509_3_lut (.I0(n2218), .I1(n2285), 
            .I2(n2247), .I3(GND_net), .O(n2317));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2005 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [4]), 
            .O(n56854));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2005.LUT_INIT = 16'h2300;
    SB_LUT4 i1_3_lut_adj_2006 (.I0(n1820), .I1(n1821), .I2(n1822_adj_5809), 
            .I3(GND_net), .O(n61412));
    defparam i1_3_lut_adj_2006.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_30__I_0_i1508_3_lut (.I0(n2217), .I1(n2284), 
            .I2(n2247), .I3(GND_net), .O(n2316));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1525_3_lut (.I0(n947), .I1(n2301), 
            .I2(n2247), .I3(GND_net), .O(n2333));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2007 (.I0(n1829), .I1(n61406), .I2(n43566), .I3(n1830), 
            .O(n61408));
    defparam i1_4_lut_adj_2007.LUT_INIT = 16'heccc;
    SB_LUT4 encoder0_position_30__I_0_i1524_3_lut (.I0(n2233), .I1(n2300), 
            .I2(n2247), .I3(GND_net), .O(n2332));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1523_3_lut (.I0(n2232), .I1(n2299), 
            .I2(n2247), .I3(GND_net), .O(n2331));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1523_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1097_11 (.CI(n49272), .I0(GND_net), .I1(n12208), .CO(n49273));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2008 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [5]), 
            .O(n56853));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2008.LUT_INIT = 16'h2300;
    SB_LUT4 mux_4310_i10_3_lut (.I0(encoder0_position[9]), .I1(n23_adj_5691), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n948));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53198_4_lut (.I0(n1818), .I1(n61408), .I2(n61412), .I3(n1819), 
            .O(n1851));
    defparam i53198_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i1516_3_lut (.I0(n2225), .I1(n2292), 
            .I2(n2247), .I3(GND_net), .O(n2324));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1518_3_lut (.I0(n2227), .I1(n2294), 
            .I2(n2247), .I3(GND_net), .O(n2326));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1520_3_lut (.I0(n2229), .I1(n2296), 
            .I2(n2247), .I3(GND_net), .O(n2328));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2009 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [6]), 
            .O(n56852));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2009.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2010 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [7]), 
            .O(n56851));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2010.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1519_3_lut (.I0(n2228), .I1(n2295), 
            .I2(n2247), .I3(GND_net), .O(n2327));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1185_3_lut (.I0(n942), .I1(n1801), 
            .I2(n1752), .I3(GND_net), .O(n1833));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_add_766_9_lut (.I0(GND_net), .I1(n1127), 
            .I2(VCC_net), .I3(n49493), .O(n1194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_8 (.CI(n49714), .I0(n1828), 
            .I1(VCC_net), .CO(n49715));
    SB_CARRY encoder0_position_30__I_0_add_766_9 (.CI(n49493), .I0(n1127), 
            .I1(VCC_net), .CO(n49494));
    SB_LUT4 i52923_1_lut (.I0(n2346), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68609));
    defparam i52923_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_2011 (.I0(n2327), .I1(n2328), .I2(n2326), .I3(n2324), 
            .O(n61274));
    defparam i1_4_lut_adj_2011.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_2012 (.I0(n61274), .I1(n2325), .I2(n2323), .I3(GND_net), 
            .O(n61276));
    defparam i1_3_lut_adj_2012.LUT_INIT = 16'hfefe;
    SB_LUT4 i29675_4_lut (.I0(n948), .I1(n2331), .I2(n2332), .I3(n2333), 
            .O(n43584));
    defparam i29675_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2013 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [0]), 
            .O(n56850));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2013.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_2014 (.I0(n2320), .I1(n2321), .I2(n61276), .I3(n2322), 
            .O(n61282));
    defparam i1_4_lut_adj_2014.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_1235_7_lut (.I0(GND_net), .I1(n1829), 
            .I2(GND_net), .I3(n49713), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_7 (.CI(n49713), .I0(n1829), 
            .I1(GND_net), .CO(n49714));
    SB_LUT4 i1_2_lut_adj_2015 (.I0(n2329), .I1(n2330), .I2(GND_net), .I3(GND_net), 
            .O(n61478));
    defparam i1_2_lut_adj_2015.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_add_766_8_lut (.I0(GND_net), .I1(n1128), 
            .I2(VCC_net), .I3(n49492), .O(n1195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_8 (.CI(n49492), .I0(n1128), 
            .I1(VCC_net), .CO(n49493));
    SB_LUT4 i1_4_lut_adj_2016 (.I0(n2319), .I1(n61478), .I2(n61282), .I3(n43584), 
            .O(n61286));
    defparam i1_4_lut_adj_2016.LUT_INIT = 16'hfefa;
    SB_LUT4 encoder0_position_30__I_0_add_1235_6_lut (.I0(GND_net), .I1(n1830), 
            .I2(GND_net), .I3(n49712), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_766_7_lut (.I0(GND_net), .I1(n1129), 
            .I2(GND_net), .I3(n49491), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_2017 (.I0(n2316), .I1(n2317), .I2(n2318), .I3(n61286), 
            .O(n61292));
    defparam i1_4_lut_adj_2017.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_add_1235_6 (.CI(n49712), .I0(n1830), 
            .I1(GND_net), .CO(n49713));
    SB_LUT4 encoder0_position_30__I_0_add_1235_5_lut (.I0(GND_net), .I1(n1831), 
            .I2(VCC_net), .I3(n49711), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2018 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [1]), 
            .O(n56849));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2018.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2019 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [2]), 
            .O(n56775));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2019.LUT_INIT = 16'h2300;
    SB_LUT4 i3_4_lut_adj_2020 (.I0(\data_in_frame[12] [6]), .I1(n25864), 
            .I2(\data_in_frame[10] [1]), .I3(\data_in_frame[12] [5]), .O(n57361));
    defparam i3_4_lut_adj_2020.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_2021 (.I0(\data_in_frame[14] [5]), .I1(n57720), 
            .I2(n57503), .I3(n57361), .O(n57717));
    defparam i3_4_lut_adj_2021.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2022 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [3]), 
            .O(n56777));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2022.LUT_INIT = 16'h2300;
    SB_LUT4 i4_4_lut_adj_2023 (.I0(n57473), .I1(\data_in_frame[14] [6]), 
            .I2(\data_in_frame[17] [1]), .I3(n57717), .O(n10_adj_5903));
    defparam i4_4_lut_adj_2023.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2024 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [4]), 
            .O(n56778));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2024.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1235_5 (.CI(n49711), .I0(n1831), 
            .I1(VCC_net), .CO(n49712));
    SB_LUT4 i52926_4_lut (.I0(n2314), .I1(n2313), .I2(n2315), .I3(n61292), 
            .O(n2346));
    defparam i52926_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2025 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [5]), 
            .O(n56779));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2025.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_adj_2026 (.I0(\data_in_frame[14] [5]), .I1(n26482), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5892));
    defparam i1_2_lut_adj_2026.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_2027 (.I0(\data_in_frame[10] [1]), .I1(\data_in_frame[12] [4]), 
            .I2(n57503), .I3(n6_adj_5892), .O(n59574));
    defparam i4_4_lut_adj_2027.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2028 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [6]), 
            .O(n56780));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2028.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2029 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [7]), 
            .O(n56781));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2029.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1235_4_lut (.I0(GND_net), .I1(n1832), 
            .I2(GND_net), .I3(n49710), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_4 (.CI(n49710), .I0(n1832), 
            .I1(GND_net), .CO(n49711));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2030 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [0]), 
            .O(n56783));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2030.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2031 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [1]), 
            .O(n56784));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2031.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1235_3_lut (.I0(GND_net), .I1(n1833), 
            .I2(VCC_net), .I3(n49709), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1235_3 (.CI(n49709), .I0(n1833), 
            .I1(VCC_net), .CO(n49710));
    SB_LUT4 encoder0_position_30__I_0_add_1235_2_lut (.I0(GND_net), .I1(n943), 
            .I2(GND_net), .I3(VCC_net), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1235_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1439_3_lut (.I0(n2116), .I1(n2183), 
            .I2(n2148), .I3(GND_net), .O(n2215));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i53171_1_lut (.I0(n2247), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68857));
    defparam i53171_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1235_2 (.CI(VCC_net), .I0(n943), 
            .I1(GND_net), .CO(n49709));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2032 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [2]), 
            .O(n56785));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2032.LUT_INIT = 16'h2300;
    SB_LUT4 i16390_3_lut_4_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30398));   // verilog/coms.v(130[12] 305[6])
    defparam i16390_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_4_lut_adj_2033 (.I0(n2223), .I1(n2227), .I2(n2224), .I3(n2226), 
            .O(n61456));
    defparam i1_4_lut_adj_2033.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(\data_in_frame[13] [6]), .I1(\data_in_frame[16] [1]), 
            .I2(\data_in_frame[15] [6]), .I3(GND_net), .O(n57780));
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_2034 (.I0(n2222), .I1(n2225), .I2(n2228), .I3(GND_net), 
            .O(n61458));
    defparam i1_3_lut_adj_2034.LUT_INIT = 16'hfefe;
    SB_LUT4 i29677_4_lut (.I0(n947), .I1(n2231), .I2(n2232), .I3(n2233), 
            .O(n43586));
    defparam i29677_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_2035 (.I0(n2220), .I1(n2221), .I2(n61458), .I3(n61456), 
            .O(n61464));
    defparam i1_4_lut_adj_2035.LUT_INIT = 16'hfffe;
    SB_LUT4 i16388_3_lut_4_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30396));   // verilog/coms.v(130[12] 305[6])
    defparam i16388_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_4_lut_adj_2036 (.I0(n2229), .I1(n61464), .I2(n43586), .I3(n2230), 
            .O(n61466));
    defparam i1_4_lut_adj_2036.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_2037 (.I0(n2217), .I1(n2218), .I2(n61466), .I3(n2219), 
            .O(n61472));
    defparam i1_4_lut_adj_2037.LUT_INIT = 16'hfffe;
    SB_LUT4 i53174_4_lut (.I0(n2215), .I1(n2214), .I2(n2216), .I3(n61472), 
            .O(n2247));
    defparam i53174_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i16387_3_lut_4_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30395));   // verilog/coms.v(130[12] 305[6])
    defparam i16387_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i4_4_lut_adj_2038 (.I0(n57701), .I1(n57125), .I2(\data_in_frame[13] [4]), 
            .I3(n57780), .O(n10_adj_5899));
    defparam i4_4_lut_adj_2038.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2039 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [3]), 
            .O(n56786));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2039.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2040 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [4]), 
            .O(n56787));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2040.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2041 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [5]), 
            .O(n56788));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2041.LUT_INIT = 16'h2300;
    SB_DFF reset_198 (.Q(reset), .C(clk16MHz), .D(n55417));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 add_2510_25_lut (.I0(n69078), .I1(n2_adj_5851), .I2(n1059), 
            .I3(n50149), .O(encoder0_position_scaled_23__N_43[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_2510_24_lut (.I0(n69065), .I1(n2_adj_5851), .I2(n1158), 
            .I3(n50148), .O(encoder0_position_scaled_23__N_43[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_24 (.CI(n50148), .I0(n2_adj_5851), .I1(n1158), .CO(n50149));
    SB_LUT4 add_2510_23_lut (.I0(n69005), .I1(n2_adj_5851), .I2(n1257), 
            .I3(n50147), .O(encoder0_position_scaled_23__N_43[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_23 (.CI(n50147), .I0(n2_adj_5851), .I1(n1257), .CO(n50148));
    SB_LUT4 add_2510_22_lut (.I0(n69032), .I1(n2_adj_5851), .I2(n1356), 
            .I3(n50146), .O(encoder0_position_scaled_23__N_43[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_22 (.CI(n50146), .I0(n2_adj_5851), .I1(n1356), .CO(n50147));
    SB_LUT4 add_2510_21_lut (.I0(n69051), .I1(n2_adj_5851), .I2(n1455), 
            .I3(n50145), .O(encoder0_position_scaled_23__N_43[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_21 (.CI(n50145), .I0(n2_adj_5851), .I1(n1455), .CO(n50146));
    SB_LUT4 add_2510_20_lut (.I0(n68902), .I1(n2_adj_5851), .I2(n1554), 
            .I3(n50144), .O(encoder0_position_scaled_23__N_43[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_20 (.CI(n50144), .I0(n2_adj_5851), .I1(n1554), .CO(n50145));
    SB_CARRY encoder0_position_30__I_0_add_766_7 (.CI(n49491), .I0(n1129), 
            .I1(GND_net), .CO(n49492));
    SB_LUT4 add_2510_19_lut (.I0(n68923), .I1(n2_adj_5851), .I2(n1653), 
            .I3(n50143), .O(encoder0_position_scaled_23__N_43[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2042 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [6]), 
            .O(n56789));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2042.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2043 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [7]), 
            .O(n56790));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2043.LUT_INIT = 16'h2300;
    SB_LUT4 add_1097_10_lut (.I0(GND_net), .I1(GND_net), .I2(n12210), 
            .I3(n49271), .O(n4920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53122_1_lut (.I0(n2049), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68808));
    defparam i53122_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53099_1_lut (.I0(n1950), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68785));
    defparam i53099_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2510_19 (.CI(n50143), .I0(n2_adj_5851), .I1(n1653), .CO(n50144));
    SB_LUT4 add_2510_18_lut (.I0(n68943), .I1(n2_adj_5851), .I2(n1752), 
            .I3(n50142), .O(encoder0_position_scaled_23__N_43[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2044 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [0]), 
            .O(n56791));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2044.LUT_INIT = 16'h2300;
    SB_CARRY add_2510_18 (.CI(n50142), .I0(n2_adj_5851), .I1(n1752), .CO(n50143));
    SB_LUT4 i16376_3_lut_4_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30384));   // verilog/coms.v(130[12] 305[6])
    defparam i16376_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2045 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [1]), 
            .O(n56792));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2045.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2046 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [2]), 
            .O(n56793));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2046.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_766_6_lut (.I0(GND_net), .I1(n1130), 
            .I2(GND_net), .I3(n49490), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2510_17_lut (.I0(n68881), .I1(n2_adj_5851), .I2(n1851), 
            .I3(n50141), .O(encoder0_position_scaled_23__N_43[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_30__I_0_add_766_6 (.CI(n49490), .I0(n1130), 
            .I1(GND_net), .CO(n49491));
    SB_CARRY add_2510_17 (.CI(n50141), .I0(n2_adj_5851), .I1(n1851), .CO(n50142));
    SB_LUT4 add_2510_16_lut (.I0(n68785), .I1(n2_adj_5851), .I2(n1950), 
            .I3(n50140), .O(encoder0_position_scaled_23__N_43[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2047 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [3]), 
            .O(n56774));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2047.LUT_INIT = 16'h2300;
    SB_CARRY add_2510_16 (.CI(n50140), .I0(n2_adj_5851), .I1(n1950), .CO(n50141));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2048 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [4]), 
            .O(n56794));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2048.LUT_INIT = 16'h2300;
    SB_LUT4 i53195_1_lut (.I0(n1851), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68881));
    defparam i53195_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53257_1_lut (.I0(n1752), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68943));
    defparam i53257_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2510_15_lut (.I0(n68808), .I1(n2_adj_5851), .I2(n2049), 
            .I3(n50139), .O(encoder0_position_scaled_23__N_43[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2049 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [5]), 
            .O(n56795));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2049.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2050 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [6]), 
            .O(n56796));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2050.LUT_INIT = 16'h2300;
    SB_CARRY add_2510_15 (.CI(n50139), .I0(n2_adj_5851), .I1(n2049), .CO(n50140));
    SB_LUT4 add_2510_14_lut (.I0(n68812), .I1(n2_adj_5851), .I2(n2148), 
            .I3(n50138), .O(encoder0_position_scaled_23__N_43[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_14 (.CI(n50138), .I0(n2_adj_5851), .I1(n2148), .CO(n50139));
    SB_LUT4 add_2510_13_lut (.I0(n68857), .I1(n2_adj_5851), .I2(n2247), 
            .I3(n50137), .O(encoder0_position_scaled_23__N_43[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_13 (.CI(n50137), .I0(n2_adj_5851), .I1(n2247), .CO(n50138));
    SB_LUT4 mux_1584_i9_3_lut (.I0(duty[11]), .I1(duty[8]), .I2(n260), 
            .I3(GND_net), .O(n12210));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2051 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [7]), 
            .O(n56797));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2051.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2052 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [0]), 
            .O(n56798));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2052.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2053 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [1]), 
            .O(n56799));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2053.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2054 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [2]), 
            .O(n56800));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2054.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2055 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [3]), 
            .O(n56801));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2055.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2056 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [4]), 
            .O(n56802));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2056.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2057 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [5]), 
            .O(n56803));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2057.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2058 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [6]), 
            .O(n56804));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2058.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2059 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [7]), 
            .O(n56805));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2059.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2060 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [0]), 
            .O(n56806));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2060.LUT_INIT = 16'h2300;
    \quadrature_decoder(1)_U0  quad_counter0 (.b_prev(b_prev), .GND_net(GND_net), 
            .a_new({a_new[1], Open_3}), .position_31__N_3827(position_31__N_3827), 
            .ENCODER0_B_N_keep(ENCODER0_B_N), .n1779(clk16MHz), .ENCODER0_A_N_keep(ENCODER0_A_N), 
            .n29724(n29724), .n1742(n1742), .n1744(n1744), .\encoder0_position[30] (encoder0_position[30]), 
            .\encoder0_position[29] (encoder0_position[29]), .\encoder0_position[28] (encoder0_position[28]), 
            .\encoder0_position[27] (encoder0_position[27]), .\encoder0_position[26] (encoder0_position[26]), 
            .\encoder0_position[25] (encoder0_position[25]), .\encoder0_position[24] (encoder0_position[24]), 
            .\encoder0_position[23] (encoder0_position[23]), .\encoder0_position[22] (encoder0_position[22]), 
            .\encoder0_position[21] (encoder0_position[21]), .\encoder0_position[20] (encoder0_position[20]), 
            .\encoder0_position[19] (encoder0_position[19]), .\encoder0_position[18] (encoder0_position[18]), 
            .\encoder0_position[17] (encoder0_position[17]), .\encoder0_position[16] (encoder0_position[16]), 
            .\encoder0_position[15] (encoder0_position[15]), .\encoder0_position[14] (encoder0_position[14]), 
            .\encoder0_position[13] (encoder0_position[13]), .\encoder0_position[12] (encoder0_position[12]), 
            .\encoder0_position[11] (encoder0_position[11]), .\encoder0_position[10] (encoder0_position[10]), 
            .\encoder0_position[9] (encoder0_position[9]), .\encoder0_position[8] (encoder0_position[8]), 
            .\encoder0_position[7] (encoder0_position[7]), .\encoder0_position[6] (encoder0_position[6]), 
            .\encoder0_position[5] (encoder0_position[5]), .\encoder0_position[4] (encoder0_position[4]), 
            .\encoder0_position[3] (encoder0_position[3]), .\encoder0_position[2] (encoder0_position[2]), 
            .\encoder0_position[1] (encoder0_position[1]), .\encoder0_position[0] (encoder0_position[0]), 
            .VCC_net(VCC_net)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(304[49] 310[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2061 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [1]), 
            .O(n28989));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2061.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2062 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [2]), 
            .O(n56807));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2062.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2510_12_lut (.I0(n68609), .I1(n2_adj_5851), .I2(n2346), 
            .I3(n50136), .O(encoder0_position_scaled_23__N_43[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_12_lut.LUT_INIT = 16'h8BB8;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .clk16MHz(clk16MHz), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    SB_CARRY add_2510_12 (.CI(n50136), .I0(n2_adj_5851), .I1(n2346), .CO(n50137));
    SB_LUT4 add_2510_11_lut (.I0(n68703), .I1(n2_adj_5851), .I2(n2445), 
            .I3(n50135), .O(encoder0_position_scaled_23__N_43[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_11_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2063 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [3]), 
            .O(n28987));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2063.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2064 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [4]), 
            .O(n56808));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2064.LUT_INIT = 16'h2300;
    SB_CARRY add_2510_11 (.CI(n50135), .I0(n2_adj_5851), .I1(n2445), .CO(n50136));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2065 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [5]), 
            .O(n56809));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2065.LUT_INIT = 16'h2300;
    SB_LUT4 add_2510_10_lut (.I0(n68734), .I1(n2_adj_5851), .I2(n2544), 
            .I3(n50134), .O(encoder0_position_scaled_23__N_43[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_10 (.CI(n50134), .I0(n2_adj_5851), .I1(n2544), .CO(n50135));
    SB_LUT4 n69342_bdd_4_lut (.I0(n69342), .I1(duty[0]), .I2(n4928), .I3(n11577), 
            .O(pwm_setpoint_23__N_3[0]));
    defparam n69342_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_2510_9_lut (.I0(n68763), .I1(n2_adj_5851), .I2(n2643), 
            .I3(n50133), .O(encoder0_position_scaled_23__N_43[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2066 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [6]), 
            .O(n56810));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2066.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2067 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [7]), 
            .O(n56811));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2067.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_766_5_lut (.I0(GND_net), .I1(n1131), 
            .I2(VCC_net), .I3(n49489), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2510_9 (.CI(n50133), .I0(n2_adj_5851), .I1(n2643), .CO(n50134));
    SB_LUT4 add_2510_8_lut (.I0(n68676), .I1(n2_adj_5851), .I2(n2742), 
            .I3(n50132), .O(encoder0_position_scaled_23__N_43[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_8 (.CI(n50132), .I0(n2_adj_5851), .I1(n2742), .CO(n50133));
    SB_LUT4 add_2510_7_lut (.I0(n68643), .I1(n2_adj_5851), .I2(n2841), 
            .I3(n50131), .O(encoder0_position_scaled_23__N_43[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_7 (.CI(n50131), .I0(n2_adj_5851), .I1(n2841), .CO(n50132));
    SB_LUT4 add_2510_6_lut (.I0(n68583), .I1(n2_adj_5851), .I2(n2940), 
            .I3(n50130), .O(encoder0_position_scaled_23__N_43[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_6 (.CI(n50130), .I0(n2_adj_5851), .I1(n2940), .CO(n50131));
    SB_CARRY encoder0_position_30__I_0_add_766_5 (.CI(n49489), .I0(n1131), 
            .I1(VCC_net), .CO(n49490));
    SB_CARRY add_1097_10 (.CI(n49271), .I0(GND_net), .I1(n12210), .CO(n49272));
    SB_LUT4 add_2510_5_lut (.I0(n68551), .I1(n2_adj_5851), .I2(n3039), 
            .I3(n50129), .O(encoder0_position_scaled_23__N_43[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_5_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_30__I_0_add_766_4_lut (.I0(GND_net), .I1(n1132), 
            .I2(GND_net), .I3(n49488), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2510_5 (.CI(n50129), .I0(n2_adj_5851), .I1(n3039), .CO(n50130));
    SB_LUT4 add_2510_4_lut (.I0(n68512), .I1(n2_adj_5851), .I2(n3138), 
            .I3(n50128), .O(encoder0_position_scaled_23__N_43[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_4 (.CI(n50128), .I0(n2_adj_5851), .I1(n3138), .CO(n50129));
    SB_LUT4 add_2510_3_lut (.I0(n68450), .I1(n2_adj_5851), .I2(n3237), 
            .I3(n50127), .O(encoder0_position_scaled_23__N_43[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_30__I_0_add_766_4 (.CI(n49488), .I0(n1132), 
            .I1(GND_net), .CO(n49489));
    SB_LUT4 add_1097_9_lut (.I0(GND_net), .I1(GND_net), .I2(n12212), .I3(n49270), 
            .O(n4921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2510_3 (.CI(n50127), .I0(n2_adj_5851), .I1(n3237), .CO(n50128));
    SB_LUT4 add_2510_2_lut (.I0(n68442), .I1(n2_adj_5851), .I2(n43530), 
            .I3(VCC_net), .O(encoder0_position_scaled_23__N_43[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2510_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2510_2 (.CI(VCC_net), .I0(n2_adj_5851), .I1(n43530), 
            .CO(n50127));
    SB_LUT4 encoder0_position_30__I_0_add_2173_33_lut (.I0(n68450), .I1(n3204), 
            .I2(VCC_net), .I3(n50126), .O(n62365)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_2173_32_lut (.I0(GND_net), .I1(n3205), 
            .I2(VCC_net), .I3(n50125), .O(n3272)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_32 (.CI(n50125), .I0(n3205), 
            .I1(VCC_net), .CO(n50126));
    SB_LUT4 encoder0_position_30__I_0_add_2173_31_lut (.I0(GND_net), .I1(n3206), 
            .I2(VCC_net), .I3(n50124), .O(n3273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_31 (.CI(n50124), .I0(n3206), 
            .I1(VCC_net), .CO(n50125));
    SB_LUT4 encoder0_position_30__I_0_add_2173_30_lut (.I0(GND_net), .I1(n3207), 
            .I2(VCC_net), .I3(n50123), .O(n3274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_30 (.CI(n50123), .I0(n3207), 
            .I1(VCC_net), .CO(n50124));
    SB_LUT4 encoder0_position_30__I_0_add_2173_29_lut (.I0(GND_net), .I1(n3208), 
            .I2(VCC_net), .I3(n50122), .O(n3275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_29 (.CI(n50122), .I0(n3208), 
            .I1(VCC_net), .CO(n50123));
    SB_LUT4 encoder0_position_30__I_0_add_2173_28_lut (.I0(GND_net), .I1(n3209), 
            .I2(VCC_net), .I3(n50121), .O(n3276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_766_3_lut (.I0(GND_net), .I1(n1133), 
            .I2(VCC_net), .I3(n49487), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_28 (.CI(n50121), .I0(n3209), 
            .I1(VCC_net), .CO(n50122));
    SB_LUT4 encoder0_position_30__I_0_add_2173_27_lut (.I0(GND_net), .I1(n3210), 
            .I2(VCC_net), .I3(n50120), .O(n3277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_27 (.CI(n50120), .I0(n3210), 
            .I1(VCC_net), .CO(n50121));
    SB_LUT4 encoder0_position_30__I_0_add_2173_26_lut (.I0(GND_net), .I1(n3211), 
            .I2(VCC_net), .I3(n50119), .O(n3278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_26 (.CI(n50119), .I0(n3211), 
            .I1(VCC_net), .CO(n50120));
    SB_LUT4 encoder0_position_30__I_0_add_2173_25_lut (.I0(GND_net), .I1(n3212), 
            .I2(VCC_net), .I3(n50118), .O(n3279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i53237_1_lut (.I0(n1653), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68923));
    defparam i53237_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_2173_25 (.CI(n50118), .I0(n3212), 
            .I1(VCC_net), .CO(n50119));
    SB_LUT4 encoder0_position_30__I_0_add_2173_24_lut (.I0(GND_net), .I1(n3213), 
            .I2(VCC_net), .I3(n50117), .O(n3280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_24 (.CI(n50117), .I0(n3213), 
            .I1(VCC_net), .CO(n50118));
    SB_LUT4 encoder0_position_30__I_0_add_2173_23_lut (.I0(GND_net), .I1(n3214), 
            .I2(VCC_net), .I3(n50116), .O(n3281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_23 (.CI(n50116), .I0(n3214), 
            .I1(VCC_net), .CO(n50117));
    SB_LUT4 encoder0_position_30__I_0_add_2173_22_lut (.I0(GND_net), .I1(n3215), 
            .I2(VCC_net), .I3(n50115), .O(n3282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_22 (.CI(n50115), .I0(n3215), 
            .I1(VCC_net), .CO(n50116));
    SB_LUT4 encoder0_position_30__I_0_add_2173_21_lut (.I0(GND_net), .I1(n3216), 
            .I2(VCC_net), .I3(n50114), .O(n3283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_21 (.CI(n50114), .I0(n3216), 
            .I1(VCC_net), .CO(n50115));
    SB_CARRY encoder0_position_30__I_0_add_766_3 (.CI(n49487), .I0(n1133), 
            .I1(VCC_net), .CO(n49488));
    SB_LUT4 encoder0_position_30__I_0_add_2173_20_lut (.I0(GND_net), .I1(n3217), 
            .I2(VCC_net), .I3(n50113), .O(n3284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_20 (.CI(n50113), .I0(n3217), 
            .I1(VCC_net), .CO(n50114));
    SB_LUT4 encoder0_position_30__I_0_add_2173_19_lut (.I0(GND_net), .I1(n3218), 
            .I2(VCC_net), .I3(n50112), .O(n3285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2068 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [0]), 
            .O(n56812));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2068.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_2173_19 (.CI(n50112), .I0(n3218), 
            .I1(VCC_net), .CO(n50113));
    SB_LUT4 encoder0_position_30__I_0_add_2173_18_lut (.I0(GND_net), .I1(n3219), 
            .I2(VCC_net), .I3(n50111), .O(n3286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_18 (.CI(n50111), .I0(n3219), 
            .I1(VCC_net), .CO(n50112));
    SB_LUT4 encoder0_position_30__I_0_add_2173_17_lut (.I0(GND_net), .I1(n3220), 
            .I2(VCC_net), .I3(n50110), .O(n3287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_17 (.CI(n50110), .I0(n3220), 
            .I1(VCC_net), .CO(n50111));
    SB_LUT4 encoder0_position_30__I_0_add_2173_16_lut (.I0(GND_net), .I1(n3221), 
            .I2(VCC_net), .I3(n50109), .O(n3288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2069 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [1]), 
            .O(n28981));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2069.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_766_2_lut (.I0(GND_net), .I1(n522), 
            .I2(GND_net), .I3(VCC_net), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_766_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_16 (.CI(n50109), .I0(n3221), 
            .I1(VCC_net), .CO(n50110));
    SB_LUT4 encoder0_position_30__I_0_add_2173_15_lut (.I0(GND_net), .I1(n3222), 
            .I2(VCC_net), .I3(n50108), .O(n3289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_766_2 (.CI(VCC_net), .I0(n522), 
            .I1(GND_net), .CO(n49487));
    SB_CARRY encoder0_position_30__I_0_add_2173_15 (.CI(n50108), .I0(n3222), 
            .I1(VCC_net), .CO(n50109));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2070 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [2]), 
            .O(n56813));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2070.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2071 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [3]), 
            .O(n56814));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2071.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_2173_14_lut (.I0(GND_net), .I1(n3223), 
            .I2(VCC_net), .I3(n50107), .O(n3290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15470_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n22726), .I3(GND_net), .O(n29478));   // verilog/coms.v(130[12] 305[6])
    defparam i15470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53216_1_lut (.I0(n1554), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n68902));
    defparam i53216_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_2173_14 (.CI(n50107), .I0(n3223), 
            .I1(VCC_net), .CO(n50108));
    SB_LUT4 i53365_1_lut (.I0(n1455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69051));
    defparam i53365_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR delay_counter__i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n27698), 
            .D(n1239), .R(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    SB_LUT4 i53346_1_lut (.I0(n1356), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69032));
    defparam i53346_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53379_1_lut (.I0(n1158), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69065));
    defparam i53379_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_2173_13_lut (.I0(GND_net), .I1(n3224), 
            .I2(VCC_net), .I3(n50106), .O(n3291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_13 (.CI(n50106), .I0(n3224), 
            .I1(VCC_net), .CO(n50107));
    SB_LUT4 i53392_1_lut (.I0(n1059), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n69078));
    defparam i53392_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_add_2173_12_lut (.I0(GND_net), .I1(n3225), 
            .I2(VCC_net), .I3(n50105), .O(n3292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_12 (.CI(n50105), .I0(n3225), 
            .I1(VCC_net), .CO(n50106));
    SB_LUT4 encoder0_position_30__I_0_add_2173_11_lut (.I0(GND_net), .I1(n3226), 
            .I2(VCC_net), .I3(n50104), .O(n3293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_11 (.CI(n50104), .I0(n3226), 
            .I1(VCC_net), .CO(n50105));
    SB_LUT4 encoder0_position_30__I_0_add_2173_10_lut (.I0(GND_net), .I1(n3227), 
            .I2(VCC_net), .I3(n50103), .O(n3294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_10 (.CI(n50103), .I0(n3227), 
            .I1(VCC_net), .CO(n50104));
    SB_LUT4 encoder0_position_30__I_0_add_2173_9_lut (.I0(GND_net), .I1(n3228), 
            .I2(VCC_net), .I3(n50102), .O(n3295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_2072 (.I0(n1926), .I1(n1927), .I2(n1928), .I3(n1925), 
            .O(n61012));
    defparam i1_4_lut_adj_2072.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_30__I_0_add_2173_9 (.CI(n50102), .I0(n3228), 
            .I1(VCC_net), .CO(n50103));
    SB_LUT4 encoder0_position_30__I_0_add_2173_8_lut (.I0(GND_net), .I1(n3229), 
            .I2(GND_net), .I3(n50101), .O(n3296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_8 (.CI(n50101), .I0(n3229), 
            .I1(GND_net), .CO(n50102));
    SB_LUT4 encoder0_position_30__I_0_add_2173_7_lut (.I0(n3298), .I1(n3230), 
            .I2(GND_net), .I3(n50100), .O(n65401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_30__I_0_add_2173_7 (.CI(n50100), .I0(n3230), 
            .I1(GND_net), .CO(n50101));
    SB_LUT4 encoder0_position_30__I_0_add_2173_6_lut (.I0(GND_net), .I1(n3231), 
            .I2(VCC_net), .I3(n50099), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_6 (.CI(n50099), .I0(n3231), 
            .I1(VCC_net), .CO(n50100));
    SB_LUT4 encoder0_position_30__I_0_add_2173_5_lut (.I0(n6_adj_5826), .I1(n3232), 
            .I2(GND_net), .I3(n50098), .O(n65412)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_5_lut.LUT_INIT = 16'hebbe;
    SB_CARRY encoder0_position_30__I_0_add_2173_5 (.CI(n50098), .I0(n3232), 
            .I1(GND_net), .CO(n50099));
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk16MHz), .D(displacement_23__N_67[23]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFFESR GHC_192 (.Q(GHC), .C(clk16MHz), .E(n27646), .D(GHC_N_391), 
            .R(n28878));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GHB_190 (.Q(GHB), .C(clk16MHz), .E(n27646), .D(GHB_N_377), 
            .R(n28878));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFFESR GHA_188 (.Q(GHA), .C(clk16MHz), .E(n27646), .D(GHA_N_355), 
            .R(n28878));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk16MHz), .D(displacement_23__N_67[22]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk16MHz), .D(displacement_23__N_67[21]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(clk16MHz), 
            .E(n7_adj_5916), .D(commutation_state_7__N_208[0]), .S(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk16MHz), .D(displacement_23__N_67[20]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFFESR GLA_189 (.Q(INLA_c_0), .C(clk16MHz), .E(n27646), .D(GLA_N_372), 
            .R(n28878));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk16MHz), .D(displacement_23__N_67[19]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk16MHz), .D(displacement_23__N_67[18]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk16MHz), .D(displacement_23__N_67[17]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk16MHz), .D(displacement_23__N_67[16]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk16MHz), .D(displacement_23__N_67[15]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk16MHz), .D(displacement_23__N_67[14]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk16MHz), .D(displacement_23__N_67[13]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk16MHz), .D(displacement_23__N_67[12]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk16MHz), .D(displacement_23__N_67[11]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk16MHz), .D(displacement_23__N_67[10]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk16MHz), .D(displacement_23__N_67[9]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk16MHz), .D(displacement_23__N_67[8]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk16MHz), .D(displacement_23__N_67[7]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk16MHz), .D(displacement_23__N_67[6]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk16MHz), .D(displacement_23__N_67[5]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk16MHz), .D(displacement_23__N_67[4]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk16MHz), .D(displacement_23__N_67[3]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk16MHz), .D(displacement_23__N_67[2]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk16MHz), .D(displacement_23__N_67[1]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(clk16MHz), .D(encoder1_position[25]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(clk16MHz), .D(encoder1_position[24]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(clk16MHz), .D(encoder1_position[23]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(clk16MHz), .D(encoder1_position[22]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(clk16MHz), .D(encoder1_position[21]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(clk16MHz), .D(encoder1_position[20]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(clk16MHz), .D(encoder1_position[19]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(clk16MHz), .D(encoder1_position[18]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(clk16MHz), .D(encoder1_position[17]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(clk16MHz), .D(encoder1_position[16]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(clk16MHz), .D(encoder1_position[15]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(clk16MHz), .D(encoder1_position[14]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(clk16MHz), .D(encoder1_position[13]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(clk16MHz), .D(encoder1_position[12]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(clk16MHz), 
           .D(encoder1_position[11]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(clk16MHz), 
           .D(encoder1_position[10]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(clk16MHz), 
           .D(encoder1_position[9]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(clk16MHz), 
           .D(encoder1_position[8]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(clk16MHz), 
           .D(encoder1_position[7]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(clk16MHz), 
           .D(encoder1_position[6]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(clk16MHz), 
           .D(encoder1_position[5]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(clk16MHz), 
           .D(encoder1_position[4]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(clk16MHz), 
           .D(encoder1_position[3]));   // verilog/TinyFPGA_B.v(320[10] 324[6])
    SB_DFFESR GLB_191 (.Q(INLB_c_0), .C(clk16MHz), .E(n27646), .D(GLB_N_386), 
            .R(n28878));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 encoder0_position_30__I_0_add_2173_4_lut (.I0(n3301), .I1(n3233), 
            .I2(VCC_net), .I3(n50097), .O(n6_adj_5826)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_4_lut.LUT_INIT = 16'h8228;
    SB_DFFESR GLC_193 (.Q(INLC_c_0), .C(clk16MHz), .E(n27646), .D(GLC_N_400), 
            .R(n28878));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    SB_LUT4 i16561_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [0]), 
            .O(n30569));   // verilog/coms.v(130[12] 305[6])
    defparam i16561_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    GND i1 (.Y(GND_net));
    SB_CARRY encoder0_position_30__I_0_add_2173_4 (.CI(n50097), .I0(n3233), 
            .I1(VCC_net), .CO(n50098));
    SB_LUT4 encoder0_position_30__I_0_add_2173_3_lut (.I0(GND_net), .I1(n957), 
            .I2(GND_net), .I3(n50096), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2173_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2173_3 (.CI(n50096), .I0(n957), 
            .I1(GND_net), .CO(n50097));
    SB_CARRY encoder0_position_30__I_0_add_2173_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(VCC_net), .CO(n50096));
    SB_LUT4 encoder0_position_30__I_0_add_2106_31_lut (.I0(n68512), .I1(n3105), 
            .I2(VCC_net), .I3(n50095), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_2106_30_lut (.I0(GND_net), .I1(n3106), 
            .I2(VCC_net), .I3(n50094), .O(n3173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_30 (.CI(n50094), .I0(n3106), 
            .I1(VCC_net), .CO(n50095));
    SB_LUT4 encoder0_position_30__I_0_add_2106_29_lut (.I0(GND_net), .I1(n3107), 
            .I2(VCC_net), .I3(n50093), .O(n3174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_29 (.CI(n50093), .I0(n3107), 
            .I1(VCC_net), .CO(n50094));
    SB_LUT4 encoder0_position_30__I_0_add_2106_28_lut (.I0(GND_net), .I1(n3108), 
            .I2(VCC_net), .I3(n50092), .O(n3175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_28 (.CI(n50092), .I0(n3108), 
            .I1(VCC_net), .CO(n50093));
    SB_LUT4 encoder0_position_30__I_0_add_2106_27_lut (.I0(GND_net), .I1(n3109), 
            .I2(VCC_net), .I3(n50091), .O(n3176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_27 (.CI(n50091), .I0(n3109), 
            .I1(VCC_net), .CO(n50092));
    SB_LUT4 encoder0_position_30__I_0_add_2106_26_lut (.I0(GND_net), .I1(n3110), 
            .I2(VCC_net), .I3(n50090), .O(n3177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n49169), .O(n1216)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_26 (.CI(n50090), .I0(n3110), 
            .I1(VCC_net), .CO(n50091));
    SB_LUT4 encoder0_position_30__I_0_add_2106_25_lut (.I0(GND_net), .I1(n3111), 
            .I2(VCC_net), .I3(n50089), .O(n3178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_25 (.CI(n50089), .I0(n3111), 
            .I1(VCC_net), .CO(n50090));
    SB_LUT4 encoder0_position_30__I_0_add_2106_24_lut (.I0(GND_net), .I1(n3112), 
            .I2(VCC_net), .I3(n50088), .O(n3179)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_24 (.CI(n50088), .I0(n3112), 
            .I1(VCC_net), .CO(n50089));
    SB_LUT4 encoder0_position_30__I_0_add_2106_23_lut (.I0(GND_net), .I1(n3113), 
            .I2(VCC_net), .I3(n50087), .O(n3180)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2073 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [4]), 
            .O(n56815));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2073.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_2106_23 (.CI(n50087), .I0(n3113), 
            .I1(VCC_net), .CO(n50088));
    SB_LUT4 encoder0_position_30__I_0_add_2106_22_lut (.I0(GND_net), .I1(n3114), 
            .I2(VCC_net), .I3(n50086), .O(n3181)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_22 (.CI(n50086), .I0(n3114), 
            .I1(VCC_net), .CO(n50087));
    SB_LUT4 encoder0_position_30__I_0_add_2106_21_lut (.I0(GND_net), .I1(n3115), 
            .I2(VCC_net), .I3(n50085), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_21 (.CI(n50085), .I0(n3115), 
            .I1(VCC_net), .CO(n50086));
    SB_CARRY add_1097_9 (.CI(n49270), .I0(GND_net), .I1(n12212), .CO(n49271));
    SB_LUT4 encoder0_position_30__I_0_add_2106_20_lut (.I0(GND_net), .I1(n3116), 
            .I2(VCC_net), .I3(n50084), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_20 (.CI(n50084), .I0(n3116), 
            .I1(VCC_net), .CO(n50085));
    SB_LUT4 add_1097_8_lut (.I0(GND_net), .I1(GND_net), .I2(n12214), .I3(n49269), 
            .O(n4922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2106_19_lut (.I0(GND_net), .I1(n3117), 
            .I2(VCC_net), .I3(n50083), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_19 (.CI(n50083), .I0(n3117), 
            .I1(VCC_net), .CO(n50084));
    SB_LUT4 encoder0_position_30__I_0_add_2106_18_lut (.I0(GND_net), .I1(n3118), 
            .I2(VCC_net), .I3(n50082), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_18 (.CI(n50082), .I0(n3118), 
            .I1(VCC_net), .CO(n50083));
    SB_LUT4 encoder0_position_30__I_0_add_2106_17_lut (.I0(GND_net), .I1(n3119), 
            .I2(VCC_net), .I3(n50081), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_17 (.CI(n50081), .I0(n3119), 
            .I1(VCC_net), .CO(n50082));
    SB_LUT4 encoder0_position_30__I_0_add_2106_16_lut (.I0(GND_net), .I1(n3120), 
            .I2(VCC_net), .I3(n50080), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_16 (.CI(n50080), .I0(n3120), 
            .I1(VCC_net), .CO(n50081));
    SB_LUT4 encoder0_position_30__I_0_add_2106_15_lut (.I0(GND_net), .I1(n3121), 
            .I2(VCC_net), .I3(n50079), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_15 (.CI(n50079), .I0(n3121), 
            .I1(VCC_net), .CO(n50080));
    SB_LUT4 encoder0_position_30__I_0_add_2106_14_lut (.I0(GND_net), .I1(n3122), 
            .I2(VCC_net), .I3(n50078), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_14 (.CI(n50078), .I0(n3122), 
            .I1(VCC_net), .CO(n50079));
    SB_CARRY add_1097_8 (.CI(n49269), .I0(GND_net), .I1(n12214), .CO(n49270));
    SB_LUT4 encoder0_position_30__I_0_add_2106_13_lut (.I0(GND_net), .I1(n3123), 
            .I2(VCC_net), .I3(n50077), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_13 (.CI(n50077), .I0(n3123), 
            .I1(VCC_net), .CO(n50078));
    SB_LUT4 encoder0_position_30__I_0_add_2106_12_lut (.I0(GND_net), .I1(n3124), 
            .I2(VCC_net), .I3(n50076), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_12 (.CI(n50076), .I0(n3124), 
            .I1(VCC_net), .CO(n50077));
    SB_LUT4 encoder0_position_30__I_0_add_2106_11_lut (.I0(GND_net), .I1(n3125), 
            .I2(VCC_net), .I3(n50075), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_11 (.CI(n50075), .I0(n3125), 
            .I1(VCC_net), .CO(n50076));
    SB_LUT4 encoder0_position_30__I_0_add_2106_10_lut (.I0(GND_net), .I1(n3126), 
            .I2(VCC_net), .I3(n50074), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_10 (.CI(n50074), .I0(n3126), 
            .I1(VCC_net), .CO(n50075));
    SB_LUT4 encoder0_position_30__I_0_add_2106_9_lut (.I0(GND_net), .I1(n3127), 
            .I2(VCC_net), .I3(n50073), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1097_7_lut (.I0(GND_net), .I1(GND_net), .I2(n12216), .I3(n49268), 
            .O(n4923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_9 (.CI(n50073), .I0(n3127), 
            .I1(VCC_net), .CO(n50074));
    SB_LUT4 encoder0_position_30__I_0_add_2106_8_lut (.I0(GND_net), .I1(n3128), 
            .I2(VCC_net), .I3(n50072), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_8 (.CI(n50072), .I0(n3128), 
            .I1(VCC_net), .CO(n50073));
    SB_LUT4 encoder0_position_30__I_0_add_2106_7_lut (.I0(GND_net), .I1(n3129), 
            .I2(GND_net), .I3(n50071), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_7 (.CI(n50071), .I0(n3129), 
            .I1(GND_net), .CO(n50072));
    SB_LUT4 encoder0_position_30__I_0_add_2106_6_lut (.I0(GND_net), .I1(n3130), 
            .I2(GND_net), .I3(n50070), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_6 (.CI(n50070), .I0(n3130), 
            .I1(GND_net), .CO(n50071));
    SB_LUT4 encoder0_position_30__I_0_add_2106_5_lut (.I0(GND_net), .I1(n3131), 
            .I2(VCC_net), .I3(n50069), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_5 (.CI(n50069), .I0(n3131), 
            .I1(VCC_net), .CO(n50070));
    SB_LUT4 encoder0_position_30__I_0_add_2106_4_lut (.I0(GND_net), .I1(n3132), 
            .I2(GND_net), .I3(n50068), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_4 (.CI(n50068), .I0(n3132), 
            .I1(GND_net), .CO(n50069));
    SB_LUT4 encoder0_position_30__I_0_add_2106_3_lut (.I0(GND_net), .I1(n3133), 
            .I2(VCC_net), .I3(n50067), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_3 (.CI(n50067), .I0(n3133), 
            .I1(VCC_net), .CO(n50068));
    SB_LUT4 encoder0_position_30__I_0_add_2106_2_lut (.I0(GND_net), .I1(n956), 
            .I2(GND_net), .I3(VCC_net), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2106_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2106_2 (.CI(VCC_net), .I0(n956), 
            .I1(GND_net), .CO(n50067));
    SB_LUT4 encoder0_position_30__I_0_add_2039_30_lut (.I0(n68551), .I1(n3006), 
            .I2(VCC_net), .I3(n50066), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_151_25 (.CI(n49169), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n49170));
    SB_LUT4 encoder0_position_30__I_0_add_2039_29_lut (.I0(GND_net), .I1(n3007), 
            .I2(VCC_net), .I3(n50065), .O(n3074)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1097_7 (.CI(n49268), .I0(GND_net), .I1(n12216), .CO(n49269));
    SB_CARRY encoder0_position_30__I_0_add_2039_29 (.CI(n50065), .I0(n3007), 
            .I1(VCC_net), .CO(n50066));
    SB_LUT4 encoder0_position_30__I_0_add_2039_28_lut (.I0(GND_net), .I1(n3008), 
            .I2(VCC_net), .I3(n50064), .O(n3075)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_28 (.CI(n50064), .I0(n3008), 
            .I1(VCC_net), .CO(n50065));
    SB_LUT4 encoder0_position_30__I_0_add_2039_27_lut (.I0(GND_net), .I1(n3009), 
            .I2(VCC_net), .I3(n50063), .O(n3076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n49168), .O(n1217)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_27 (.CI(n50063), .I0(n3009), 
            .I1(VCC_net), .CO(n50064));
    SB_LUT4 encoder0_position_30__I_0_add_2039_26_lut (.I0(GND_net), .I1(n3010), 
            .I2(VCC_net), .I3(n50062), .O(n3077)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_26 (.CI(n50062), .I0(n3010), 
            .I1(VCC_net), .CO(n50063));
    SB_LUT4 encoder0_position_30__I_0_add_2039_25_lut (.I0(GND_net), .I1(n3011), 
            .I2(VCC_net), .I3(n50061), .O(n3078)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_25 (.CI(n50061), .I0(n3011), 
            .I1(VCC_net), .CO(n50062));
    SB_CARRY add_151_24 (.CI(n49168), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n49169));
    SB_LUT4 encoder0_position_30__I_0_add_2039_24_lut (.I0(GND_net), .I1(n3012), 
            .I2(VCC_net), .I3(n50060), .O(n3079)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_24 (.CI(n50060), .I0(n3012), 
            .I1(VCC_net), .CO(n50061));
    SB_LUT4 encoder0_position_30__I_0_add_2039_23_lut (.I0(GND_net), .I1(n3013), 
            .I2(VCC_net), .I3(n50059), .O(n3080)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_23 (.CI(n50059), .I0(n3013), 
            .I1(VCC_net), .CO(n50060));
    SB_LUT4 encoder0_position_30__I_0_add_2039_22_lut (.I0(GND_net), .I1(n3014), 
            .I2(VCC_net), .I3(n50058), .O(n3081)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_22 (.CI(n50058), .I0(n3014), 
            .I1(VCC_net), .CO(n50059));
    SB_LUT4 encoder0_position_30__I_0_add_2039_21_lut (.I0(GND_net), .I1(n3015), 
            .I2(VCC_net), .I3(n50057), .O(n3082)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_21 (.CI(n50057), .I0(n3015), 
            .I1(VCC_net), .CO(n50058));
    SB_LUT4 encoder0_position_30__I_0_add_2039_20_lut (.I0(GND_net), .I1(n3016), 
            .I2(VCC_net), .I3(n50056), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_20 (.CI(n50056), .I0(n3016), 
            .I1(VCC_net), .CO(n50057));
    SB_LUT4 encoder0_position_30__I_0_add_2039_19_lut (.I0(GND_net), .I1(n3017), 
            .I2(VCC_net), .I3(n50055), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_19 (.CI(n50055), .I0(n3017), 
            .I1(VCC_net), .CO(n50056));
    SB_LUT4 i15472_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n22726), .I3(GND_net), .O(n29480));   // verilog/coms.v(130[12] 305[6])
    defparam i15472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2074 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [5]), 
            .O(n56816));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2074.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_2039_18_lut (.I0(GND_net), .I1(n3018), 
            .I2(VCC_net), .I3(n50054), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_18 (.CI(n50054), .I0(n3018), 
            .I1(VCC_net), .CO(n50055));
    SB_LUT4 encoder0_position_30__I_0_add_2039_17_lut (.I0(GND_net), .I1(n3019), 
            .I2(VCC_net), .I3(n50053), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_17 (.CI(n50053), .I0(n3019), 
            .I1(VCC_net), .CO(n50054));
    SB_LUT4 encoder0_position_30__I_0_add_2039_16_lut (.I0(GND_net), .I1(n3020), 
            .I2(VCC_net), .I3(n50052), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_16 (.CI(n50052), .I0(n3020), 
            .I1(VCC_net), .CO(n50053));
    SB_LUT4 encoder0_position_30__I_0_add_2039_15_lut (.I0(GND_net), .I1(n3021), 
            .I2(VCC_net), .I3(n50051), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_15 (.CI(n50051), .I0(n3021), 
            .I1(VCC_net), .CO(n50052));
    SB_LUT4 encoder0_position_30__I_0_add_2039_14_lut (.I0(GND_net), .I1(n3022), 
            .I2(VCC_net), .I3(n50050), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_14 (.CI(n50050), .I0(n3022), 
            .I1(VCC_net), .CO(n50051));
    SB_LUT4 encoder0_position_30__I_0_add_2039_13_lut (.I0(GND_net), .I1(n3023), 
            .I2(VCC_net), .I3(n50049), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_13 (.CI(n50049), .I0(n3023), 
            .I1(VCC_net), .CO(n50050));
    SB_LUT4 add_1097_6_lut (.I0(GND_net), .I1(GND_net), .I2(n12218), .I3(n49267), 
            .O(n4924)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_12_lut (.I0(GND_net), .I1(n3024), 
            .I2(VCC_net), .I3(n50048), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_12 (.CI(n50048), .I0(n3024), 
            .I1(VCC_net), .CO(n50049));
    SB_LUT4 encoder0_position_30__I_0_add_2039_11_lut (.I0(GND_net), .I1(n3025), 
            .I2(VCC_net), .I3(n50047), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_11 (.CI(n50047), .I0(n3025), 
            .I1(VCC_net), .CO(n50048));
    SB_LUT4 encoder0_position_30__I_0_add_2039_10_lut (.I0(GND_net), .I1(n3026), 
            .I2(VCC_net), .I3(n50046), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_10 (.CI(n50046), .I0(n3026), 
            .I1(VCC_net), .CO(n50047));
    SB_LUT4 add_151_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n49167), .O(n1218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_2039_9_lut (.I0(GND_net), .I1(n3027), 
            .I2(VCC_net), .I3(n50045), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1097_6 (.CI(n49267), .I0(GND_net), .I1(n12218), .CO(n49268));
    SB_CARRY encoder0_position_30__I_0_add_2039_9 (.CI(n50045), .I0(n3027), 
            .I1(VCC_net), .CO(n50046));
    SB_LUT4 encoder0_position_30__I_0_add_2039_8_lut (.I0(GND_net), .I1(n3028), 
            .I2(VCC_net), .I3(n50044), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_8 (.CI(n50044), .I0(n3028), 
            .I1(VCC_net), .CO(n50045));
    SB_LUT4 encoder0_position_30__I_0_add_2039_7_lut (.I0(GND_net), .I1(n3029), 
            .I2(GND_net), .I3(n50043), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_7 (.CI(n50043), .I0(n3029), 
            .I1(GND_net), .CO(n50044));
    SB_LUT4 encoder0_position_30__I_0_add_2039_6_lut (.I0(GND_net), .I1(n3030), 
            .I2(GND_net), .I3(n50042), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2075 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [6]), 
            .O(n56817));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2075.LUT_INIT = 16'h2300;
    SB_LUT4 add_1097_5_lut (.I0(GND_net), .I1(GND_net), .I2(n12220), .I3(n49266), 
            .O(n4925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_6 (.CI(n50042), .I0(n3030), 
            .I1(GND_net), .CO(n50043));
    SB_LUT4 encoder0_position_30__I_0_add_2039_5_lut (.I0(GND_net), .I1(n3031), 
            .I2(VCC_net), .I3(n50041), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_5 (.CI(n50041), .I0(n3031), 
            .I1(VCC_net), .CO(n50042));
    SB_LUT4 encoder0_position_30__I_0_add_2039_4_lut (.I0(GND_net), .I1(n3032), 
            .I2(GND_net), .I3(n50040), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_4 (.CI(n50040), .I0(n3032), 
            .I1(GND_net), .CO(n50041));
    SB_LUT4 encoder0_position_30__I_0_add_2039_3_lut (.I0(GND_net), .I1(n3033), 
            .I2(VCC_net), .I3(n50039), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1097_5 (.CI(n49266), .I0(GND_net), .I1(n12220), .CO(n49267));
    SB_CARRY encoder0_position_30__I_0_add_2039_3 (.CI(n50039), .I0(n3033), 
            .I1(VCC_net), .CO(n50040));
    SB_LUT4 encoder0_position_30__I_0_add_2039_2_lut (.I0(GND_net), .I1(n955), 
            .I2(GND_net), .I3(VCC_net), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_2039_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_2039_2 (.CI(VCC_net), .I0(n955), 
            .I1(GND_net), .CO(n50039));
    SB_LUT4 encoder0_position_30__I_0_add_1972_29_lut (.I0(GND_net), .I1(n2907), 
            .I2(VCC_net), .I3(n50038), .O(n2974)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_28_lut (.I0(GND_net), .I1(n2908), 
            .I2(VCC_net), .I3(n50037), .O(n2975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_28 (.CI(n50037), .I0(n2908), 
            .I1(VCC_net), .CO(n50038));
    SB_LUT4 encoder0_position_30__I_0_add_1972_27_lut (.I0(GND_net), .I1(n2909), 
            .I2(VCC_net), .I3(n50036), .O(n2976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_27 (.CI(n50036), .I0(n2909), 
            .I1(VCC_net), .CO(n50037));
    SB_LUT4 encoder0_position_30__I_0_add_1972_26_lut (.I0(GND_net), .I1(n2910), 
            .I2(VCC_net), .I3(n50035), .O(n2977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_23 (.CI(n49167), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n49168));
    SB_CARRY encoder0_position_30__I_0_add_1972_26 (.CI(n50035), .I0(n2910), 
            .I1(VCC_net), .CO(n50036));
    SB_LUT4 encoder0_position_30__I_0_add_1972_25_lut (.I0(GND_net), .I1(n2911), 
            .I2(VCC_net), .I3(n50034), .O(n2978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_25 (.CI(n50034), .I0(n2911), 
            .I1(VCC_net), .CO(n50035));
    SB_LUT4 add_1097_4_lut (.I0(GND_net), .I1(GND_net), .I2(n12222), .I3(n49265), 
            .O(n4926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_10 (.CI(n49154), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n49155));
    SB_LUT4 encoder0_position_30__I_0_add_1972_24_lut (.I0(GND_net), .I1(n2912), 
            .I2(VCC_net), .I3(n50033), .O(n2979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2076 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [7]), 
            .O(n56818));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2076.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1972_24 (.CI(n50033), .I0(n2912), 
            .I1(VCC_net), .CO(n50034));
    SB_LUT4 encoder0_position_30__I_0_add_1168_17_lut (.I0(n68943), .I1(n1719), 
            .I2(VCC_net), .I3(n49681), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1168_16_lut (.I0(GND_net), .I1(n1720), 
            .I2(VCC_net), .I3(n49680), .O(n1787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n49166), .O(n1219)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_23_lut (.I0(GND_net), .I1(n2913), 
            .I2(VCC_net), .I3(n50032), .O(n2980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_16 (.CI(n49680), .I0(n1720), 
            .I1(VCC_net), .CO(n49681));
    SB_CARRY encoder0_position_30__I_0_add_1972_23 (.CI(n50032), .I0(n2913), 
            .I1(VCC_net), .CO(n50033));
    SB_LUT4 encoder0_position_30__I_0_add_1972_22_lut (.I0(GND_net), .I1(n2914), 
            .I2(VCC_net), .I3(n50031), .O(n2981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_22 (.CI(n50031), .I0(n2914), 
            .I1(VCC_net), .CO(n50032));
    SB_LUT4 encoder0_position_30__I_0_add_1972_21_lut (.I0(GND_net), .I1(n2915), 
            .I2(VCC_net), .I3(n50030), .O(n2982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_15_lut (.I0(GND_net), .I1(n1721), 
            .I2(VCC_net), .I3(n49679), .O(n1788_adj_5804)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_21 (.CI(n50030), .I0(n2915), 
            .I1(VCC_net), .CO(n50031));
    SB_LUT4 encoder0_position_30__I_0_add_1972_20_lut (.I0(GND_net), .I1(n2916), 
            .I2(VCC_net), .I3(n50029), .O(n2983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1097_4 (.CI(n49265), .I0(GND_net), .I1(n12222), .CO(n49266));
    SB_CARRY encoder0_position_30__I_0_add_1972_20 (.CI(n50029), .I0(n2916), 
            .I1(VCC_net), .CO(n50030));
    SB_LUT4 encoder0_position_30__I_0_add_1972_19_lut (.I0(GND_net), .I1(n2917), 
            .I2(VCC_net), .I3(n50028), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_15 (.CI(n49679), .I0(n1721), 
            .I1(VCC_net), .CO(n49680));
    SB_CARRY encoder0_position_30__I_0_add_1972_19 (.CI(n50028), .I0(n2917), 
            .I1(VCC_net), .CO(n50029));
    SB_LUT4 encoder0_position_30__I_0_add_1972_18_lut (.I0(GND_net), .I1(n2918), 
            .I2(VCC_net), .I3(n50027), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_14_lut (.I0(GND_net), .I1(n1722), 
            .I2(VCC_net), .I3(n49678), .O(n1789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_14 (.CI(n49678), .I0(n1722), 
            .I1(VCC_net), .CO(n49679));
    SB_CARRY encoder0_position_30__I_0_add_1972_18 (.CI(n50027), .I0(n2918), 
            .I1(VCC_net), .CO(n50028));
    SB_LUT4 encoder0_position_30__I_0_add_1168_13_lut (.I0(GND_net), .I1(n1723), 
            .I2(VCC_net), .I3(n49677), .O(n1790_adj_5805)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_17_lut (.I0(GND_net), .I1(n2919), 
            .I2(VCC_net), .I3(n50026), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_17 (.CI(n50026), .I0(n2919), 
            .I1(VCC_net), .CO(n50027));
    SB_LUT4 encoder0_position_30__I_0_add_1972_16_lut (.I0(GND_net), .I1(n2920), 
            .I2(VCC_net), .I3(n50025), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_16 (.CI(n50025), .I0(n2920), 
            .I1(VCC_net), .CO(n50026));
    SB_LUT4 encoder0_position_30__I_0_add_1972_15_lut (.I0(GND_net), .I1(n2921), 
            .I2(VCC_net), .I3(n50024), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_15 (.CI(n50024), .I0(n2921), 
            .I1(VCC_net), .CO(n50025));
    SB_LUT4 encoder0_position_30__I_0_add_1972_14_lut (.I0(GND_net), .I1(n2922), 
            .I2(VCC_net), .I3(n50023), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_14 (.CI(n50023), .I0(n2922), 
            .I1(VCC_net), .CO(n50024));
    SB_LUT4 encoder0_position_30__I_0_add_1972_13_lut (.I0(GND_net), .I1(n2923), 
            .I2(VCC_net), .I3(n50022), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_13 (.CI(n49677), .I0(n1723), 
            .I1(VCC_net), .CO(n49678));
    SB_LUT4 encoder0_position_30__I_0_add_1168_12_lut (.I0(GND_net), .I1(n1724), 
            .I2(VCC_net), .I3(n49676), .O(n1791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_13 (.CI(n50022), .I0(n2923), 
            .I1(VCC_net), .CO(n50023));
    SB_CARRY encoder0_position_30__I_0_add_1168_12 (.CI(n49676), .I0(n1724), 
            .I1(VCC_net), .CO(n49677));
    SB_LUT4 encoder0_position_30__I_0_add_1168_11_lut (.I0(GND_net), .I1(n1725), 
            .I2(VCC_net), .I3(n49675), .O(n1792_adj_5806)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1097_3_lut (.I0(GND_net), .I1(GND_net), .I2(n12224), .I3(n49264), 
            .O(n4927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1097_3 (.CI(n49264), .I0(GND_net), .I1(n12224), .CO(n49265));
    SB_LUT4 encoder0_position_30__I_0_add_699_10_lut (.I0(GND_net), .I1(n1026), 
            .I2(VCC_net), .I3(n49474), .O(n1093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_11 (.CI(n49675), .I0(n1725), 
            .I1(VCC_net), .CO(n49676));
    SB_LUT4 encoder0_position_30__I_0_add_1168_10_lut (.I0(GND_net), .I1(n1726), 
            .I2(VCC_net), .I3(n49674), .O(n1793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_10 (.CI(n49674), .I0(n1726), 
            .I1(VCC_net), .CO(n49675));
    SB_LUT4 encoder0_position_30__I_0_add_1168_9_lut (.I0(GND_net), .I1(n1727), 
            .I2(VCC_net), .I3(n49673), .O(n1794_adj_5807)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_9_lut (.I0(GND_net), .I1(n1027), 
            .I2(VCC_net), .I3(n49473), .O(n1094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_9 (.CI(n49673), .I0(n1727), 
            .I1(VCC_net), .CO(n49674));
    SB_LUT4 encoder0_position_30__I_0_add_1972_12_lut (.I0(GND_net), .I1(n2924), 
            .I2(VCC_net), .I3(n50021), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_12 (.CI(n50021), .I0(n2924), 
            .I1(VCC_net), .CO(n50022));
    SB_CARRY encoder0_position_30__I_0_add_699_9 (.CI(n49473), .I0(n1027), 
            .I1(VCC_net), .CO(n49474));
    SB_CARRY add_151_22 (.CI(n49166), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n49167));
    SB_LUT4 encoder0_position_30__I_0_add_699_8_lut (.I0(GND_net), .I1(n1028), 
            .I2(VCC_net), .I3(n49472), .O(n1095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_8_lut (.I0(GND_net), .I1(n1728), 
            .I2(VCC_net), .I3(n49672), .O(n1795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1972_11_lut (.I0(GND_net), .I1(n2925), 
            .I2(VCC_net), .I3(n50020), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_8 (.CI(n49672), .I0(n1728), 
            .I1(VCC_net), .CO(n49673));
    SB_LUT4 add_1097_2_lut (.I0(GND_net), .I1(GND_net), .I2(n11642), .I3(VCC_net), 
            .O(n4928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1097_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_8 (.CI(n49472), .I0(n1028), 
            .I1(VCC_net), .CO(n49473));
    SB_CARRY encoder0_position_30__I_0_add_1972_11 (.CI(n50020), .I0(n2925), 
            .I1(VCC_net), .CO(n50021));
    SB_LUT4 encoder0_position_30__I_0_add_699_7_lut (.I0(GND_net), .I1(n1029), 
            .I2(GND_net), .I3(n49471), .O(n1096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_7_lut (.I0(GND_net), .I1(n1729), 
            .I2(GND_net), .I3(n49671), .O(n1796_adj_5808)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_7 (.CI(n49471), .I0(n1029), 
            .I1(GND_net), .CO(n49472));
    SB_LUT4 encoder0_position_30__I_0_add_1972_10_lut (.I0(GND_net), .I1(n2926), 
            .I2(VCC_net), .I3(n50019), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_10 (.CI(n50019), .I0(n2926), 
            .I1(VCC_net), .CO(n50020));
    SB_LUT4 encoder0_position_30__I_0_add_1972_9_lut (.I0(GND_net), .I1(n2927), 
            .I2(VCC_net), .I3(n50018), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_7 (.CI(n49671), .I0(n1729), 
            .I1(GND_net), .CO(n49672));
    SB_LUT4 encoder0_position_30__I_0_add_699_6_lut (.I0(GND_net), .I1(n1030), 
            .I2(GND_net), .I3(n49470), .O(n1097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_9 (.CI(n50018), .I0(n2927), 
            .I1(VCC_net), .CO(n50019));
    SB_LUT4 encoder0_position_30__I_0_add_1972_8_lut (.I0(GND_net), .I1(n2928), 
            .I2(VCC_net), .I3(n50017), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n49147), .O(n1238)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_8 (.CI(n50017), .I0(n2928), 
            .I1(VCC_net), .CO(n50018));
    SB_LUT4 encoder0_position_30__I_0_add_1972_7_lut (.I0(GND_net), .I1(n2929), 
            .I2(GND_net), .I3(n50016), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_6_lut (.I0(GND_net), .I1(n1730), 
            .I2(GND_net), .I3(n49670), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_6 (.CI(n49470), .I0(n1030), 
            .I1(GND_net), .CO(n49471));
    SB_CARRY encoder0_position_30__I_0_add_1168_6 (.CI(n49670), .I0(n1730), 
            .I1(GND_net), .CO(n49671));
    SB_LUT4 encoder0_position_30__I_0_add_699_5_lut (.I0(GND_net), .I1(n1031), 
            .I2(VCC_net), .I3(n49469), .O(n1098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_7 (.CI(n50016), .I0(n2929), 
            .I1(GND_net), .CO(n50017));
    SB_CARRY add_1097_2 (.CI(VCC_net), .I0(GND_net), .I1(n11642), .CO(n49264));
    SB_LUT4 encoder0_position_30__I_0_add_1972_6_lut (.I0(GND_net), .I1(n2930), 
            .I2(GND_net), .I3(n50015), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_6 (.CI(n50015), .I0(n2930), 
            .I1(GND_net), .CO(n50016));
    SB_LUT4 encoder0_position_30__I_0_add_1168_5_lut (.I0(GND_net), .I1(n1731), 
            .I2(VCC_net), .I3(n49669), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_5 (.CI(n49669), .I0(n1731), 
            .I1(VCC_net), .CO(n49670));
    SB_LUT4 encoder0_position_30__I_0_add_1972_5_lut (.I0(GND_net), .I1(n2931), 
            .I2(VCC_net), .I3(n50014), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1168_4_lut (.I0(GND_net), .I1(n1732), 
            .I2(GND_net), .I3(n49668), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_5 (.CI(n49469), .I0(n1031), 
            .I1(VCC_net), .CO(n49470));
    SB_CARRY encoder0_position_30__I_0_add_1972_5 (.CI(n50014), .I0(n2931), 
            .I1(VCC_net), .CO(n50015));
    SB_LUT4 encoder0_position_30__I_0_add_1972_4_lut (.I0(GND_net), .I1(n2932), 
            .I2(GND_net), .I3(n50013), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_4_lut (.I0(GND_net), .I1(n1032), 
            .I2(GND_net), .I3(n49468), .O(n1099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_4 (.CI(n49468), .I0(n1032), 
            .I1(GND_net), .CO(n49469));
    SB_CARRY encoder0_position_30__I_0_add_1972_4 (.CI(n50013), .I0(n2932), 
            .I1(GND_net), .CO(n50014));
    SB_CARRY encoder0_position_30__I_0_add_1168_4 (.CI(n49668), .I0(n1732), 
            .I1(GND_net), .CO(n49669));
    SB_LUT4 encoder0_position_30__I_0_add_1972_3_lut (.I0(GND_net), .I1(n2933), 
            .I2(VCC_net), .I3(n50012), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n49153), .O(n1232)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_699_3_lut (.I0(GND_net), .I1(n1033), 
            .I2(VCC_net), .I3(n49467), .O(n1100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_3 (.CI(n49467), .I0(n1033), 
            .I1(VCC_net), .CO(n49468));
    SB_CARRY encoder0_position_30__I_0_add_1972_3 (.CI(n50012), .I0(n2933), 
            .I1(VCC_net), .CO(n50013));
    SB_LUT4 encoder0_position_30__I_0_add_1168_3_lut (.I0(GND_net), .I1(n1733), 
            .I2(VCC_net), .I3(n49667), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1168_3 (.CI(n49667), .I0(n1733), 
            .I1(VCC_net), .CO(n49668));
    SB_LUT4 encoder0_position_30__I_0_add_1972_2_lut (.I0(GND_net), .I1(n954), 
            .I2(GND_net), .I3(VCC_net), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1972_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1972_2 (.CI(VCC_net), .I0(n954), 
            .I1(GND_net), .CO(n50012));
    SB_LUT4 encoder0_position_30__I_0_add_699_2_lut (.I0(GND_net), .I1(n521), 
            .I2(GND_net), .I3(VCC_net), .O(n1101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_699_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_699_2 (.CI(VCC_net), .I0(n521), 
            .I1(GND_net), .CO(n49467));
    SB_LUT4 encoder0_position_30__I_0_add_1168_2_lut (.I0(GND_net), .I1(n942), 
            .I2(GND_net), .I3(VCC_net), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1168_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_28_lut (.I0(n68643), .I1(n2808), 
            .I2(VCC_net), .I3(n50011), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1905_27_lut (.I0(GND_net), .I1(n2809), 
            .I2(VCC_net), .I3(n50010), .O(n2876)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_27 (.CI(n50010), .I0(n2809), 
            .I1(VCC_net), .CO(n50011));
    SB_LUT4 encoder0_position_30__I_0_add_1905_26_lut (.I0(GND_net), .I1(n2810), 
            .I2(VCC_net), .I3(n50009), .O(n2877)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_26 (.CI(n50009), .I0(n2810), 
            .I1(VCC_net), .CO(n50010));
    SB_CARRY encoder0_position_30__I_0_add_1168_2 (.CI(VCC_net), .I0(n942), 
            .I1(GND_net), .CO(n49667));
    SB_LUT4 encoder0_position_30__I_0_add_632_9_lut (.I0(n960), .I1(n927), 
            .I2(VCC_net), .I3(n49466), .O(n1026)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1905_25_lut (.I0(GND_net), .I1(n2811), 
            .I2(VCC_net), .I3(n50008), .O(n2878)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_632_8_lut (.I0(GND_net), .I1(n928), 
            .I2(VCC_net), .I3(n49465), .O(n995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n49165), .O(n1220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_25 (.CI(n50008), .I0(n2811), 
            .I1(VCC_net), .CO(n50009));
    SB_LUT4 encoder0_position_30__I_0_add_1905_24_lut (.I0(GND_net), .I1(n2812), 
            .I2(VCC_net), .I3(n50007), .O(n2879)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_24 (.CI(n50007), .I0(n2812), 
            .I1(VCC_net), .CO(n50008));
    SB_LUT4 encoder0_position_30__I_0_add_1905_23_lut (.I0(GND_net), .I1(n2813), 
            .I2(VCC_net), .I3(n50006), .O(n2880)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_8 (.CI(n49465), .I0(n928), 
            .I1(VCC_net), .CO(n49466));
    SB_CARRY encoder0_position_30__I_0_add_1905_23 (.CI(n50006), .I0(n2813), 
            .I1(VCC_net), .CO(n50007));
    SB_LUT4 encoder0_position_30__I_0_add_1905_22_lut (.I0(GND_net), .I1(n2814), 
            .I2(VCC_net), .I3(n50005), .O(n2881)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_632_7_lut (.I0(GND_net), .I1(n929), 
            .I2(GND_net), .I3(n49464), .O(n996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_22 (.CI(n50005), .I0(n2814), 
            .I1(VCC_net), .CO(n50006));
    SB_CARRY add_151_21 (.CI(n49165), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n49166));
    SB_LUT4 encoder0_position_30__I_0_add_1905_21_lut (.I0(GND_net), .I1(n2815), 
            .I2(VCC_net), .I3(n50004), .O(n2882)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_21 (.CI(n50004), .I0(n2815), 
            .I1(VCC_net), .CO(n50005));
    SB_CARRY encoder0_position_30__I_0_add_632_7 (.CI(n49464), .I0(n929), 
            .I1(GND_net), .CO(n49465));
    SB_LUT4 encoder0_position_30__I_0_add_632_6_lut (.I0(GND_net), .I1(n930), 
            .I2(GND_net), .I3(n49463), .O(n997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_20_lut (.I0(GND_net), .I1(n2816), 
            .I2(VCC_net), .I3(n50003), .O(n2883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_20 (.CI(n50003), .I0(n2816), 
            .I1(VCC_net), .CO(n50004));
    SB_CARRY encoder0_position_30__I_0_add_632_6 (.CI(n49463), .I0(n930), 
            .I1(GND_net), .CO(n49464));
    SB_LUT4 encoder0_position_30__I_0_add_1905_19_lut (.I0(GND_net), .I1(n2817), 
            .I2(VCC_net), .I3(n50002), .O(n2884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_632_5_lut (.I0(GND_net), .I1(n931), 
            .I2(VCC_net), .I3(n49462), .O(n998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_19 (.CI(n50002), .I0(n2817), 
            .I1(VCC_net), .CO(n50003));
    SB_LUT4 encoder0_position_30__I_0_add_1905_18_lut (.I0(GND_net), .I1(n2818), 
            .I2(VCC_net), .I3(n50001), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_5 (.CI(n49462), .I0(n931), 
            .I1(VCC_net), .CO(n49463));
    SB_LUT4 encoder0_position_30__I_0_add_632_4_lut (.I0(GND_net), .I1(n932), 
            .I2(GND_net), .I3(n49461), .O(n999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_18 (.CI(n50001), .I0(n2818), 
            .I1(VCC_net), .CO(n50002));
    SB_CARRY encoder0_position_30__I_0_add_632_4 (.CI(n49461), .I0(n932), 
            .I1(GND_net), .CO(n49462));
    SB_LUT4 encoder0_position_30__I_0_add_1905_17_lut (.I0(GND_net), .I1(n2819), 
            .I2(VCC_net), .I3(n50000), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_17 (.CI(n50000), .I0(n2819), 
            .I1(VCC_net), .CO(n50001));
    SB_LUT4 encoder0_position_30__I_0_add_632_3_lut (.I0(GND_net), .I1(n933), 
            .I2(VCC_net), .I3(n49460), .O(n1000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_16_lut (.I0(GND_net), .I1(n2820_adj_5813), 
            .I2(VCC_net), .I3(n49999), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_16 (.CI(n49999), .I0(n2820_adj_5813), 
            .I1(VCC_net), .CO(n50000));
    SB_CARRY encoder0_position_30__I_0_add_632_3 (.CI(n49460), .I0(n933), 
            .I1(VCC_net), .CO(n49461));
    SB_LUT4 encoder0_position_30__I_0_add_632_2_lut (.I0(GND_net), .I1(n520), 
            .I2(GND_net), .I3(VCC_net), .O(n1001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_632_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_15_lut (.I0(GND_net), .I1(n2821), 
            .I2(VCC_net), .I3(n49998), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_632_2 (.CI(VCC_net), .I0(n520), 
            .I1(GND_net), .CO(n49460));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2077 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [0]), 
            .O(n56819));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2077.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_565_8_lut (.I0(n861), .I1(n828), 
            .I2(VCC_net), .I3(n49459), .O(n927)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_565_7_lut (.I0(GND_net), .I1(n829), 
            .I2(GND_net), .I3(n49458), .O(n896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_15 (.CI(n49998), .I0(n2821), 
            .I1(VCC_net), .CO(n49999));
    SB_LUT4 encoder0_position_30__I_0_add_1101_16_lut (.I0(n68923), .I1(n1620), 
            .I2(VCC_net), .I3(n49648), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1101_15_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n49647), .O(n1688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_15 (.CI(n49647), .I0(n1621), 
            .I1(VCC_net), .CO(n49648));
    SB_LUT4 encoder0_position_30__I_0_add_1101_14_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n49646), .O(n1689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_7 (.CI(n49458), .I0(n829), 
            .I1(GND_net), .CO(n49459));
    SB_LUT4 encoder0_position_30__I_0_add_1905_14_lut (.I0(GND_net), .I1(n2822), 
            .I2(VCC_net), .I3(n49997), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_14 (.CI(n49997), .I0(n2822), 
            .I1(VCC_net), .CO(n49998));
    SB_LUT4 encoder0_position_30__I_0_add_565_6_lut (.I0(GND_net), .I1(n830), 
            .I2(GND_net), .I3(n49457), .O(n897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_6 (.CI(n49457), .I0(n830), 
            .I1(GND_net), .CO(n49458));
    SB_LUT4 encoder0_position_30__I_0_add_565_5_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n49456), .O(n898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_14 (.CI(n49646), .I0(n1622), 
            .I1(VCC_net), .CO(n49647));
    SB_CARRY encoder0_position_30__I_0_add_565_5 (.CI(n49456), .I0(n831), 
            .I1(VCC_net), .CO(n49457));
    SB_LUT4 encoder0_position_30__I_0_add_1101_13_lut (.I0(GND_net), .I1(n1623), 
            .I2(VCC_net), .I3(n49645), .O(n1690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_13 (.CI(n49645), .I0(n1623), 
            .I1(VCC_net), .CO(n49646));
    SB_LUT4 add_151_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n49164), .O(n1221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_565_4_lut (.I0(GND_net), .I1(n832), 
            .I2(GND_net), .I3(n49455), .O(n899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_13_lut (.I0(GND_net), .I1(n2823), 
            .I2(VCC_net), .I3(n49996), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_4 (.CI(n49455), .I0(n832), 
            .I1(GND_net), .CO(n49456));
    SB_LUT4 encoder0_position_30__I_0_add_1101_12_lut (.I0(GND_net), .I1(n1624), 
            .I2(VCC_net), .I3(n49644), .O(n1691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_13 (.CI(n49996), .I0(n2823), 
            .I1(VCC_net), .CO(n49997));
    SB_CARRY encoder0_position_30__I_0_add_1101_12 (.CI(n49644), .I0(n1624), 
            .I1(VCC_net), .CO(n49645));
    SB_LUT4 encoder0_position_30__I_0_add_1905_12_lut (.I0(GND_net), .I1(n2824), 
            .I2(VCC_net), .I3(n49995), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_11_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n49643), .O(n1692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_565_3_lut (.I0(GND_net), .I1(n833), 
            .I2(VCC_net), .I3(n49454), .O(n900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_11 (.CI(n49643), .I0(n1625), 
            .I1(VCC_net), .CO(n49644));
    SB_LUT4 encoder0_position_30__I_0_add_1101_10_lut (.I0(GND_net), .I1(n1626), 
            .I2(VCC_net), .I3(n49642), .O(n1693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_10 (.CI(n49642), .I0(n1626), 
            .I1(VCC_net), .CO(n49643));
    SB_LUT4 encoder0_position_30__I_0_add_1101_9_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n49641), .O(n1694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_565_3 (.CI(n49454), .I0(n833), 
            .I1(VCC_net), .CO(n49455));
    SB_CARRY encoder0_position_30__I_0_add_1905_12 (.CI(n49995), .I0(n2824), 
            .I1(VCC_net), .CO(n49996));
    SB_LUT4 encoder0_position_30__I_0_add_1905_11_lut (.I0(GND_net), .I1(n2825), 
            .I2(VCC_net), .I3(n49994), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_565_2_lut (.I0(GND_net), .I1(n519), 
            .I2(GND_net), .I3(VCC_net), .O(n901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_9 (.CI(n49641), .I0(n1627), 
            .I1(VCC_net), .CO(n49642));
    SB_CARRY encoder0_position_30__I_0_add_1905_11 (.CI(n49994), .I0(n2825), 
            .I1(VCC_net), .CO(n49995));
    SB_LUT4 encoder0_position_30__I_0_add_1101_8_lut (.I0(GND_net), .I1(n1628), 
            .I2(VCC_net), .I3(n49640), .O(n1695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_10_lut (.I0(GND_net), .I1(n2826), 
            .I2(VCC_net), .I3(n49993), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_10 (.CI(n49993), .I0(n2826), 
            .I1(VCC_net), .CO(n49994));
    SB_LUT4 encoder0_position_30__I_0_add_1905_9_lut (.I0(GND_net), .I1(n2827), 
            .I2(VCC_net), .I3(n49992), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_8 (.CI(n49640), .I0(n1628), 
            .I1(VCC_net), .CO(n49641));
    SB_CARRY encoder0_position_30__I_0_add_1905_9 (.CI(n49992), .I0(n2827), 
            .I1(VCC_net), .CO(n49993));
    SB_LUT4 encoder0_position_30__I_0_add_1101_7_lut (.I0(GND_net), .I1(n1629), 
            .I2(GND_net), .I3(n49639), .O(n1696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_8_lut (.I0(GND_net), .I1(n2828), 
            .I2(VCC_net), .I3(n49991), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_8 (.CI(n49991), .I0(n2828), 
            .I1(VCC_net), .CO(n49992));
    SB_CARRY add_151_20 (.CI(n49164), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n49165));
    SB_LUT4 encoder0_position_30__I_0_add_1905_7_lut (.I0(GND_net), .I1(n2829), 
            .I2(GND_net), .I3(n49990), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_7 (.CI(n49639), .I0(n1629), 
            .I1(GND_net), .CO(n49640));
    SB_CARRY encoder0_position_30__I_0_add_565_2 (.CI(VCC_net), .I0(n519), 
            .I1(GND_net), .CO(n49454));
    SB_LUT4 i23860_3_lut_4_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30350));
    defparam i23860_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY encoder0_position_30__I_0_add_1905_7 (.CI(n49990), .I0(n2829), 
            .I1(GND_net), .CO(n49991));
    SB_LUT4 encoder0_position_30__I_0_add_1101_6_lut (.I0(GND_net), .I1(n1630), 
            .I2(GND_net), .I3(n49638), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_6_lut (.I0(GND_net), .I1(n2830), 
            .I2(GND_net), .I3(n49989), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_6 (.CI(n49989), .I0(n2830), 
            .I1(GND_net), .CO(n49990));
    SB_LUT4 add_2460_7_lut (.I0(GND_net), .I1(n621), .I2(GND_net), .I3(n49453), 
            .O(n7450)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2460_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1905_5_lut (.I0(GND_net), .I1(n2831), 
            .I2(VCC_net), .I3(n49988), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_6 (.CI(n49638), .I0(n1630), 
            .I1(GND_net), .CO(n49639));
    SB_CARRY encoder0_position_30__I_0_add_1905_5 (.CI(n49988), .I0(n2831), 
            .I1(VCC_net), .CO(n49989));
    SB_LUT4 encoder0_position_30__I_0_add_1905_4_lut (.I0(GND_net), .I1(n2832), 
            .I2(GND_net), .I3(n49987), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2460_6_lut (.I0(GND_net), .I1(n622), .I2(GND_net), .I3(n49452), 
            .O(n7451)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2460_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_4 (.CI(n49987), .I0(n2832), 
            .I1(GND_net), .CO(n49988));
    SB_LUT4 encoder0_position_30__I_0_add_1101_5_lut (.I0(GND_net), .I1(n1631), 
            .I2(VCC_net), .I3(n49637), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_5 (.CI(n49637), .I0(n1631), 
            .I1(VCC_net), .CO(n49638));
    SB_LUT4 encoder0_position_30__I_0_add_1905_3_lut (.I0(GND_net), .I1(n2833), 
            .I2(VCC_net), .I3(n49986), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_3 (.CI(n49986), .I0(n2833), 
            .I1(VCC_net), .CO(n49987));
    SB_CARRY add_2460_6 (.CI(n49452), .I0(n622), .I1(GND_net), .CO(n49453));
    SB_LUT4 encoder0_position_30__I_0_add_1905_2_lut (.I0(GND_net), .I1(n953), 
            .I2(GND_net), .I3(VCC_net), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1905_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1905_2 (.CI(VCC_net), .I0(n953), 
            .I1(GND_net), .CO(n49986));
    SB_LUT4 encoder0_position_30__I_0_add_1838_27_lut (.I0(n68676), .I1(n2709), 
            .I2(VCC_net), .I3(n49985), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1838_26_lut (.I0(GND_net), .I1(n2710), 
            .I2(VCC_net), .I3(n49984), .O(n2777)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1101_4_lut (.I0(GND_net), .I1(n1632), 
            .I2(GND_net), .I3(n49636), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_26 (.CI(n49984), .I0(n2710), 
            .I1(VCC_net), .CO(n49985));
    SB_CARRY encoder0_position_30__I_0_add_1101_4 (.CI(n49636), .I0(n1632), 
            .I1(GND_net), .CO(n49637));
    SB_LUT4 encoder0_position_30__I_0_add_1838_25_lut (.I0(GND_net), .I1(n2711), 
            .I2(VCC_net), .I3(n49983), .O(n2778)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_25 (.CI(n49983), .I0(n2711), 
            .I1(VCC_net), .CO(n49984));
    SB_LUT4 encoder0_position_30__I_0_add_1101_3_lut (.I0(GND_net), .I1(n1633), 
            .I2(VCC_net), .I3(n49635), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_24_lut (.I0(GND_net), .I1(n2712), 
            .I2(VCC_net), .I3(n49982), .O(n2779)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1101_3 (.CI(n49635), .I0(n1633), 
            .I1(VCC_net), .CO(n49636));
    SB_LUT4 encoder0_position_30__I_0_add_1101_2_lut (.I0(GND_net), .I1(n941), 
            .I2(GND_net), .I3(VCC_net), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1101_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_24 (.CI(n49982), .I0(n2712), 
            .I1(VCC_net), .CO(n49983));
    SB_CARRY encoder0_position_30__I_0_add_1101_2 (.CI(VCC_net), .I0(n941), 
            .I1(GND_net), .CO(n49635));
    SB_LUT4 encoder0_position_30__I_0_add_1838_23_lut (.I0(GND_net), .I1(n2713), 
            .I2(VCC_net), .I3(n49981), .O(n2780)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_23 (.CI(n49981), .I0(n2713), 
            .I1(VCC_net), .CO(n49982));
    SB_LUT4 add_2460_5_lut (.I0(GND_net), .I1(n623), .I2(VCC_net), .I3(n49451), 
            .O(n7452)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2460_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_22_lut (.I0(GND_net), .I1(n2714), 
            .I2(VCC_net), .I3(n49980), .O(n2781)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_22 (.CI(n49980), .I0(n2714), 
            .I1(VCC_net), .CO(n49981));
    SB_LUT4 encoder0_position_30__I_0_add_1838_21_lut (.I0(GND_net), .I1(n2715), 
            .I2(VCC_net), .I3(n49979), .O(n2782)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2460_5 (.CI(n49451), .I0(n623), .I1(VCC_net), .CO(n49452));
    SB_CARRY encoder0_position_30__I_0_add_1838_21 (.CI(n49979), .I0(n2715), 
            .I1(VCC_net), .CO(n49980));
    SB_LUT4 add_2460_4_lut (.I0(GND_net), .I1(n516), .I2(GND_net), .I3(n49450), 
            .O(n7453)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2460_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1838_20_lut (.I0(GND_net), .I1(n2716), 
            .I2(VCC_net), .I3(n49978), .O(n2783)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2460_4 (.CI(n49450), .I0(n516), .I1(GND_net), .CO(n49451));
    SB_LUT4 add_2460_3_lut (.I0(GND_net), .I1(n625), .I2(VCC_net), .I3(n49449), 
            .O(n7454)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2460_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16341_3_lut_4_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30349));   // verilog/coms.v(130[12] 305[6])
    defparam i16341_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_CARRY add_2460_3 (.CI(n49449), .I0(n625), .I1(VCC_net), .CO(n49450));
    SB_CARRY encoder0_position_30__I_0_add_1838_20 (.CI(n49978), .I0(n2716), 
            .I1(VCC_net), .CO(n49979));
    SB_LUT4 encoder0_position_30__I_0_add_1838_19_lut (.I0(GND_net), .I1(n2717), 
            .I2(VCC_net), .I3(n49977), .O(n2784)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_19 (.CI(n49977), .I0(n2717), 
            .I1(VCC_net), .CO(n49978));
    SB_LUT4 encoder0_position_30__I_0_add_1838_18_lut (.I0(GND_net), .I1(n2718), 
            .I2(VCC_net), .I3(n49976), .O(n2785)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_18 (.CI(n49976), .I0(n2718), 
            .I1(VCC_net), .CO(n49977));
    SB_LUT4 encoder0_position_30__I_0_add_1838_17_lut (.I0(GND_net), .I1(n2719), 
            .I2(VCC_net), .I3(n49975), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2460_2_lut (.I0(GND_net), .I1(n518), .I2(GND_net), .I3(VCC_net), 
            .O(n7455)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2460_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_17 (.CI(n49975), .I0(n2719), 
            .I1(VCC_net), .CO(n49976));
    SB_LUT4 encoder0_position_30__I_0_add_1838_16_lut (.I0(GND_net), .I1(n2720), 
            .I2(VCC_net), .I3(n49974), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_16 (.CI(n49974), .I0(n2720), 
            .I1(VCC_net), .CO(n49975));
    SB_LUT4 encoder0_position_30__I_0_add_1838_15_lut (.I0(GND_net), .I1(n2721), 
            .I2(VCC_net), .I3(n49973), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2460_2 (.CI(VCC_net), .I0(n518), .I1(GND_net), .CO(n49449));
    SB_CARRY encoder0_position_30__I_0_add_1838_15 (.CI(n49973), .I0(n2721), 
            .I1(VCC_net), .CO(n49974));
    SB_LUT4 encoder0_position_30__I_0_add_1838_14_lut (.I0(GND_net), .I1(n2722), 
            .I2(VCC_net), .I3(n49972), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_14 (.CI(n49972), .I0(n2722), 
            .I1(VCC_net), .CO(n49973));
    SB_LUT4 i16339_3_lut_4_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30347));   // verilog/coms.v(130[12] 305[6])
    defparam i16339_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_add_1838_13_lut (.I0(GND_net), .I1(n2723), 
            .I2(VCC_net), .I3(n49971), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_13 (.CI(n49971), .I0(n2723), 
            .I1(VCC_net), .CO(n49972));
    SB_LUT4 encoder0_position_30__I_0_add_1838_12_lut (.I0(GND_net), .I1(n2724), 
            .I2(VCC_net), .I3(n49970), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_12 (.CI(n49970), .I0(n2724), 
            .I1(VCC_net), .CO(n49971));
    SB_LUT4 encoder0_position_30__I_0_add_1838_11_lut (.I0(GND_net), .I1(n2725), 
            .I2(VCC_net), .I3(n49969), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2078 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [1]), 
            .O(n56820));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2078.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1838_11 (.CI(n49969), .I0(n2725), 
            .I1(VCC_net), .CO(n49970));
    SB_LUT4 encoder0_position_30__I_0_add_1838_10_lut (.I0(GND_net), .I1(n2726), 
            .I2(VCC_net), .I3(n49968), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_10 (.CI(n49968), .I0(n2726), 
            .I1(VCC_net), .CO(n49969));
    SB_LUT4 encoder0_position_30__I_0_add_1838_9_lut (.I0(GND_net), .I1(n2727), 
            .I2(VCC_net), .I3(n49967), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_9 (.CI(n49967), .I0(n2727), 
            .I1(VCC_net), .CO(n49968));
    SB_LUT4 encoder0_position_30__I_0_add_1838_8_lut (.I0(GND_net), .I1(n2728), 
            .I2(VCC_net), .I3(n49966), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_8 (.CI(n49966), .I0(n2728), 
            .I1(VCC_net), .CO(n49967));
    SB_LUT4 encoder0_position_30__I_0_add_1838_7_lut (.I0(GND_net), .I1(n2729), 
            .I2(GND_net), .I3(n49965), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_7 (.CI(n49965), .I0(n2729), 
            .I1(GND_net), .CO(n49966));
    SB_LUT4 encoder0_position_30__I_0_add_1838_6_lut (.I0(GND_net), .I1(n2730), 
            .I2(GND_net), .I3(n49964), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_6 (.CI(n49964), .I0(n2730), 
            .I1(GND_net), .CO(n49965));
    SB_LUT4 encoder0_position_30__I_0_add_1838_5_lut (.I0(GND_net), .I1(n2731), 
            .I2(VCC_net), .I3(n49963), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_5 (.CI(n49963), .I0(n2731), 
            .I1(VCC_net), .CO(n49964));
    SB_LUT4 encoder0_position_30__I_0_add_1838_4_lut (.I0(GND_net), .I1(n2732), 
            .I2(GND_net), .I3(n49962), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_4 (.CI(n49962), .I0(n2732), 
            .I1(GND_net), .CO(n49963));
    SB_LUT4 encoder0_position_30__I_0_add_1838_3_lut (.I0(GND_net), .I1(n2733), 
            .I2(VCC_net), .I3(n49961), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_3 (.CI(n49961), .I0(n2733), 
            .I1(VCC_net), .CO(n49962));
    SB_LUT4 encoder0_position_30__I_0_add_1838_2_lut (.I0(GND_net), .I1(n952), 
            .I2(GND_net), .I3(VCC_net), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1838_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1838_2 (.CI(VCC_net), .I0(n952), 
            .I1(GND_net), .CO(n49961));
    SB_LUT4 encoder0_position_30__I_0_add_1771_26_lut (.I0(GND_net), .I1(n2610), 
            .I2(VCC_net), .I3(n49960), .O(n2677)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1771_25_lut (.I0(GND_net), .I1(n2611), 
            .I2(VCC_net), .I3(n49959), .O(n2678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n49163), .O(n1222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_25 (.CI(n49959), .I0(n2611), 
            .I1(VCC_net), .CO(n49960));
    SB_LUT4 encoder0_position_30__I_0_add_1771_24_lut (.I0(GND_net), .I1(n2612), 
            .I2(VCC_net), .I3(n49958), .O(n2679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_24 (.CI(n49958), .I0(n2612), 
            .I1(VCC_net), .CO(n49959));
    SB_CARRY add_151_9 (.CI(n49153), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n49154));
    SB_LUT4 encoder0_position_30__I_0_add_1771_23_lut (.I0(GND_net), .I1(n2613), 
            .I2(VCC_net), .I3(n49957), .O(n2680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_23 (.CI(n49957), .I0(n2613), 
            .I1(VCC_net), .CO(n49958));
    SB_LUT4 encoder0_position_30__I_0_add_1771_22_lut (.I0(GND_net), .I1(n2614), 
            .I2(VCC_net), .I3(n49956), .O(n2681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_22 (.CI(n49956), .I0(n2614), 
            .I1(VCC_net), .CO(n49957));
    SB_LUT4 encoder0_position_30__I_0_add_1771_21_lut (.I0(GND_net), .I1(n2615), 
            .I2(VCC_net), .I3(n49955), .O(n2682)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_21 (.CI(n49955), .I0(n2615), 
            .I1(VCC_net), .CO(n49956));
    SB_LUT4 encoder0_position_30__I_0_add_1771_20_lut (.I0(GND_net), .I1(n2616), 
            .I2(VCC_net), .I3(n49954), .O(n2683)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_20 (.CI(n49954), .I0(n2616), 
            .I1(VCC_net), .CO(n49955));
    SB_LUT4 encoder0_position_30__I_0_add_1771_19_lut (.I0(GND_net), .I1(n2617), 
            .I2(VCC_net), .I3(n49953), .O(n2684)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_19 (.CI(n49953), .I0(n2617), 
            .I1(VCC_net), .CO(n49954));
    SB_LUT4 encoder0_position_30__I_0_add_1771_18_lut (.I0(GND_net), .I1(n2618), 
            .I2(VCC_net), .I3(n49952), .O(n2685)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_18 (.CI(n49952), .I0(n2618), 
            .I1(VCC_net), .CO(n49953));
    SB_LUT4 encoder0_position_30__I_0_add_1771_17_lut (.I0(GND_net), .I1(n2619), 
            .I2(VCC_net), .I3(n49951), .O(n2686)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_17 (.CI(n49951), .I0(n2619), 
            .I1(VCC_net), .CO(n49952));
    SB_LUT4 encoder0_position_30__I_0_add_1771_16_lut (.I0(GND_net), .I1(n2620), 
            .I2(VCC_net), .I3(n49950), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_16 (.CI(n49950), .I0(n2620), 
            .I1(VCC_net), .CO(n49951));
    SB_CARRY add_151_19 (.CI(n49163), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n49164));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2079 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [2]), 
            .O(n56821));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2079.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1771_15_lut (.I0(GND_net), .I1(n2621), 
            .I2(VCC_net), .I3(n49949), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_15 (.CI(n49949), .I0(n2621), 
            .I1(VCC_net), .CO(n49950));
    SB_LUT4 encoder0_position_30__I_0_add_1771_14_lut (.I0(GND_net), .I1(n2622), 
            .I2(VCC_net), .I3(n49948), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n49162), .O(n1223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_14 (.CI(n49948), .I0(n2622), 
            .I1(VCC_net), .CO(n49949));
    SB_LUT4 encoder0_position_30__I_0_add_1771_13_lut (.I0(GND_net), .I1(n2623), 
            .I2(VCC_net), .I3(n49947), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_13 (.CI(n49947), .I0(n2623), 
            .I1(VCC_net), .CO(n49948));
    SB_LUT4 encoder0_position_30__I_0_add_1771_12_lut (.I0(GND_net), .I1(n2624), 
            .I2(VCC_net), .I3(n49946), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_12 (.CI(n49946), .I0(n2624), 
            .I1(VCC_net), .CO(n49947));
    SB_LUT4 encoder0_position_30__I_0_add_1771_11_lut (.I0(GND_net), .I1(n2625), 
            .I2(VCC_net), .I3(n49945), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_11 (.CI(n49945), .I0(n2625), 
            .I1(VCC_net), .CO(n49946));
    SB_LUT4 encoder0_position_30__I_0_add_1771_10_lut (.I0(GND_net), .I1(n2626), 
            .I2(VCC_net), .I3(n49944), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_10 (.CI(n49944), .I0(n2626), 
            .I1(VCC_net), .CO(n49945));
    SB_LUT4 encoder0_position_30__I_0_add_1771_9_lut (.I0(GND_net), .I1(n2627), 
            .I2(VCC_net), .I3(n49943), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_9 (.CI(n49943), .I0(n2627), 
            .I1(VCC_net), .CO(n49944));
    SB_LUT4 encoder0_position_30__I_0_add_1771_8_lut (.I0(GND_net), .I1(n2628), 
            .I2(VCC_net), .I3(n49942), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_8 (.CI(n49942), .I0(n2628), 
            .I1(VCC_net), .CO(n49943));
    SB_CARRY add_151_18 (.CI(n49162), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n49163));
    SB_LUT4 encoder0_position_30__I_0_add_1771_7_lut (.I0(GND_net), .I1(n2629), 
            .I2(GND_net), .I3(n49941), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n49161), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_7 (.CI(n49941), .I0(n2629), 
            .I1(GND_net), .CO(n49942));
    SB_LUT4 encoder0_position_30__I_0_add_1771_6_lut (.I0(GND_net), .I1(n2630), 
            .I2(GND_net), .I3(n49940), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_6 (.CI(n49940), .I0(n2630), 
            .I1(GND_net), .CO(n49941));
    SB_CARRY add_151_17 (.CI(n49161), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n49162));
    SB_LUT4 encoder0_position_30__I_0_add_1771_5_lut (.I0(GND_net), .I1(n2631), 
            .I2(VCC_net), .I3(n49939), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_5 (.CI(n49939), .I0(n2631), 
            .I1(VCC_net), .CO(n49940));
    SB_LUT4 add_151_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n49152), .O(n1233)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_8 (.CI(n49152), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n49153));
    SB_LUT4 encoder0_position_30__I_0_add_1771_4_lut (.I0(GND_net), .I1(n2632), 
            .I2(GND_net), .I3(n49938), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_4 (.CI(n49938), .I0(n2632), 
            .I1(GND_net), .CO(n49939));
    SB_LUT4 encoder0_position_30__I_0_add_1771_3_lut (.I0(GND_net), .I1(n2633), 
            .I2(VCC_net), .I3(n49937), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_3 (.CI(n49937), .I0(n2633), 
            .I1(VCC_net), .CO(n49938));
    SB_LUT4 encoder0_position_30__I_0_add_1771_2_lut (.I0(GND_net), .I1(n951), 
            .I2(GND_net), .I3(VCC_net), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1771_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1771_2 (.CI(VCC_net), .I0(n951), 
            .I1(GND_net), .CO(n49937));
    SB_LUT4 encoder0_position_30__I_0_add_1704_25_lut (.I0(n68734), .I1(n2511), 
            .I2(VCC_net), .I3(n49936), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_151_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n49160), .O(n1225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1704_24_lut (.I0(GND_net), .I1(n2512), 
            .I2(VCC_net), .I3(n49935), .O(n2579)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_24 (.CI(n49935), .I0(n2512), 
            .I1(VCC_net), .CO(n49936));
    SB_LUT4 encoder0_position_30__I_0_add_1704_23_lut (.I0(GND_net), .I1(n2513), 
            .I2(VCC_net), .I3(n49934), .O(n2580)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_23 (.CI(n49934), .I0(n2513), 
            .I1(VCC_net), .CO(n49935));
    SB_LUT4 encoder0_position_30__I_0_add_1704_22_lut (.I0(GND_net), .I1(n2514), 
            .I2(VCC_net), .I3(n49933), .O(n2581)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_22 (.CI(n49933), .I0(n2514), 
            .I1(VCC_net), .CO(n49934));
    SB_CARRY add_151_16 (.CI(n49160), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n49161));
    SB_LUT4 encoder0_position_30__I_0_add_1704_21_lut (.I0(GND_net), .I1(n2515), 
            .I2(VCC_net), .I3(n49932), .O(n2582)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_21 (.CI(n49932), .I0(n2515), 
            .I1(VCC_net), .CO(n49933));
    SB_LUT4 encoder0_position_30__I_0_add_1704_20_lut (.I0(GND_net), .I1(n2516), 
            .I2(VCC_net), .I3(n49931), .O(n2583)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_20 (.CI(n49931), .I0(n2516), 
            .I1(VCC_net), .CO(n49932));
    SB_LUT4 encoder0_position_30__I_0_add_1704_19_lut (.I0(GND_net), .I1(n2517), 
            .I2(VCC_net), .I3(n49930), .O(n2584)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_19 (.CI(n49930), .I0(n2517), 
            .I1(VCC_net), .CO(n49931));
    SB_LUT4 encoder0_position_30__I_0_add_1704_18_lut (.I0(GND_net), .I1(n2518), 
            .I2(VCC_net), .I3(n49929), .O(n2585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_3 (.CI(n49147), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n49148));
    SB_CARRY encoder0_position_30__I_0_add_1704_18 (.CI(n49929), .I0(n2518), 
            .I1(VCC_net), .CO(n49930));
    SB_LUT4 encoder0_position_30__I_0_add_1704_17_lut (.I0(GND_net), .I1(n2519), 
            .I2(VCC_net), .I3(n49928), .O(n2586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_17 (.CI(n49928), .I0(n2519), 
            .I1(VCC_net), .CO(n49929));
    SB_LUT4 encoder0_position_30__I_0_add_1704_16_lut (.I0(GND_net), .I1(n2520), 
            .I2(VCC_net), .I3(n49927), .O(n2587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_16 (.CI(n49927), .I0(n2520), 
            .I1(VCC_net), .CO(n49928));
    SB_LUT4 encoder0_position_30__I_0_add_1704_15_lut (.I0(GND_net), .I1(n2521), 
            .I2(VCC_net), .I3(n49926), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_15 (.CI(n49926), .I0(n2521), 
            .I1(VCC_net), .CO(n49927));
    SB_LUT4 encoder0_position_30__I_0_add_1704_14_lut (.I0(GND_net), .I1(n2522), 
            .I2(VCC_net), .I3(n49925), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_14 (.CI(n49925), .I0(n2522), 
            .I1(VCC_net), .CO(n49926));
    SB_LUT4 encoder0_position_30__I_0_add_1704_13_lut (.I0(GND_net), .I1(n2523), 
            .I2(VCC_net), .I3(n49924), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_13 (.CI(n49924), .I0(n2523), 
            .I1(VCC_net), .CO(n49925));
    SB_LUT4 encoder0_position_30__I_0_add_1704_12_lut (.I0(GND_net), .I1(n2524), 
            .I2(VCC_net), .I3(n49923), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_12 (.CI(n49923), .I0(n2524), 
            .I1(VCC_net), .CO(n49924));
    SB_LUT4 encoder0_position_30__I_0_add_1704_11_lut (.I0(GND_net), .I1(n2525), 
            .I2(VCC_net), .I3(n49922), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_11 (.CI(n49922), .I0(n2525), 
            .I1(VCC_net), .CO(n49923));
    SB_LUT4 encoder0_position_30__I_0_add_1704_10_lut (.I0(GND_net), .I1(n2526), 
            .I2(VCC_net), .I3(n49921), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_10 (.CI(n49921), .I0(n2526), 
            .I1(VCC_net), .CO(n49922));
    SB_LUT4 encoder0_position_30__I_0_add_1704_9_lut (.I0(GND_net), .I1(n2527), 
            .I2(VCC_net), .I3(n49920), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_9 (.CI(n49920), .I0(n2527), 
            .I1(VCC_net), .CO(n49921));
    SB_LUT4 encoder0_position_30__I_0_add_1704_8_lut (.I0(GND_net), .I1(n2528), 
            .I2(VCC_net), .I3(n49919), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n49159), .O(n1226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_8 (.CI(n49919), .I0(n2528), 
            .I1(VCC_net), .CO(n49920));
    SB_LUT4 encoder0_position_30__I_0_add_1704_7_lut (.I0(GND_net), .I1(n2529), 
            .I2(GND_net), .I3(n49918), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_7 (.CI(n49918), .I0(n2529), 
            .I1(GND_net), .CO(n49919));
    SB_LUT4 encoder0_position_30__I_0_add_1704_6_lut (.I0(GND_net), .I1(n2530), 
            .I2(GND_net), .I3(n49917), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_6 (.CI(n49917), .I0(n2530), 
            .I1(GND_net), .CO(n49918));
    SB_LUT4 encoder0_position_30__I_0_add_1704_5_lut (.I0(GND_net), .I1(n2531), 
            .I2(VCC_net), .I3(n49916), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_5 (.CI(n49916), .I0(n2531), 
            .I1(VCC_net), .CO(n49917));
    SB_LUT4 encoder0_position_30__I_0_add_1704_4_lut (.I0(GND_net), .I1(n2532), 
            .I2(GND_net), .I3(n49915), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_4 (.CI(n49915), .I0(n2532), 
            .I1(GND_net), .CO(n49916));
    SB_LUT4 encoder0_position_30__I_0_add_1704_3_lut (.I0(GND_net), .I1(n2533), 
            .I2(VCC_net), .I3(n49914), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_3 (.CI(n49914), .I0(n2533), 
            .I1(VCC_net), .CO(n49915));
    SB_LUT4 encoder0_position_30__I_0_add_1704_2_lut (.I0(GND_net), .I1(n950), 
            .I2(GND_net), .I3(VCC_net), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1704_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1704_2 (.CI(VCC_net), .I0(n950), 
            .I1(GND_net), .CO(n49914));
    SB_LUT4 encoder0_position_30__I_0_add_1637_24_lut (.I0(n68703), .I1(n2412), 
            .I2(VCC_net), .I3(n49913), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_30__I_0_add_1637_23_lut (.I0(GND_net), .I1(n2413), 
            .I2(VCC_net), .I3(n49912), .O(n2480)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_23 (.CI(n49912), .I0(n2413), 
            .I1(VCC_net), .CO(n49913));
    SB_LUT4 add_151_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n49151), .O(n1234)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_22_lut (.I0(GND_net), .I1(n2414), 
            .I2(VCC_net), .I3(n49911), .O(n2481)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_22 (.CI(n49911), .I0(n2414), 
            .I1(VCC_net), .CO(n49912));
    SB_LUT4 encoder0_position_30__I_0_add_1637_21_lut (.I0(GND_net), .I1(n2415), 
            .I2(VCC_net), .I3(n49910), .O(n2482)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_21 (.CI(n49910), .I0(n2415), 
            .I1(VCC_net), .CO(n49911));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2080 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [3]), 
            .O(n56822));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2080.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2081 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [4]), 
            .O(n56823));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2081.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1637_20_lut (.I0(GND_net), .I1(n2416), 
            .I2(VCC_net), .I3(n49909), .O(n2483)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_20 (.CI(n49909), .I0(n2416), 
            .I1(VCC_net), .CO(n49910));
    SB_LUT4 encoder0_position_30__I_0_add_1637_19_lut (.I0(GND_net), .I1(n2417), 
            .I2(VCC_net), .I3(n49908), .O(n2484)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_19 (.CI(n49908), .I0(n2417), 
            .I1(VCC_net), .CO(n49909));
    SB_LUT4 encoder0_position_30__I_0_add_1637_18_lut (.I0(GND_net), .I1(n2418), 
            .I2(VCC_net), .I3(n49907), .O(n2485)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_18 (.CI(n49907), .I0(n2418), 
            .I1(VCC_net), .CO(n49908));
    SB_LUT4 encoder0_position_30__I_0_add_1637_17_lut (.I0(GND_net), .I1(n2419), 
            .I2(VCC_net), .I3(n49906), .O(n2486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_17 (.CI(n49906), .I0(n2419), 
            .I1(VCC_net), .CO(n49907));
    SB_LUT4 encoder0_position_30__I_0_add_1637_16_lut (.I0(GND_net), .I1(n2420), 
            .I2(VCC_net), .I3(n49905), .O(n2487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_16 (.CI(n49905), .I0(n2420), 
            .I1(VCC_net), .CO(n49906));
    SB_LUT4 encoder0_position_30__I_0_add_1637_15_lut (.I0(GND_net), .I1(n2421), 
            .I2(VCC_net), .I3(n49904), .O(n2488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_15 (.CI(n49904), .I0(n2421), 
            .I1(VCC_net), .CO(n49905));
    SB_LUT4 encoder0_position_30__I_0_add_1637_14_lut (.I0(GND_net), .I1(n2422), 
            .I2(VCC_net), .I3(n49903), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2082 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [5]), 
            .O(n56824));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2082.LUT_INIT = 16'h2300;
    SB_LUT4 add_151_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1239)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_14 (.CI(n49903), .I0(n2422), 
            .I1(VCC_net), .CO(n49904));
    SB_LUT4 encoder0_position_30__I_0_add_1637_13_lut (.I0(GND_net), .I1(n2423), 
            .I2(VCC_net), .I3(n49902), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_13 (.CI(n49902), .I0(n2423), 
            .I1(VCC_net), .CO(n49903));
    SB_LUT4 encoder0_position_30__I_0_add_1637_12_lut (.I0(GND_net), .I1(n2424), 
            .I2(VCC_net), .I3(n49901), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_12 (.CI(n49901), .I0(n2424), 
            .I1(VCC_net), .CO(n49902));
    SB_LUT4 encoder0_position_30__I_0_add_1637_11_lut (.I0(GND_net), .I1(n2425), 
            .I2(VCC_net), .I3(n49900), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_11 (.CI(n49900), .I0(n2425), 
            .I1(VCC_net), .CO(n49901));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2083 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [6]), 
            .O(n56825));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2083.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1637_10_lut (.I0(GND_net), .I1(n2426), 
            .I2(VCC_net), .I3(n49899), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29492_3_lut (.I0(n944), .I1(n1932), .I2(n1933), .I3(GND_net), 
            .O(n43398));
    defparam i29492_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY encoder0_position_30__I_0_add_1637_10 (.CI(n49899), .I0(n2426), 
            .I1(VCC_net), .CO(n49900));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2084 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [7]), 
            .O(n56826));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2084.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1637_9_lut (.I0(GND_net), .I1(n2427), 
            .I2(VCC_net), .I3(n49898), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2085 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [0]), 
            .O(n56827));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2085.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16335_3_lut_4_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30343));   // verilog/coms.v(130[12] 305[6])
    defparam i16335_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2086 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [1]), 
            .O(n56828));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2086.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2087 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [2]), 
            .O(n56829));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2087.LUT_INIT = 16'h2300;
    SB_CARRY encoder0_position_30__I_0_add_1637_9 (.CI(n49898), .I0(n2427), 
            .I1(VCC_net), .CO(n49899));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2088 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [3]), 
            .O(n56830));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2088.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1637_8_lut (.I0(GND_net), .I1(n2428), 
            .I2(VCC_net), .I3(n49897), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15723_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[1] [1]), 
            .I3(control_mode[1]), .O(n29731));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15723_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15708_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[20] [1]), 
            .I3(current_limit[9]), .O(n29716));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15708_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY encoder0_position_30__I_0_add_1637_8 (.CI(n49897), .I0(n2428), 
            .I1(VCC_net), .CO(n49898));
    SB_LUT4 i15704_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[20] [2]), 
            .I3(current_limit[10]), .O(n29712));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15704_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15700_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[20] [3]), 
            .I3(current_limit[11]), .O(n29708));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15700_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 encoder0_position_30__I_0_add_1637_7_lut (.I0(GND_net), .I1(n2429), 
            .I2(GND_net), .I3(n49896), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_7 (.CI(n49896), .I0(n2429), 
            .I1(GND_net), .CO(n49897));
    SB_LUT4 encoder0_position_30__I_0_add_1637_6_lut (.I0(GND_net), .I1(n2430), 
            .I2(GND_net), .I3(n49895), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21765_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[20] [5]), 
            .I3(current_limit[13]), .O(n29706));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i21765_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16273_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[21] [4]), 
            .I3(current_limit[4]), .O(n30281));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i16273_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16242_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[21] [5]), 
            .I3(current_limit[5]), .O(n30250));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i16242_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15482_3_lut_4_lut (.I0(\data_in_frame[16] [3]), .I1(rx_data[3]), 
            .I2(reset), .I3(n92), .O(n29490));   // verilog/coms.v(130[12] 305[6])
    defparam i15482_3_lut_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY encoder0_position_30__I_0_add_1637_6 (.CI(n49895), .I0(n2430), 
            .I1(GND_net), .CO(n49896));
    SB_LUT4 encoder0_position_30__I_0_add_1637_5_lut (.I0(GND_net), .I1(n2431), 
            .I2(VCC_net), .I3(n49894), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21764_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[20] [7]), 
            .I3(current_limit[15]), .O(n29662));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i21764_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16224_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[21] [6]), 
            .I3(current_limit[6]), .O(n30232));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i16224_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY add_151_7 (.CI(n49151), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n49152));
    SB_CARRY add_151_15 (.CI(n49159), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n49160));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2089 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [4]), 
            .O(n56831));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2089.LUT_INIT = 16'h2300;
    SB_LUT4 add_151_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n49150), .O(n1235)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_5 (.CI(n49894), .I0(n2431), 
            .I1(VCC_net), .CO(n49895));
    SB_LUT4 i15699_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[20] [4]), 
            .I3(current_limit[12]), .O(n29707));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15699_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 encoder0_position_30__I_0_add_1637_4_lut (.I0(GND_net), .I1(n2432), 
            .I2(GND_net), .I3(n49893), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_4 (.CI(n49893), .I0(n2432), 
            .I1(GND_net), .CO(n49894));
    SB_LUT4 encoder0_position_30__I_0_add_1637_3_lut (.I0(GND_net), .I1(n2433), 
            .I2(VCC_net), .I3(n49892), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2090 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [2]), 
            .O(n56951));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2090.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1034_15_lut (.I0(n68902), .I1(n1521), 
            .I2(VCC_net), .I3(n49610), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15485_3_lut_4_lut (.I0(\data_in_frame[16] [4]), .I1(rx_data[4]), 
            .I2(reset), .I3(n92), .O(n29493));   // verilog/coms.v(130[12] 305[6])
    defparam i15485_3_lut_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i15488_3_lut_4_lut (.I0(\data_in_frame[16] [5]), .I1(rx_data[5]), 
            .I2(reset), .I3(n92), .O(n29496));   // verilog/coms.v(130[12] 305[6])
    defparam i15488_3_lut_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 encoder0_position_30__I_0_add_1034_14_lut (.I0(GND_net), .I1(n1522), 
            .I2(VCC_net), .I3(n49609), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_14 (.CI(n49609), .I0(n1522), 
            .I1(VCC_net), .CO(n49610));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5752));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_30__I_0_add_1637_3 (.CI(n49892), .I0(n2433), 
            .I1(VCC_net), .CO(n49893));
    SB_LUT4 add_151_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n49158), .O(n1227)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1637_2_lut (.I0(GND_net), .I1(n949), 
            .I2(GND_net), .I3(VCC_net), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1637_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n49147));
    SB_LUT4 encoder0_position_30__I_0_add_1034_13_lut (.I0(GND_net), .I1(n1523), 
            .I2(VCC_net), .I3(n49608), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1637_2 (.CI(VCC_net), .I0(n949), 
            .I1(GND_net), .CO(n49892));
    SB_LUT4 i16274_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[21] [3]), 
            .I3(current_limit[3]), .O(n30282));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i16274_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 encoder0_position_30__I_0_add_1570_23_lut (.I0(n68609), .I1(n2313), 
            .I2(VCC_net), .I3(n49891), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i16291_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[21] [2]), 
            .I3(current_limit[2]), .O(n30299));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i16291_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15726_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[1] [4]), 
            .I3(control_mode[4]), .O(n29734));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15726_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 encoder0_position_30__I_0_add_1570_22_lut (.I0(GND_net), .I1(n2314), 
            .I2(VCC_net), .I3(n49890), .O(n2381)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_22 (.CI(n49890), .I0(n2314), 
            .I1(VCC_net), .CO(n49891));
    SB_CARRY encoder0_position_30__I_0_add_1034_13 (.CI(n49608), .I0(n1523), 
            .I1(VCC_net), .CO(n49609));
    SB_LUT4 encoder0_position_30__I_0_add_1570_21_lut (.I0(GND_net), .I1(n2315), 
            .I2(VCC_net), .I3(n49889), .O(n2382)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_21 (.CI(n49889), .I0(n2315), 
            .I1(VCC_net), .CO(n49890));
    SB_LUT4 encoder0_position_30__I_0_add_1570_20_lut (.I0(GND_net), .I1(n2316), 
            .I2(VCC_net), .I3(n49888), .O(n2383)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15491_3_lut_4_lut (.I0(\data_in_frame[16] [6]), .I1(rx_data[6]), 
            .I2(reset), .I3(n92), .O(n29499));   // verilog/coms.v(130[12] 305[6])
    defparam i15491_3_lut_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY encoder0_position_30__I_0_add_1570_20 (.CI(n49888), .I0(n2316), 
            .I1(VCC_net), .CO(n49889));
    SB_LUT4 encoder0_position_30__I_0_add_1570_19_lut (.I0(GND_net), .I1(n2317), 
            .I2(VCC_net), .I3(n49887), .O(n2384)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_19 (.CI(n49887), .I0(n2317), 
            .I1(VCC_net), .CO(n49888));
    SB_LUT4 encoder0_position_30__I_0_add_1570_18_lut (.I0(GND_net), .I1(n2318), 
            .I2(VCC_net), .I3(n49886), .O(n2385)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_18 (.CI(n49886), .I0(n2318), 
            .I1(VCC_net), .CO(n49887));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2091 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [3]), 
            .O(n56950));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2091.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1570_17_lut (.I0(GND_net), .I1(n2319), 
            .I2(VCC_net), .I3(n49885), .O(n2386)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_17 (.CI(n49885), .I0(n2319), 
            .I1(VCC_net), .CO(n49886));
    SB_LUT4 encoder0_position_30__I_0_add_1570_16_lut (.I0(GND_net), .I1(n2320), 
            .I2(VCC_net), .I3(n49884), .O(n2387)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_12_lut (.I0(GND_net), .I1(n1524), 
            .I2(VCC_net), .I3(n49607), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_16 (.CI(n49884), .I0(n2320), 
            .I1(VCC_net), .CO(n49885));
    SB_LUT4 encoder0_position_30__I_0_add_1570_15_lut (.I0(GND_net), .I1(n2321), 
            .I2(VCC_net), .I3(n49883), .O(n2388)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_15 (.CI(n49883), .I0(n2321), 
            .I1(VCC_net), .CO(n49884));
    SB_CARRY encoder0_position_30__I_0_add_1034_12 (.CI(n49607), .I0(n1524), 
            .I1(VCC_net), .CO(n49608));
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2092 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [4]), 
            .O(n56949));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2092.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1034_11_lut (.I0(GND_net), .I1(n1525), 
            .I2(VCC_net), .I3(n49606), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_11 (.CI(n49606), .I0(n1525), 
            .I1(VCC_net), .CO(n49607));
    SB_LUT4 encoder0_position_30__I_0_add_1570_14_lut (.I0(GND_net), .I1(n2322), 
            .I2(VCC_net), .I3(n49882), .O(n2389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_10_lut (.I0(GND_net), .I1(n1526), 
            .I2(VCC_net), .I3(n49605), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_14 (.CI(n49882), .I0(n2322), 
            .I1(VCC_net), .CO(n49883));
    SB_CARRY encoder0_position_30__I_0_add_1034_10 (.CI(n49605), .I0(n1526), 
            .I1(VCC_net), .CO(n49606));
    SB_LUT4 encoder0_position_30__I_0_add_1570_13_lut (.I0(GND_net), .I1(n2323), 
            .I2(VCC_net), .I3(n49881), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_13 (.CI(n49881), .I0(n2323), 
            .I1(VCC_net), .CO(n49882));
    SB_LUT4 encoder0_position_30__I_0_add_1034_9_lut (.I0(GND_net), .I1(n1527), 
            .I2(VCC_net), .I3(n49604), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1570_12_lut (.I0(GND_net), .I1(n2324), 
            .I2(VCC_net), .I3(n49880), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_i1445_3_lut (.I0(n2122), .I1(n2189), 
            .I2(n2148), .I3(GND_net), .O(n2221));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1445_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_30__I_0_add_1034_9 (.CI(n49604), .I0(n1527), 
            .I1(VCC_net), .CO(n49605));
    SB_CARRY encoder0_position_30__I_0_add_1570_12 (.CI(n49880), .I0(n2324), 
            .I1(VCC_net), .CO(n49881));
    SB_LUT4 encoder0_position_30__I_0_add_1570_11_lut (.I0(GND_net), .I1(n2325), 
            .I2(VCC_net), .I3(n49879), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_11 (.CI(n49879), .I0(n2325), 
            .I1(VCC_net), .CO(n49880));
    SB_LUT4 encoder0_position_30__I_0_add_1034_8_lut (.I0(GND_net), .I1(n1528), 
            .I2(VCC_net), .I3(n49603), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_8 (.CI(n49603), .I0(n1528), 
            .I1(VCC_net), .CO(n49604));
    SB_LUT4 encoder0_position_30__I_0_add_1570_10_lut (.I0(GND_net), .I1(n2326), 
            .I2(VCC_net), .I3(n49878), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_10 (.CI(n49878), .I0(n2326), 
            .I1(VCC_net), .CO(n49879));
    SB_LUT4 encoder0_position_30__I_0_add_1570_9_lut (.I0(GND_net), .I1(n2327), 
            .I2(VCC_net), .I3(n49877), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16459_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[1] [5]), 
            .I3(control_mode[5]), .O(n30467));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i16459_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY encoder0_position_30__I_0_add_1570_9 (.CI(n49877), .I0(n2327), 
            .I1(VCC_net), .CO(n49878));
    SB_LUT4 encoder0_position_30__I_0_add_1570_8_lut (.I0(GND_net), .I1(n2328), 
            .I2(VCC_net), .I3(n49876), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_2093 (.I0(n1929), .I1(n43398), .I2(n1930), .I3(n1931), 
            .O(n58681));
    defparam i1_4_lut_adj_2093.LUT_INIT = 16'ha080;
    SB_CARRY encoder0_position_30__I_0_add_1570_8 (.CI(n49876), .I0(n2328), 
            .I1(VCC_net), .CO(n49877));
    SB_LUT4 encoder0_position_30__I_0_add_1570_7_lut (.I0(GND_net), .I1(n2329), 
            .I2(GND_net), .I3(n49875), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_7 (.CI(n49875), .I0(n2329), 
            .I1(GND_net), .CO(n49876));
    SB_LUT4 i1_4_lut_adj_2094 (.I0(n1918), .I1(n1920), .I2(n1922), .I3(n61012), 
            .O(n61018));
    defparam i1_4_lut_adj_2094.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_1570_6_lut (.I0(GND_net), .I1(n2330), 
            .I2(GND_net), .I3(n49874), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2095 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [0]), 
            .O(n56948));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2095.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_add_1034_7_lut (.I0(GND_net), .I1(n1529), 
            .I2(GND_net), .I3(n49602), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_6 (.CI(n49874), .I0(n2330), 
            .I1(GND_net), .CO(n49875));
    SB_LUT4 encoder0_position_30__I_0_add_1570_5_lut (.I0(GND_net), .I1(n2331), 
            .I2(VCC_net), .I3(n49873), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_7 (.CI(n49602), .I0(n1529), 
            .I1(GND_net), .CO(n49603));
    SB_CARRY encoder0_position_30__I_0_add_1570_5 (.CI(n49873), .I0(n2331), 
            .I1(VCC_net), .CO(n49874));
    SB_LUT4 encoder0_position_30__I_0_add_1570_4_lut (.I0(GND_net), .I1(n2332), 
            .I2(GND_net), .I3(n49872), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_30__I_0_add_1034_6_lut (.I0(GND_net), .I1(n1530), 
            .I2(GND_net), .I3(n49601), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_4 (.CI(n49872), .I0(n2332), 
            .I1(GND_net), .CO(n49873));
    SB_LUT4 encoder0_position_30__I_0_add_1570_3_lut (.I0(GND_net), .I1(n2333), 
            .I2(VCC_net), .I3(n49871), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_3 (.CI(n49871), .I0(n2333), 
            .I1(VCC_net), .CO(n49872));
    SB_CARRY encoder0_position_30__I_0_add_1034_6 (.CI(n49601), .I0(n1530), 
            .I1(GND_net), .CO(n49602));
    SB_LUT4 encoder0_position_30__I_0_add_1570_2_lut (.I0(GND_net), .I1(n948), 
            .I2(GND_net), .I3(VCC_net), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1570_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1570_2 (.CI(VCC_net), .I0(n948), 
            .I1(GND_net), .CO(n49871));
    SB_LUT4 encoder0_position_30__I_0_add_1503_22_lut (.I0(n68857), .I1(n2214), 
            .I2(VCC_net), .I3(n49870), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_151_6 (.CI(n49150), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n49151));
    SB_LUT4 encoder0_position_30__I_0_add_1034_5_lut (.I0(GND_net), .I1(n1531), 
            .I2(VCC_net), .I3(n49600), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1034_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_30__I_0_add_1034_5 (.CI(n49600), .I0(n1531), 
            .I1(VCC_net), .CO(n49601));
    SB_LUT4 i1_4_lut_adj_2096 (.I0(n58681), .I1(n1921), .I2(n1923), .I3(n1924), 
            .O(n61328));
    defparam i1_4_lut_adj_2096.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_add_1503_21_lut (.I0(GND_net), .I1(n2215), 
            .I2(VCC_net), .I3(n49869), .O(n2282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_30__I_0_add_1503_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_1086_i15_2_lut (.I0(r_Clock_Count_adj_5987[7]), .I1(o_Rx_DV_N_3488[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5838));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1086_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY encoder0_position_30__I_0_add_1503_21 (.CI(n49869), .I0(n2215), 
            .I1(VCC_net), .CO(n49870));
    SB_LUT4 LessThan_1086_i9_2_lut (.I0(r_Clock_Count_adj_5987[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5835));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1086_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1086_i13_2_lut (.I0(r_Clock_Count_adj_5987[6]), .I1(o_Rx_DV_N_3488[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5837));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1086_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2097 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [1]), 
            .O(n56947));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2097.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_1086_i11_2_lut (.I0(r_Clock_Count_adj_5987[5]), .I1(o_Rx_DV_N_3488[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5836));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1086_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2098 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [3]), 
            .O(n56946));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2098.LUT_INIT = 16'h2300;
    SB_LUT4 i47172_3_lut (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[17] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n62858));
    defparam i47172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2099 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [5]), 
            .O(n56945));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2099.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2100 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [6]), 
            .O(n56944));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2100.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2101 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [7]), 
            .O(n56943));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2101.LUT_INIT = 16'h2300;
    SB_LUT4 i47173_3_lut (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[19] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n62859));
    defparam i47173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2102 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [1]), 
            .O(n56942));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2102.LUT_INIT = 16'h2300;
    SB_LUT4 i47026_3_lut (.I0(\data_out_frame[22] [3]), .I1(\data_out_frame[23] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n62712));
    defparam i47026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5753));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2103 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [3]), 
            .O(n56941));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2103.LUT_INIT = 16'h2300;
    SB_LUT4 i47025_3_lut (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[21] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n62711));
    defparam i47025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2104 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [4]), 
            .O(n56940));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2104.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2105 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [6]), 
            .O(n56771));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2105.LUT_INIT = 16'h2300;
    SB_LUT4 i15501_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n22726), .I3(GND_net), .O(n29509));   // verilog/coms.v(130[12] 305[6])
    defparam i15501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2106 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [7]), 
            .O(n56939));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2106.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_1086_i4_4_lut (.I0(r_Clock_Count_adj_5987[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count_adj_5987[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5832));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1086_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i51952_3_lut (.I0(n4_adj_5832), .I1(o_Rx_DV_N_3488[5]), .I2(n11_adj_5836), 
            .I3(GND_net), .O(n67638));   // verilog/uart_tx.v(117[17:57])
    defparam i51952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51953_3_lut (.I0(n67638), .I1(o_Rx_DV_N_3488[6]), .I2(n13_adj_5837), 
            .I3(GND_net), .O(n67639));   // verilog/uart_tx.v(117[17:57])
    defparam i51953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2107 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [0]), 
            .O(n56938));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2107.LUT_INIT = 16'h2300;
    SB_LUT4 i21760_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[20] [6]), 
            .I3(current_limit[14]), .O(n29705));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i21760_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2108 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [1]), 
            .O(n29117));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2108.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2109 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [2]), 
            .O(n29116));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2109.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5754));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2110 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [3]), 
            .O(n29115));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2110.LUT_INIT = 16'h2300;
    SB_LUT4 i51365_4_lut (.I0(n13_adj_5837), .I1(n11_adj_5836), .I2(n9_adj_5835), 
            .I3(n66171), .O(n67051));
    defparam i51365_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2111 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [4]), 
            .O(n56937));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2111.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_1086_i8_3_lut (.I0(n6_adj_5833), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5835), .I3(GND_net), .O(n8_adj_5834));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1086_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50992_3_lut (.I0(n67639), .I1(o_Rx_DV_N_3488[7]), .I2(n15_adj_5838), 
            .I3(GND_net), .O(n66678));   // verilog/uart_tx.v(117[17:57])
    defparam i50992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15845_3_lut (.I0(\data_in_frame[1] [0]), .I1(rx_data[0]), .I2(n57044), 
            .I3(GND_net), .O(n29853));   // verilog/coms.v(130[12] 305[6])
    defparam i15845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i51956_4_lut (.I0(n66678), .I1(n8_adj_5834), .I2(n15_adj_5838), 
            .I3(n67051), .O(n67642));   // verilog/uart_tx.v(117[17:57])
    defparam i51956_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51957_3_lut (.I0(n67642), .I1(o_Rx_DV_N_3488[8]), .I2(r_Clock_Count_adj_5987[8]), 
            .I3(GND_net), .O(n4940));   // verilog/uart_tx.v(117[17:57])
    defparam i51957_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2112 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [5]), 
            .O(n56936));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2112.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2113 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [6]), 
            .O(n56935));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2113.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2114 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [7]), 
            .O(n56934));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2114.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2115 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [0]), 
            .O(n56933));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2115.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2116 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [1]), 
            .O(n56932));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2116.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5759));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_4310_i13_3_lut (.I0(encoder0_position[12]), .I1(n20_adj_5694), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n945));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2117 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [2]), 
            .O(n56931));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2117.LUT_INIT = 16'h2300;
    SB_LUT4 i27697_4_lut_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15_adj_5681), .I3(n15), .O(n41621));
    defparam i27697_4_lut_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 i15727_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[21] [7]), 
            .I3(current_limit[7]), .O(n29735));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15727_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2118 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [3]), 
            .O(n56930));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2118.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2119 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [4]), 
            .O(n56929));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2119.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2120 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [5]), 
            .O(n56928));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2120.LUT_INIT = 16'h2300;
    SB_LUT4 mux_4310_i14_3_lut (.I0(encoder0_position[13]), .I1(n19_adj_5695), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n944));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2121 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [6]), 
            .O(n56927));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2121.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_30__I_0_i1321_3_lut (.I0(n944), .I1(n2001), 
            .I2(n1950), .I3(GND_net), .O(n2033));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i15_3_lut (.I0(encoder0_position[14]), .I1(n18_adj_5696), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n943));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1253_3_lut (.I0(n943), .I1(n1901), 
            .I2(n1851), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1253_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1320_3_lut (.I0(n1933), .I1(n2000), 
            .I2(n1950), .I3(GND_net), .O(n2032));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i42298_2_lut (.I0(r_SM_Main_adj_5986[2]), .I1(r_SM_Main_adj_5986[0]), 
            .I2(GND_net), .I3(GND_net), .O(n57935));
    defparam i42298_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2122 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [7]), 
            .O(n56926));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2122.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2123 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [0]), 
            .O(n56925));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2123.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2124 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [1]), 
            .O(n56924));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2124.LUT_INIT = 16'h2300;
    SB_LUT4 i16192_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n60708), 
            .I3(n27_adj_5781), .O(n30200));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16192_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2125 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [2]), 
            .O(n56923));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2125.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2126 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [3]), 
            .O(n56922));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2126.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2127 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [4]), 
            .O(n56921));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2127.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2128 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [5]), 
            .O(n56920));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2128.LUT_INIT = 16'h2300;
    SB_LUT4 i16193_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n60692), 
            .I3(n27_adj_5781), .O(n30201));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16193_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2129 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [6]), 
            .O(n56919));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2129.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2130 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [5]), 
            .O(n56832));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2130.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2131 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [6]), 
            .O(n56833));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2131.LUT_INIT = 16'h2300;
    SB_LUT4 i12_4_lut_adj_2132 (.I0(\data_in_frame[19] [6]), .I1(n28379), 
            .I2(n28434), .I3(rx_data[6]), .O(n56037));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2132.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5761));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12_4_lut_adj_2133 (.I0(\data_in_frame[19] [5]), .I1(n28379), 
            .I2(n28434), .I3(rx_data[5]), .O(n56041));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2133.LUT_INIT = 16'h3a0a;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(current[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5711));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut_adj_2134 (.I0(\data_in_frame[19] [4]), .I1(n28379), 
            .I2(n28434), .I3(rx_data[4]), .O(n56045));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2134.LUT_INIT = 16'h3a0a;
    SB_LUT4 LessThan_11_i7_2_lut (.I0(current[3]), .I1(duty[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5724));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15709_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[20] [0]), 
            .I3(current_limit[8]), .O(n29717));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15709_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2135 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [7]), 
            .O(n56834));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2135.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2136 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [0]), 
            .O(n56835));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2136.LUT_INIT = 16'h2300;
    SB_LUT4 i53102_4_lut (.I0(n61328), .I1(n61018), .I2(n1919), .I3(n1917), 
            .O(n1950));
    defparam i53102_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(current[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5722));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i27085_4_lut (.I0(n65433), .I1(n65432), .I2(rx_data[3]), .I3(\data_in_frame[19] [3]), 
            .O(n41018));   // verilog/coms.v(94[13:20])
    defparam i27085_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i27086_3_lut (.I0(n41018), .I1(\data_in_frame[19] [3]), .I2(reset), 
            .I3(GND_net), .O(n30207));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i27086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_2137 (.I0(\data_in_frame[19] [2]), .I1(n28379), 
            .I2(n28434), .I3(rx_data[2]), .O(n56049));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2137.LUT_INIT = 16'h3a0a;
    SB_LUT4 i2_2_lut (.I0(dti_counter[1]), .I1(dti_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_5902));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i16367_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[1] [6]), 
            .I3(control_mode[6]), .O(n30375));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i16367_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(current[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5716));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15630_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[1] [0]), 
            .I3(control_mode[0]), .O(n29638));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15630_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 encoder0_position_30__I_0_i1252_3_lut (.I0(n1833), .I1(n1900), 
            .I2(n1851), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1252_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16202_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5966[1]), 
            .I2(n10_adj_5844), .I3(n25535), .O(n30210));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16202_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i6_4_lut_adj_2138 (.I0(dti_counter[7]), .I1(dti_counter[4]), 
            .I2(dti_counter[5]), .I3(dti_counter[6]), .O(n14_adj_5901));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i6_4_lut_adj_2138.LUT_INIT = 16'hfffe;
    SB_LUT4 i16203_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5966[2]), 
            .I2(n4_adj_5727), .I3(n25540), .O(n30211));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16203_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16340_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[1] [7]), 
            .I3(control_mode[7]), .O(n30348));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i16340_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16204_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5966[3]), 
            .I2(n4_adj_5727), .I3(n25535), .O(n30212));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16204_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16205_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5966[4]), 
            .I2(n4_adj_5728), .I3(n25540), .O(n30213));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16205_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(current[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5713));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16206_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5966[5]), 
            .I2(n4_adj_5728), .I3(n25535), .O(n30214));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16206_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_30__I_0_i1319_3_lut (.I0(n1932), .I1(n1999), 
            .I2(n1950), .I3(GND_net), .O(n2031));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(current[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5712));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(current[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5720));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_2139 (.I0(n2026), .I1(n2025), .I2(n2028), .I3(GND_net), 
            .O(n61426));
    defparam i1_3_lut_adj_2139.LUT_INIT = 16'hfefe;
    SB_LUT4 i16207_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5966[6]), 
            .I2(n42804), .I3(n25540), .O(n30215));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16207_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2140 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [1]), 
            .O(n56836));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2140.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(current[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5719));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(current[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5718));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_2141 (.I0(n2023), .I1(n2024), .I2(n2027), .I3(GND_net), 
            .O(n61428));
    defparam i1_3_lut_adj_2141.LUT_INIT = 16'hfefe;
    SB_LUT4 i16208_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5966[7]), 
            .I2(n42804), .I3(n25535), .O(n30216));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16208_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_2_lut_adj_2142 (.I0(state[0]), .I1(n23_adj_5913), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5815));
    defparam i1_2_lut_adj_2142.LUT_INIT = 16'h2222;
    SB_LUT4 i13_4_lut (.I0(n111), .I1(n43462), .I2(state[1]), .I3(n4_adj_5815), 
            .O(n5_adj_5904));   // verilog/neopixel.v(34[12] 116[6])
    defparam i13_4_lut.LUT_INIT = 16'hcafa;
    SB_LUT4 i12_4_lut_adj_2143 (.I0(\data_in_frame[19] [1]), .I1(n28379), 
            .I2(n28434), .I3(rx_data[1]), .O(n56053));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2143.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2144 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [2]), 
            .O(n56837));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2144.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2145 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [3]), 
            .O(n56838));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2145.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2146 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [4]), 
            .O(n56839));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2146.LUT_INIT = 16'h2300;
    SB_LUT4 i12_4_lut_adj_2147 (.I0(\data_in_frame[19] [0]), .I1(n28379), 
            .I2(n28434), .I3(rx_data[0]), .O(n56057));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2147.LUT_INIT = 16'h3a0a;
    SB_LUT4 i28319_4_lut_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15_adj_5681), .I3(n15), .O(n42234));
    defparam i28319_4_lut_4_lut.LUT_INIT = 16'hf535;
    SB_LUT4 i12_4_lut_adj_2148 (.I0(\data_in_frame[18] [7]), .I1(n28381), 
            .I2(n28436), .I3(rx_data[7]), .O(n56061));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2148.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_2149 (.I0(\data_in_frame[18] [6]), .I1(n28381), 
            .I2(n28436), .I3(rx_data[6]), .O(n56065));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2149.LUT_INIT = 16'h3a0a;
    SB_LUT4 i15724_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[1] [2]), 
            .I3(control_mode[2]), .O(n29732));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15724_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2150 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [5]), 
            .O(n56840));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2150.LUT_INIT = 16'h2300;
    SB_LUT4 i12_4_lut_adj_2151 (.I0(\data_in_frame[18] [2]), .I1(n28381), 
            .I2(n28436), .I3(rx_data[2]), .O(n56071));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2151.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2152 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [6]), 
            .O(n56772));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2152.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2153 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [7]), 
            .O(n56782));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2153.LUT_INIT = 16'h2300;
    SB_LUT4 i12_4_lut_adj_2154 (.I0(\data_in_frame[18] [1]), .I1(n28381), 
            .I2(n28436), .I3(rx_data[1]), .O(n56075));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2154.LUT_INIT = 16'h3a0a;
    SB_LUT4 LessThan_14_i15_2_lut (.I0(current[7]), .I1(current_limit[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5660));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i13_2_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16731_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [1]), 
            .O(n30739));   // verilog/coms.v(130[12] 305[6])
    defparam i16731_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i46831_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n62508));
    defparam i46831_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53423_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n6617), .I2(n62508), 
            .I3(n25_adj_5897), .O(n17_adj_5896));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i53423_4_lut.LUT_INIT = 16'h88ba;
    SB_LUT4 encoder0_position_30__I_0_i971_3_lut (.I0(n1424), .I1(n1491), 
            .I2(n1455), .I3(GND_net), .O(n1523));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16188_3_lut (.I0(\data_in_frame[13] [6]), .I1(rx_data[6]), 
            .I2(n59230), .I3(GND_net), .O(n30196));   // verilog/coms.v(130[12] 305[6])
    defparam i16188_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16184_3_lut (.I0(\data_in_frame[13] [5]), .I1(rx_data[5]), 
            .I2(n59230), .I3(GND_net), .O(n30192));   // verilog/coms.v(130[12] 305[6])
    defparam i16184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i969_3_lut (.I0(n1422), .I1(n1489), 
            .I2(n1455), .I3(GND_net), .O(n1521));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i969_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16181_3_lut (.I0(\data_in_frame[13] [4]), .I1(rx_data[4]), 
            .I2(n59230), .I3(GND_net), .O(n30189));   // verilog/coms.v(130[12] 305[6])
    defparam i16181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16178_3_lut (.I0(\data_in_frame[13] [3]), .I1(rx_data[3]), 
            .I2(n59230), .I3(GND_net), .O(n30186));   // verilog/coms.v(130[12] 305[6])
    defparam i16178_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5762));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i977_3_lut (.I0(n1430), .I1(n1497), 
            .I2(n1455), .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i19_2_lut (.I0(current[9]), .I1(current_limit[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16174_3_lut (.I0(\data_in_frame[13] [2]), .I1(rx_data[2]), 
            .I2(n59230), .I3(GND_net), .O(n30182));   // verilog/coms.v(130[12] 305[6])
    defparam i16174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16171_3_lut (.I0(\data_in_frame[13] [1]), .I1(rx_data[1]), 
            .I2(n59230), .I3(GND_net), .O(n30179));   // verilog/coms.v(130[12] 305[6])
    defparam i16171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1044_3_lut (.I0(n1529), .I1(n1596), 
            .I2(n1554), .I3(GND_net), .O(n1628));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i7_2_lut (.I0(current[3]), .I1(current_limit[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5661));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i1111_3_lut (.I0(n1628), .I1(n1695), 
            .I2(n1653), .I3(GND_net), .O(n1727));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16168_3_lut (.I0(\data_in_frame[13] [0]), .I1(rx_data[0]), 
            .I2(n59230), .I3(GND_net), .O(n30176));   // verilog/coms.v(130[12] 305[6])
    defparam i16168_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i9_2_lut (.I0(current[4]), .I1(current_limit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i11_2_lut (.I0(current[5]), .I1(current_limit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16164_3_lut (.I0(\data_in_frame[12] [7]), .I1(rx_data[7]), 
            .I2(n57921), .I3(GND_net), .O(n30172));   // verilog/coms.v(130[12] 305[6])
    defparam i16164_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16161_3_lut (.I0(\data_in_frame[12] [6]), .I1(rx_data[6]), 
            .I2(n57921), .I3(GND_net), .O(n30169));   // verilog/coms.v(130[12] 305[6])
    defparam i16161_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1178_3_lut (.I0(n1727), .I1(n1794_adj_5807), 
            .I2(n1752), .I3(GND_net), .O(n1826));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1178_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16158_3_lut (.I0(\data_in_frame[12] [5]), .I1(rx_data[5]), 
            .I2(n57921), .I3(GND_net), .O(n30166));   // verilog/coms.v(130[12] 305[6])
    defparam i16158_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1245_3_lut (.I0(n1826), .I1(n1893), 
            .I2(n1851), .I3(GND_net), .O(n1925));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1245_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1312_3_lut (.I0(n1925), .I1(n1992), 
            .I2(n1950), .I3(GND_net), .O(n2024));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i52640_3_lut (.I0(rx_data[4]), .I1(\data_in_frame[12] [4]), 
            .I2(n57921), .I3(GND_net), .O(n56343));   // verilog/coms.v(94[13:20])
    defparam i52640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52639_3_lut (.I0(rx_data[3]), .I1(\data_in_frame[12] [3]), 
            .I2(n57921), .I3(GND_net), .O(n56303));   // verilog/coms.v(94[13:20])
    defparam i52639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15725_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[1] [3]), 
            .I3(control_mode[3]), .O(n29733));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15725_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 encoder0_position_30__I_0_i976_3_lut (.I0(n1429), .I1(n1496), 
            .I2(n1455), .I3(GND_net), .O(n1528));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16148_3_lut (.I0(\data_in_frame[12] [2]), .I1(rx_data[2]), 
            .I2(n57921), .I3(GND_net), .O(n30156));   // verilog/coms.v(130[12] 305[6])
    defparam i16148_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7_4_lut_adj_2155 (.I0(dti_counter[0]), .I1(n14_adj_5901), .I2(n10_adj_5902), 
            .I3(dti_counter[3]), .O(n22849));   // verilog/TinyFPGA_B.v(171[9:23])
    defparam i7_4_lut_adj_2155.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i1043_3_lut (.I0(n1528), .I1(n1595), 
            .I2(n1554), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(duty[2]), .I1(duty[3]), .I2(current[3]), 
            .I3(GND_net), .O(n6_adj_5725));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_14_i17_2_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16144_3_lut (.I0(\data_in_frame[12] [1]), .I1(rx_data[1]), 
            .I2(n57921), .I3(GND_net), .O(n30152));   // verilog/coms.v(130[12] 305[6])
    defparam i16144_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i5_2_lut (.I0(current[2]), .I1(current_limit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5663));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_30__I_0_i1110_3_lut (.I0(n1627), .I1(n1694), 
            .I2(n1653), .I3(GND_net), .O(n1726));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i50568_4_lut (.I0(n11), .I1(n9), .I2(n7_adj_5661), .I3(n5_adj_5663), 
            .O(n66254));
    defparam i50568_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 encoder0_position_30__I_0_i1177_3_lut (.I0(n1726), .I1(n1793), 
            .I2(n1752), .I3(GND_net), .O(n1825));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1244_3_lut (.I0(n1825), .I1(n1892), 
            .I2(n1851), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1244_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1311_3_lut (.I0(n1924), .I1(n1991), 
            .I2(n1950), .I3(GND_net), .O(n2023));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16141_3_lut (.I0(\data_in_frame[12] [0]), .I1(rx_data[0]), 
            .I2(n57921), .I3(GND_net), .O(n30149));   // verilog/coms.v(130[12] 305[6])
    defparam i16141_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i16_3_lut (.I0(n8), .I1(current_limit[9]), .I2(n19), 
            .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_14_i4_4_lut (.I0(current_limit[0]), .I1(current_limit[1]), 
            .I2(current[1]), .I3(current[0]), .O(n4_adj_5664));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i52075_3_lut (.I0(n4_adj_5664), .I1(current_limit[5]), .I2(n11), 
            .I3(GND_net), .O(n67761));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i52075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2156 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [0]), 
            .O(n56841));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2156.LUT_INIT = 16'h2300;
    SB_LUT4 i52076_3_lut (.I0(n67761), .I1(current_limit[6]), .I2(n13), 
            .I3(GND_net), .O(n67762));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i52076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2157 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [1]), 
            .O(n56842));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2157.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2158 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [2]), 
            .O(n56843));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2158.LUT_INIT = 16'h2300;
    SB_LUT4 i50547_4_lut (.I0(n17), .I1(n15_adj_5660), .I2(n13), .I3(n66254), 
            .O(n66233));
    defparam i50547_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i16331_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[21] [1]), 
            .I3(current_limit[1]), .O(n30339));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i16331_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i52413_4_lut (.I0(n16), .I1(n6_adj_5662), .I2(n19), .I3(n66231), 
            .O(n68099));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i52413_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50817_3_lut (.I0(n67762), .I1(current_limit[7]), .I2(n15_adj_5660), 
            .I3(GND_net), .O(n66503));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i50817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52569_4_lut (.I0(n66503), .I1(n68099), .I2(n19), .I3(n66233), 
            .O(n68255));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i52569_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52570_3_lut (.I0(n68255), .I1(current_limit[10]), .I2(current[10]), 
            .I3(GND_net), .O(n68256));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i52570_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2159 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [3]), 
            .O(n56844));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2159.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2160 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [7]), 
            .O(n56918));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2160.LUT_INIT = 16'h2300;
    SB_LUT4 i52496_3_lut (.I0(n68256), .I1(current_limit[11]), .I2(current[11]), 
            .I3(GND_net), .O(n68182));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam i52496_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_14_i26_3_lut (.I0(n68182), .I1(current_limit[12]), 
            .I2(current[15]), .I3(GND_net), .O(n26));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i15631_3_lut_4_lut (.I0(n2873), .I1(n27696), .I2(\data_in_frame[21] [0]), 
            .I3(current_limit[0]), .O(n29639));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i15631_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2161 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [0]), 
            .O(n56917));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2161.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2162 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [1]), 
            .O(n56916));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2162.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_11_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(current[6]), 
            .I3(GND_net), .O(n10_adj_5721));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2163 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [2]), 
            .O(n56915));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2163.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(duty[7]), .I1(n303), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5680));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2164 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [4]), 
            .O(n56845));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2164.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2165 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [5]), 
            .O(n56846));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2165.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(duty[6]), .I1(n304), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5685));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(duty[9]), .I1(n301), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5667));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i7_2_lut (.I0(duty[3]), .I1(n307), .I2(GND_net), 
            .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(duty[5]), .I1(n305), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5682));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i9_2_lut (.I0(duty[4]), .I1(n306), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5665));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(duty[8]), .I1(n302), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5668));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2166 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [6]), 
            .O(n56847));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2166.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2167 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [7]), 
            .O(n56848));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2167.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_11_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(current[8]), 
            .I3(GND_net), .O(n8_adj_5723));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_17_i5_2_lut (.I0(duty[2]), .I1(n308), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50311_4_lut (.I0(n11_adj_5682), .I1(n9_adj_5665), .I2(n7), 
            .I3(n5), .O(n65997));
    defparam i50311_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2168 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [3]), 
            .O(n56776));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2168.LUT_INIT = 16'h2300;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5763));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16087_3_lut (.I0(\data_in_frame[9] [7]), .I1(rx_data[7]), .I2(n57039), 
            .I3(GND_net), .O(n30095));   // verilog/coms.v(130[12] 305[6])
    defparam i16087_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_17_i8_3_lut (.I0(n306), .I1(n302), .I2(n17_adj_5668), 
            .I3(GND_net), .O(n8_adj_5666));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16084_3_lut (.I0(\data_in_frame[9] [6]), .I1(rx_data[6]), .I2(n57039), 
            .I3(GND_net), .O(n30092));   // verilog/coms.v(130[12] 305[6])
    defparam i16084_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2169 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [4]), 
            .O(n56914));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2169.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i6_3_lut (.I0(n308), .I1(n307), .I2(n7), .I3(GND_net), 
            .O(n6_adj_5659));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n8_adj_5666), .I1(n301), .I2(n19_adj_5667), 
            .I3(GND_net), .O(n16_adj_5669));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2170 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [5]), 
            .O(n56913));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2170.LUT_INIT = 16'h2300;
    SB_LUT4 i16081_3_lut (.I0(\data_in_frame[9] [5]), .I1(rx_data[5]), .I2(n57039), 
            .I3(GND_net), .O(n30089));   // verilog/coms.v(130[12] 305[6])
    defparam i16081_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_adj_2171 (.I0(duty[15]), .I1(duty[20]), .I2(n294), 
            .I3(GND_net), .O(n12_adj_5791));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i2_3_lut_adj_2171.LUT_INIT = 16'h7e7e;
    SB_LUT4 i6_4_lut_adj_2172 (.I0(duty[13]), .I1(n12_adj_5791), .I2(duty[21]), 
            .I3(n294), .O(n16_adj_5789));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i6_4_lut_adj_2172.LUT_INIT = 16'hdffe;
    SB_LUT4 i16077_3_lut (.I0(\data_in_frame[9] [4]), .I1(rx_data[4]), .I2(n57039), 
            .I3(GND_net), .O(n30085));   // verilog/coms.v(130[12] 305[6])
    defparam i16077_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_3_lut (.I0(duty[19]), .I1(duty[16]), .I2(n294), .I3(GND_net), 
            .O(n14_adj_5790));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i4_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i16074_3_lut (.I0(\data_in_frame[9] [3]), .I1(rx_data[3]), .I2(n57039), 
            .I3(GND_net), .O(n30082));   // verilog/coms.v(130[12] 305[6])
    defparam i16074_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16071_3_lut (.I0(\data_in_frame[9] [2]), .I1(rx_data[2]), .I2(n57039), 
            .I3(GND_net), .O(n30079));   // verilog/coms.v(130[12] 305[6])
    defparam i16071_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1237_3_lut (.I0(n1818), .I1(n1885), 
            .I2(n1851), .I3(GND_net), .O(n1917));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1237_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1304_3_lut (.I0(n1917), .I1(n1984), 
            .I2(n1950), .I3(GND_net), .O(n2016));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1304_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_4_lut_adj_2173 (.I0(\FRAME_MATCHER.i [3]), .I1(n57917), 
            .I2(n8_adj_5760), .I3(n134), .O(n92));
    defparam i2_3_lut_4_lut_adj_2173.LUT_INIT = 16'hfffb;
    SB_LUT4 LessThan_17_i10_3_lut (.I0(n305), .I1(n304), .I2(n13_adj_5685), 
            .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16067_3_lut (.I0(\data_in_frame[9] [1]), .I1(rx_data[1]), .I2(n57039), 
            .I3(GND_net), .O(n30075));   // verilog/coms.v(130[12] 305[6])
    defparam i16067_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2174 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [6]), 
            .O(n56912));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2174.LUT_INIT = 16'h2300;
    SB_LUT4 i16064_3_lut (.I0(\data_in_frame[9] [0]), .I1(rx_data[0]), .I2(n57039), 
            .I3(GND_net), .O(n30072));   // verilog/coms.v(130[12] 305[6])
    defparam i16064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5764));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_17_i4_3_lut (.I0(n65285), .I1(n309), .I2(duty[1]), 
            .I3(GND_net), .O(n4));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2175 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [7]), 
            .O(n56911));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2175.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i12_3_lut (.I0(n10), .I1(n303), .I2(n15_adj_5680), 
            .I3(GND_net), .O(n12_adj_5738));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam LessThan_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16061_3_lut (.I0(\data_in_frame[8] [7]), .I1(rx_data[7]), .I2(n57948), 
            .I3(GND_net), .O(n30069));   // verilog/coms.v(130[12] 305[6])
    defparam i16061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16058_3_lut (.I0(\data_in_frame[8] [6]), .I1(rx_data[6]), .I2(n57948), 
            .I3(GND_net), .O(n30066));   // verilog/coms.v(130[12] 305[6])
    defparam i16058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6572_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_400));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i6572_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 i50299_4_lut (.I0(n17_adj_5668), .I1(n15_adj_5680), .I2(n13_adj_5685), 
            .I3(n65997), .O(n65985));
    defparam i50299_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52411_4_lut (.I0(n16_adj_5669), .I1(n6_adj_5659), .I2(n19_adj_5667), 
            .I3(n65983), .O(n68097));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i52411_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51559_4_lut (.I0(n12_adj_5738), .I1(n4), .I2(n15_adj_5680), 
            .I3(n65995), .O(n67245));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51559_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i16055_3_lut (.I0(\data_in_frame[8] [5]), .I1(rx_data[5]), .I2(n57948), 
            .I3(GND_net), .O(n30063));   // verilog/coms.v(130[12] 305[6])
    defparam i16055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6570_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_391));   // verilog/TinyFPGA_B.v(200[7] 219[14])
    defparam i6570_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 i52576_4_lut (.I0(n67245), .I1(n68097), .I2(n19_adj_5667), 
            .I3(n65985), .O(n68262));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i52576_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52577_3_lut (.I0(n68262), .I1(n300), .I2(duty[10]), .I3(GND_net), 
            .O(n68263));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i52577_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i23858_3_lut (.I0(n57948), .I1(rx_data[4]), .I2(\data_in_frame[8] [4]), 
            .I3(GND_net), .O(n30280));   // verilog/coms.v(94[13:20])
    defparam i23858_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i52488_3_lut (.I0(n68263), .I1(n299), .I2(duty[11]), .I3(GND_net), 
            .O(n68174));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i52488_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2176 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [0]), 
            .O(n56910));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2176.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2177 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [1]), 
            .O(n56909));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2177.LUT_INIT = 16'h2300;
    SB_LUT4 i6562_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_355));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i6562_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 i16049_3_lut (.I0(\data_in_frame[8] [3]), .I1(rx_data[3]), .I2(n57948), 
            .I3(GND_net), .O(n30057));   // verilog/coms.v(130[12] 305[6])
    defparam i16049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16046_3_lut (.I0(\data_in_frame[8] [2]), .I1(rx_data[2]), .I2(n57948), 
            .I3(GND_net), .O(n30054));   // verilog/coms.v(130[12] 305[6])
    defparam i16046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16042_3_lut (.I0(\data_in_frame[8] [1]), .I1(rx_data[1]), .I2(n57948), 
            .I3(GND_net), .O(n30050));   // verilog/coms.v(130[12] 305[6])
    defparam i16042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8_4_lut (.I0(duty[14]), .I1(n16_adj_5789), .I2(duty[18]), 
            .I3(n294), .O(n18_adj_5787));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i8_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 i7_4_lut_adj_2178 (.I0(duty[22]), .I1(n14_adj_5790), .I2(duty[17]), 
            .I3(n294), .O(n17_adj_5788));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i7_4_lut_adj_2178.LUT_INIT = 16'hdffe;
    SB_LUT4 i6564_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_372));   // verilog/TinyFPGA_B.v(179[7] 198[15])
    defparam i6564_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 i16039_3_lut (.I0(\data_in_frame[8] [0]), .I1(rx_data[0]), .I2(n57948), 
            .I3(GND_net), .O(n30047));   // verilog/coms.v(130[12] 305[6])
    defparam i16039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6566_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_377));
    defparam i6566_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 i51884_3_lut (.I0(n68174), .I1(n298), .I2(duty[12]), .I3(GND_net), 
            .O(n67570));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51884_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i6568_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_386));
    defparam i6568_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 i51885_4_lut (.I0(n67570), .I1(n294), .I2(n17_adj_5788), .I3(n18_adj_5787), 
            .O(n67571));   // verilog/TinyFPGA_B.v(121[11:24])
    defparam i51885_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i42401_4_lut (.I0(n260), .I1(duty[23]), .I2(n294), .I3(n67571), 
            .O(n11577));
    defparam i42401_4_lut.LUT_INIT = 16'h1151;
    SB_LUT4 i51357_3_lut (.I0(n15_adj_5718), .I1(n13_adj_5719), .I2(n11_adj_5720), 
            .I3(GND_net), .O(n67043));
    defparam i51357_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_2179 (.I0(\FRAME_MATCHER.i [3]), .I1(n3470), 
            .I2(n161), .I3(n134), .O(n111_adj_5814));
    defparam i1_2_lut_3_lut_4_lut_adj_2179.LUT_INIT = 16'hffbf;
    SB_LUT4 i50309_2_lut_4_lut (.I0(duty[6]), .I1(n304), .I2(duty[5]), 
            .I3(n305), .O(n65995));
    defparam i50309_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51309_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n67043), .O(n66995));
    defparam i51309_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i50458_4_lut (.I0(n21_adj_5712), .I1(n19_adj_5713), .I2(n17_adj_5716), 
            .I3(n9_adj_5722), .O(n66144));
    defparam i50458_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mux_245_i1_4_lut (.I0(encoder1_position_scaled[0]), .I1(displacement[0]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[0]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i50297_2_lut_4_lut (.I0(duty[8]), .I1(n302), .I2(duty[4]), 
            .I3(n306), .O(n65983));
    defparam i50297_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51381_4_lut (.I0(n9_adj_5722), .I1(n7_adj_5724), .I2(current[2]), 
            .I3(duty[2]), .O(n67067));
    defparam i51381_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 mux_245_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[1]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i51791_4_lut (.I0(n15_adj_5718), .I1(n13_adj_5719), .I2(n11_adj_5720), 
            .I3(n67067), .O(n67477));
    defparam i51791_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51789_4_lut (.I0(n21_adj_5712), .I1(n19_adj_5713), .I2(n17_adj_5716), 
            .I3(n67477), .O(n67475));
    defparam i51789_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52339_4_lut (.I0(current[15]), .I1(n23_adj_5711), .I2(duty[12]), 
            .I3(n67475), .O(n68025));
    defparam i52339_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i51331_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n68025), .O(n67017));
    defparam i51331_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(current[1]), 
            .I3(current[0]), .O(n4_adj_5726));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i51263_4_lut (.I0(current[15]), .I1(duty[16]), .I2(duty[17]), 
            .I3(n15_adj_5718), .O(n66949));
    defparam i51263_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 LessThan_11_i30_4_lut (.I0(duty[7]), .I1(duty[17]), .I2(current[15]), 
            .I3(duty[16]), .O(n30_adj_5710));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i30_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i52071_3_lut (.I0(n4_adj_5726), .I1(duty[13]), .I2(current[15]), 
            .I3(GND_net), .O(n67757));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52071_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50382_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n66995), .O(n66068));
    defparam i50382_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 LessThan_11_i35_rep_172_2_lut (.I0(current[15]), .I1(duty[17]), 
            .I2(GND_net), .I3(GND_net), .O(n69682));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i35_rep_172_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52415_3_lut (.I0(n30_adj_5710), .I1(n10_adj_5721), .I2(n66949), 
            .I3(GND_net), .O(n68101));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52415_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_14_i6_3_lut_3_lut (.I0(current_limit[2]), .I1(current_limit[3]), 
            .I2(current[3]), .I3(GND_net), .O(n6_adj_5662));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50545_2_lut_4_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(current[4]), .I3(current_limit[4]), .O(n66231));
    defparam i50545_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_14_i8_3_lut_3_lut (.I0(current_limit[4]), .I1(current_limit[8]), 
            .I2(current[8]), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(118[9:30])
    defparam LessThan_14_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50825_4_lut (.I0(n67757), .I1(duty[15]), .I2(current[15]), 
            .I3(duty[14]), .O(n66511));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i50825_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i52041_3_lut (.I0(n6_adj_5725), .I1(duty[10]), .I2(n21_adj_5712), 
            .I3(GND_net), .O(n67727));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52042_3_lut (.I0(n67727), .I1(duty[11]), .I2(n23_adj_5711), 
            .I3(GND_net), .O(n67728));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_245_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[2]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i51785_4_lut (.I0(current[15]), .I1(n23_adj_5711), .I2(duty[12]), 
            .I3(n66144), .O(n67471));
    defparam i51785_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n8_adj_5723), .I1(duty[9]), .I2(n19_adj_5713), 
            .I3(GND_net), .O(n16_adj_5717));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16213_4_lut_4_lut (.I0(n27920), .I1(state[1]), .I2(bit_ctr[1]), 
            .I3(bit_ctr[0]), .O(n30221));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16213_4_lut_4_lut.LUT_INIT = 16'h5270;
    SB_LUT4 i50827_3_lut (.I0(n67728), .I1(duty[12]), .I2(current[15]), 
            .I3(GND_net), .O(n66513));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i50827_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52101_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n67017), .O(n67787));
    defparam i52101_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i15532_3_lut_4_lut (.I0(\data_in_frame[18] [3]), .I1(rx_data[3]), 
            .I2(n40973), .I3(n8_adj_5741), .O(n29540));   // verilog/coms.v(130[12] 305[6])
    defparam i15532_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i15535_3_lut_4_lut (.I0(\data_in_frame[18] [4]), .I1(rx_data[4]), 
            .I2(n40973), .I3(n8_adj_5741), .O(n29543));   // verilog/coms.v(130[12] 305[6])
    defparam i15535_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i15538_3_lut_4_lut (.I0(\data_in_frame[18] [5]), .I1(rx_data[5]), 
            .I2(n40973), .I3(n8_adj_5741), .O(n29546));   // verilog/coms.v(130[12] 305[6])
    defparam i15538_3_lut_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5775));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5776));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52571_4_lut (.I0(n66511), .I1(n68101), .I2(n69682), .I3(n66068), 
            .O(n68257));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52571_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i51571_3_lut (.I0(n66513), .I1(n16_adj_5717), .I2(n67471), 
            .I3(GND_net), .O(n67257));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i51571_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i52633_4_lut (.I0(n67257), .I1(n68257), .I2(n69682), .I3(n67787), 
            .O(n68319));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52633_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52626_4_lut (.I0(n68319), .I1(duty[19]), .I2(current[15]), 
            .I3(duty[18]), .O(n68312));   // verilog/TinyFPGA_B.v(110[10:22])
    defparam i52626_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i1_4_lut_adj_2180 (.I0(n68312), .I1(current[15]), .I2(duty[21]), 
            .I3(duty[20]), .O(n5_adj_5905));
    defparam i1_4_lut_adj_2180.LUT_INIT = 16'hfffe;
    SB_LUT4 i15987_3_lut (.I0(\data_in_frame[5] [7]), .I1(rx_data[7]), .I2(n59242), 
            .I3(GND_net), .O(n29995));   // verilog/coms.v(130[12] 305[6])
    defparam i15987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7_4_lut_adj_2181 (.I0(n5_adj_5905), .I1(duty[23]), .I2(n21_adj_5850), 
            .I3(duty[22]), .O(n11579));
    defparam i7_4_lut_adj_2181.LUT_INIT = 16'h3332;
    SB_LUT4 i15858_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n60804), 
            .I3(n27_adj_5781), .O(n29866));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i15858_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16297_3_lut (.I0(\data_in_frame[13] [7]), .I1(rx_data[7]), 
            .I2(n59230), .I3(GND_net), .O(n30305));   // verilog/coms.v(130[12] 305[6])
    defparam i16297_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5777));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16300_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30308));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16300_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5778));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_2182 (.I0(n40973), .I1(n8_adj_5741), .I2(GND_net), 
            .I3(GND_net), .O(n28436));
    defparam i1_2_lut_adj_2182.LUT_INIT = 16'h2222;
    SB_LUT4 i50285_2_lut_4_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n57917), 
            .I2(n134), .I3(n8_adj_5731), .O(n65433));   // verilog/coms.v(94[13:20])
    defparam i50285_2_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 mux_4310_i27_3_lut (.I0(encoder0_position[26]), .I1(n6_adj_5707), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n625));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_2183 (.I0(\data_in_frame[18] [0]), .I1(n28381), 
            .I2(n28436), .I3(rx_data[0]), .O(n56079));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2183.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5779));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[4]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_4_lut (.I0(n92), .I1(\data_in_frame[16] [7]), .I2(reset), 
            .I3(rx_data[7]), .O(n56249));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hcdc8;
    SB_LUT4 i12_4_lut_adj_2184 (.I0(\data_in_frame[17] [7]), .I1(n28387), 
            .I2(n28438), .I3(rx_data[7]), .O(n56083));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2184.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_2185 (.I0(\data_in_frame[17] [6]), .I1(n28387), 
            .I2(n28438), .I3(rx_data[6]), .O(n56087));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2185.LUT_INIT = 16'h3a0a;
    SB_LUT4 mux_4310_i28_3_lut (.I0(encoder0_position[27]), .I1(n5_adj_5709), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n516));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16733_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [3]), 
            .O(n30741));   // verilog/coms.v(130[12] 305[6])
    defparam i16733_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16307_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30315));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i29_3_lut (.I0(encoder0_position[28]), .I1(n4_adj_5714), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n623));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16308_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30316));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2186 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5684));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_4_lut_adj_2186.LUT_INIT = 16'h7bde;
    SB_LUT4 i16309_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30317));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i30_3_lut (.I0(encoder0_position[29]), .I1(n3), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n622));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16310_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30318));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16311_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30319));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6055_2_lut (.I0(n2_adj_5715), .I1(encoder0_position[30]), .I2(GND_net), 
            .I3(GND_net), .O(n621));
    defparam i6055_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_245_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[5]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_245_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[7]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16312_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30320));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16313_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30321));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(262[11:14])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1444_3_lut (.I0(n2121), .I1(n2188), 
            .I2(n2148), .I3(GND_net), .O(n2220));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16314_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30322));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16315_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n25_adj_5906), .I3(GND_net), .O(n30323));   // verilog/neopixel.v(34[12] 116[6])
    defparam i16315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15984_3_lut (.I0(\data_in_frame[5] [6]), .I1(rx_data[6]), .I2(n59242), 
            .I3(GND_net), .O(n29992));   // verilog/coms.v(130[12] 305[6])
    defparam i15984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15981_3_lut (.I0(\data_in_frame[5] [5]), .I1(rx_data[5]), .I2(n59242), 
            .I3(GND_net), .O(n29989));   // verilog/coms.v(130[12] 305[6])
    defparam i15981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_1083_i9_2_lut (.I0(r_Clock_Count[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5831));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1083_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15978_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n59242), 
            .I3(GND_net), .O(n29986));   // verilog/coms.v(130[12] 305[6])
    defparam i15978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15841_3_lut_4_lut (.I0(deadband[2]), .I1(\data_in_frame[16] [2]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29849));   // verilog/coms.v(130[12] 305[6])
    defparam i15841_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_3_lut_adj_2187 (.I0(n5_adj_5894), .I1(n3), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n61420));
    defparam i1_3_lut_adj_2187.LUT_INIT = 16'h8080;
    SB_LUT4 i12_4_lut_adj_2188 (.I0(\data_in_frame[17] [5]), .I1(n28387), 
            .I2(n28438), .I3(rx_data[5]), .O(n56091));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2188.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_2189 (.I0(\data_in_frame[17] [4]), .I1(n28387), 
            .I2(n28438), .I3(rx_data[4]), .O(n56095));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2189.LUT_INIT = 16'h3a0a;
    SB_LUT4 i15859_3_lut (.I0(\data_in_frame[1] [1]), .I1(rx_data[1]), .I2(n57044), 
            .I3(GND_net), .O(n29867));   // verilog/coms.v(130[12] 305[6])
    defparam i15859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22792_3_lut (.I0(n214), .I1(IntegralLimit[17]), .I2(n155), 
            .I3(GND_net), .O(n36759));
    defparam i22792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_2190 (.I0(n36759), .I1(Ki[0]), .I2(GND_net), 
            .I3(GND_net), .O(n53));
    defparam i1_2_lut_adj_2190.LUT_INIT = 16'h8888;
    SB_LUT4 i15862_3_lut (.I0(\data_in_frame[1] [2]), .I1(rx_data[2]), .I2(n57044), 
            .I3(GND_net), .O(n29870));   // verilog/coms.v(130[12] 305[6])
    defparam i15862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15840_3_lut_4_lut (.I0(deadband[3]), .I1(\data_in_frame[16] [3]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29848));   // verilog/coms.v(130[12] 305[6])
    defparam i15840_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 LessThan_1083_i4_4_lut (.I0(r_Clock_Count[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5828));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1083_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 encoder0_position_30__I_0_i500_4_lut (.I0(n2_adj_5715), .I1(n7450), 
            .I2(n61420), .I3(encoder0_position[30]), .O(n828));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i500_4_lut.LUT_INIT = 16'h8a80;
    SB_LUT4 i15839_3_lut_4_lut (.I0(deadband[4]), .I1(\data_in_frame[16] [4]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29847));   // verilog/coms.v(130[12] 305[6])
    defparam i15839_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i12_4_lut_adj_2191 (.I0(\data_in_frame[17] [3]), .I1(n28387), 
            .I2(n28438), .I3(rx_data[3]), .O(n56099));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2191.LUT_INIT = 16'h3a0a;
    SB_LUT4 i15838_3_lut_4_lut (.I0(deadband[5]), .I1(\data_in_frame[16] [5]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29846));   // verilog/coms.v(130[12] 305[6])
    defparam i15838_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i12_4_lut_adj_2192 (.I0(\data_in_frame[17] [2]), .I1(n28387), 
            .I2(n28438), .I3(rx_data[2]), .O(n56101));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2192.LUT_INIT = 16'h3a0a;
    SB_LUT4 LessThan_1083_i8_3_lut (.I0(n6_adj_5829), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5831), .I3(GND_net), .O(n8_adj_5830));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1083_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_2193 (.I0(\data_in_frame[17] [1]), .I1(n28387), 
            .I2(n28438), .I3(rx_data[1]), .O(n56103));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2193.LUT_INIT = 16'h3a0a;
    SB_LUT4 i52387_4_lut (.I0(n8_adj_5830), .I1(n4_adj_5828), .I2(n9_adj_5831), 
            .I3(n66181), .O(n68073));   // verilog/uart_rx.v(119[17:57])
    defparam i52387_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i12_4_lut_adj_2194 (.I0(\data_in_frame[17] [0]), .I1(n28387), 
            .I2(n28438), .I3(rx_data[0]), .O(n56107));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2194.LUT_INIT = 16'h3a0a;
    SB_LUT4 i12_4_lut_adj_2195 (.I0(n56988), .I1(\data_in_frame[16] [2]), 
            .I2(n142), .I3(rx_data[2]), .O(n56199));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2195.LUT_INIT = 16'hcac0;
    SB_LUT4 mux_245_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[8]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12_4_lut_adj_2196 (.I0(n56988), .I1(\data_in_frame[16] [1]), 
            .I2(n142), .I3(rx_data[1]), .O(n56201));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2196.LUT_INIT = 16'hcac0;
    SB_LUT4 i15974_3_lut (.I0(\data_in_frame[5] [3]), .I1(rx_data[3]), .I2(n59242), 
            .I3(GND_net), .O(n29982));   // verilog/coms.v(130[12] 305[6])
    defparam i15974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29496_3_lut (.I0(n945), .I1(n2032), .I2(n2033), .I3(GND_net), 
            .O(n43402));
    defparam i29496_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i15971_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n59242), 
            .I3(GND_net), .O(n29979));   // verilog/coms.v(130[12] 305[6])
    defparam i15971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15968_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n59242), 
            .I3(GND_net), .O(n29976));   // verilog/coms.v(130[12] 305[6])
    defparam i15968_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2197 (.I0(reset), .I1(n92), .I2(GND_net), .I3(GND_net), 
            .O(n142));
    defparam i1_2_lut_adj_2197.LUT_INIT = 16'heeee;
    SB_LUT4 i52388_3_lut (.I0(n68073), .I1(o_Rx_DV_N_3488[5]), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n68074));   // verilog/uart_rx.v(119[17:57])
    defparam i52388_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52251_3_lut (.I0(n68074), .I1(o_Rx_DV_N_3488[6]), .I2(r_Clock_Count[6]), 
            .I3(GND_net), .O(n67937));   // verilog/uart_rx.v(119[17:57])
    defparam i52251_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50990_3_lut (.I0(n67937), .I1(o_Rx_DV_N_3488[7]), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(n4937));   // verilog/uart_rx.v(119[17:57])
    defparam i50990_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5780));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15965_3_lut (.I0(\data_in_frame[5] [0]), .I1(rx_data[0]), .I2(n59242), 
            .I3(GND_net), .O(n29973));   // verilog/coms.v(130[12] 305[6])
    defparam i15965_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[9]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_245_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[18]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_1584_i1_3_lut (.I0(duty[3]), .I1(duty[0]), .I2(n260), 
            .I3(GND_net), .O(n11642));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1584_i2_3_lut (.I0(duty[4]), .I1(duty[1]), .I2(n260), 
            .I3(GND_net), .O(n12224));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[10]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_30__I_0_i1443_3_lut (.I0(n2120), .I1(n2187), 
            .I2(n2148), .I3(GND_net), .O(n2219));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15837_3_lut_4_lut (.I0(deadband[6]), .I1(\data_in_frame[16] [6]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29845));   // verilog/coms.v(130[12] 305[6])
    defparam i15837_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15836_3_lut_4_lut (.I0(deadband[7]), .I1(\data_in_frame[16] [7]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29844));   // verilog/coms.v(130[12] 305[6])
    defparam i15836_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15835_3_lut_4_lut (.I0(deadband[8]), .I1(\data_in_frame[15] [0]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29843));   // verilog/coms.v(130[12] 305[6])
    defparam i15835_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15834_3_lut_4_lut (.I0(deadband[9]), .I1(\data_in_frame[15] [1]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29842));   // verilog/coms.v(130[12] 305[6])
    defparam i15834_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15833_3_lut_4_lut (.I0(deadband[10]), .I1(\data_in_frame[15] [2]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29841));   // verilog/coms.v(130[12] 305[6])
    defparam i15833_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i701_3_lut (.I0(n1026), .I1(n1093), 
            .I2(n1059), .I3(GND_net), .O(n1125));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i701_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[11]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15832_3_lut_4_lut (.I0(deadband[11]), .I1(\data_in_frame[15] [3]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29840));   // verilog/coms.v(130[12] 305[6])
    defparam i15832_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15831_3_lut_4_lut (.I0(deadband[12]), .I1(\data_in_frame[15] [4]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29839));   // verilog/coms.v(130[12] 305[6])
    defparam i15831_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5785));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15829_3_lut_4_lut (.I0(deadband[14]), .I1(\data_in_frame[15] [6]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29837));   // verilog/coms.v(130[12] 305[6])
    defparam i15829_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15828_3_lut_4_lut (.I0(deadband[15]), .I1(\data_in_frame[15] [7]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29836));   // verilog/coms.v(130[12] 305[6])
    defparam i15828_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1442_3_lut (.I0(n2119), .I1(n2186), 
            .I2(n2148), .I3(GND_net), .O(n2218));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_4_lut_adj_2198 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(reset), .I3(n42632), .O(n55417));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_4_lut_4_lut_adj_2198.LUT_INIT = 16'hb1f1;
    SB_LUT4 mux_4310_i18_3_lut (.I0(encoder0_position[17]), .I1(n15_adj_5699), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n940));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_245_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[12]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15666_3_lut (.I0(\data_in_frame[22] [3]), .I1(rx_data[3]), 
            .I2(n28428), .I3(GND_net), .O(n29674));   // verilog/coms.v(130[12] 305[6])
    defparam i15666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16375_3_lut (.I0(current[11]), .I1(data_adj_5974[11]), .I2(n27706), 
            .I3(GND_net), .O(n30383));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35007_3_lut_4_lut (.I0(n36723), .I1(Ki[3]), .I2(n4_adj_5802), 
            .I3(n20195), .O(n6_adj_5827));
    defparam i35007_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i1_3_lut_4_lut (.I0(n36723), .I1(Ki[3]), .I2(n4_adj_5802), 
            .I3(n20195), .O(n20149));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i16377_3_lut (.I0(current[10]), .I1(data_adj_5974[10]), .I2(n27706), 
            .I3(GND_net), .O(n30385));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_2199 (.I0(n36723), .I1(Ki[2]), .I2(n48856), 
            .I3(n20196), .O(n20150));
    defparam i1_3_lut_4_lut_adj_2199.LUT_INIT = 16'h8778;
    SB_LUT4 i16378_3_lut (.I0(current[9]), .I1(data_adj_5974[9]), .I2(n27706), 
            .I3(GND_net), .O(n30386));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16379_3_lut (.I0(current[8]), .I1(data_adj_5974[8]), .I2(n27706), 
            .I3(GND_net), .O(n30387));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16380_3_lut (.I0(current[7]), .I1(data_adj_5974[7]), .I2(n27706), 
            .I3(GND_net), .O(n30388));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16380_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16381_3_lut (.I0(current[6]), .I1(data_adj_5974[6]), .I2(n27706), 
            .I3(GND_net), .O(n30389));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16381_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16382_3_lut (.I0(current[5]), .I1(data_adj_5974[5]), .I2(n27706), 
            .I3(GND_net), .O(n30390));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16383_3_lut (.I0(current[4]), .I1(data_adj_5974[4]), .I2(n27706), 
            .I3(GND_net), .O(n30391));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16384_3_lut (.I0(current[3]), .I1(data_adj_5974[3]), .I2(n27706), 
            .I3(GND_net), .O(n30392));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1584_i3_3_lut (.I0(duty[5]), .I1(duty[2]), .I2(n260), 
            .I3(GND_net), .O(n12222));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i16385_3_lut (.I0(current[2]), .I1(data_adj_5974[2]), .I2(n27706), 
            .I3(GND_net), .O(n30393));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16386_3_lut (.I0(current[1]), .I1(data_adj_5974[1]), .I2(n27706), 
            .I3(GND_net), .O(n30394));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16391_3_lut (.I0(baudrate[31]), .I1(data_adj_5966[7]), .I2(n27997), 
            .I3(GND_net), .O(n30399));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16392_3_lut (.I0(baudrate[30]), .I1(data_adj_5966[6]), .I2(n27997), 
            .I3(GND_net), .O(n30400));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16393_3_lut (.I0(baudrate[29]), .I1(data_adj_5966[5]), .I2(n27997), 
            .I3(GND_net), .O(n30401));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16394_3_lut (.I0(baudrate[28]), .I1(data_adj_5966[4]), .I2(n27997), 
            .I3(GND_net), .O(n30402));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5755));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15661_3_lut (.I0(\data_in_frame[22] [2]), .I1(rx_data[2]), 
            .I2(n28428), .I3(GND_net), .O(n29669));   // verilog/coms.v(130[12] 305[6])
    defparam i15661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16395_3_lut (.I0(baudrate[27]), .I1(data_adj_5966[3]), .I2(n27997), 
            .I3(GND_net), .O(n30403));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16396_3_lut (.I0(baudrate[26]), .I1(data_adj_5966[2]), .I2(n27997), 
            .I3(GND_net), .O(n30404));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_245_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[13]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16397_3_lut (.I0(baudrate[25]), .I1(data_adj_5966[1]), .I2(n27997), 
            .I3(GND_net), .O(n30405));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16398_3_lut (.I0(baudrate[24]), .I1(data_adj_5966[0]), .I2(n27997), 
            .I3(GND_net), .O(n30406));   // verilog/eeprom.v(35[8] 81[4])
    defparam i16398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_2200 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[9] [7]), 
            .I2(n57467), .I3(GND_net), .O(n57503));
    defparam i1_2_lut_3_lut_adj_2200.LUT_INIT = 16'h9696;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5756));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34999_3_lut_4_lut (.I0(n36723), .I1(Ki[2]), .I2(n48856), 
            .I3(n20196), .O(n4_adj_5802));
    defparam i34999_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5757));   // verilog/TinyFPGA_B.v(323[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i50641_2_lut (.I0(n69489), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n65487));
    defparam i50641_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_1584_i4_3_lut (.I0(duty[6]), .I1(duty[3]), .I2(n260), 
            .I3(GND_net), .O(n12220));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i15827_3_lut_4_lut (.I0(deadband[16]), .I1(\data_in_frame[14] [0]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29835));   // verilog/coms.v(130[12] 305[6])
    defparam i15827_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15826_3_lut_4_lut (.I0(deadband[17]), .I1(\data_in_frame[14] [1]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29834));   // verilog/coms.v(130[12] 305[6])
    defparam i15826_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 mux_245_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[14]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15825_3_lut_4_lut (.I0(deadband[18]), .I1(\data_in_frame[14] [2]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29833));   // verilog/coms.v(130[12] 305[6])
    defparam i15825_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15824_3_lut_4_lut (.I0(deadband[19]), .I1(\data_in_frame[14] [3]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29832));   // verilog/coms.v(130[12] 305[6])
    defparam i15824_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15823_3_lut_4_lut (.I0(deadband[20]), .I1(\data_in_frame[14] [4]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29831));   // verilog/coms.v(130[12] 305[6])
    defparam i15823_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_4_lut_adj_2201 (.I0(n2021), .I1(n2022), .I2(n61428), .I3(n61426), 
            .O(n61434));
    defparam i1_4_lut_adj_2201.LUT_INIT = 16'hfffe;
    SB_LUT4 i34986_2_lut_3_lut_4_lut (.I0(n36694), .I1(Ki[0]), .I2(Ki[1]), 
            .I3(n36723), .O(n20151));
    defparam i34986_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i15822_3_lut_4_lut (.I0(deadband[21]), .I1(\data_in_frame[14] [5]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29830));   // verilog/coms.v(130[12] 305[6])
    defparam i15822_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i34988_2_lut_3_lut_4_lut (.I0(n36694), .I1(Ki[0]), .I2(Ki[1]), 
            .I3(n36723), .O(n48856));
    defparam i34988_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i15821_3_lut_4_lut (.I0(deadband[22]), .I1(\data_in_frame[14] [6]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29829));   // verilog/coms.v(130[12] 305[6])
    defparam i15821_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15820_3_lut_4_lut (.I0(deadband[23]), .I1(\data_in_frame[14] [7]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29828));   // verilog/coms.v(130[12] 305[6])
    defparam i15820_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i35214_3_lut_4_lut (.I0(n36694), .I1(Ki[3]), .I2(n4_adj_5883), 
            .I3(n20222), .O(n6_adj_5882));
    defparam i35214_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i15819_3_lut_4_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29827));   // verilog/coms.v(130[12] 305[6])
    defparam i15819_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15818_3_lut_4_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29826));   // verilog/coms.v(130[12] 305[6])
    defparam i15818_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_3_lut_4_lut_adj_2202 (.I0(n36694), .I1(Ki[3]), .I2(n4_adj_5883), 
            .I3(n20222), .O(n20194));
    defparam i1_3_lut_4_lut_adj_2202.LUT_INIT = 16'h8778;
    SB_LUT4 mux_245_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[15]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i50305_2_lut (.I0(n69525), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n65441));
    defparam i50305_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_2203 (.I0(n2029), .I1(n43402), .I2(n2030), .I3(n2031), 
            .O(n58718));
    defparam i1_4_lut_adj_2203.LUT_INIT = 16'ha080;
    SB_LUT4 i15817_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29825));   // verilog/coms.v(130[12] 305[6])
    defparam i15817_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i53318_2_lut (.I0(n22849), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_404));
    defparam i53318_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i15816_3_lut_4_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29824));   // verilog/coms.v(130[12] 305[6])
    defparam i15816_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_4_lut_adj_2204 (.I0(n2019), .I1(n58718), .I2(n2020), .I3(n61434), 
            .O(n61440));
    defparam i1_4_lut_adj_2204.LUT_INIT = 16'hfffe;
    SB_LUT4 i15815_3_lut_4_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29823));   // verilog/coms.v(130[12] 305[6])
    defparam i15815_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1105_3_lut (.I0(n1622), .I1(n1689), 
            .I2(n1653), .I3(GND_net), .O(n1721));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15814_3_lut_4_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29822));   // verilog/coms.v(130[12] 305[6])
    defparam i15814_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i53125_4_lut (.I0(n2017), .I1(n2016), .I2(n2018), .I3(n61440), 
            .O(n2049));
    defparam i53125_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15813_3_lut_4_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29821));   // verilog/coms.v(130[12] 305[6])
    defparam i15813_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15812_3_lut_4_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29820));   // verilog/coms.v(130[12] 305[6])
    defparam i15812_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15811_3_lut_4_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29819));   // verilog/coms.v(130[12] 305[6])
    defparam i15811_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15810_3_lut_4_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29818));   // verilog/coms.v(130[12] 305[6])
    defparam i15810_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i22458_3_lut_4_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29817));
    defparam i22458_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16431_3_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(\PID_CONTROLLER.integral_23__N_3715 [23]), 
            .I2(control_update), .I3(GND_net), .O(n30439));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1172_3_lut (.I0(n1721), .I1(n1788_adj_5804), 
            .I2(n1752), .I3(GND_net), .O(n1820));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16432_3_lut (.I0(\PID_CONTROLLER.integral [22]), .I1(\PID_CONTROLLER.integral_23__N_3715 [22]), 
            .I2(control_update), .I3(GND_net), .O(n30440));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16433_3_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral_23__N_3715 [21]), 
            .I2(control_update), .I3(GND_net), .O(n30441));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16434_3_lut (.I0(\PID_CONTROLLER.integral [20]), .I1(\PID_CONTROLLER.integral_23__N_3715 [20]), 
            .I2(control_update), .I3(GND_net), .O(n30442));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22459_3_lut_4_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29816));
    defparam i22459_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i22726_3_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n36694), 
            .I2(control_update), .I3(GND_net), .O(n30443));   // verilog/motorControl.v(20[7:21])
    defparam i22726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1584_i5_3_lut (.I0(duty[7]), .I1(duty[4]), .I2(n260), 
            .I3(GND_net), .O(n12218));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i15807_3_lut_4_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29815));   // verilog/coms.v(130[12] 305[6])
    defparam i15807_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i22756_3_lut (.I0(\PID_CONTROLLER.integral [18]), .I1(n36723), 
            .I2(control_update), .I3(GND_net), .O(n30445));   // verilog/motorControl.v(20[7:21])
    defparam i22756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22793_3_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n36759), 
            .I2(control_update), .I3(GND_net), .O(n30447));   // verilog/motorControl.v(20[7:21])
    defparam i22793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16440_3_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral_23__N_3715 [16]), 
            .I2(control_update), .I3(GND_net), .O(n30448));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15806_3_lut_4_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29814));   // verilog/coms.v(130[12] 305[6])
    defparam i15806_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15866_3_lut (.I0(\data_in_frame[1] [3]), .I1(rx_data[3]), .I2(n57044), 
            .I3(GND_net), .O(n29874));   // verilog/coms.v(130[12] 305[6])
    defparam i15866_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16441_3_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(\PID_CONTROLLER.integral_23__N_3715 [15]), 
            .I2(control_update), .I3(GND_net), .O(n30449));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16442_3_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(\PID_CONTROLLER.integral_23__N_3715 [14]), 
            .I2(control_update), .I3(GND_net), .O(n30450));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16443_3_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(\PID_CONTROLLER.integral_23__N_3715 [13]), 
            .I2(control_update), .I3(GND_net), .O(n30451));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16443_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22435_3_lut (.I0(\PID_CONTROLLER.integral [12]), .I1(\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .I2(control_update), .I3(GND_net), .O(n30452));   // verilog/motorControl.v(20[7:21])
    defparam i22435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16445_3_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .I2(control_update), .I3(GND_net), .O(n30453));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16446_3_lut (.I0(\PID_CONTROLLER.integral [10]), .I1(\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .I2(control_update), .I3(GND_net), .O(n30454));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15805_3_lut_4_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29813));   // verilog/coms.v(130[12] 305[6])
    defparam i15805_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15804_3_lut_4_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29812));   // verilog/coms.v(130[12] 305[6])
    defparam i15804_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i12_4_lut_adj_2205 (.I0(\data_in_frame[22] [7]), .I1(n28375), 
            .I2(n28428), .I3(rx_data[7]), .O(n56027));   // verilog/coms.v(130[12] 305[6])
    defparam i12_4_lut_adj_2205.LUT_INIT = 16'h3a0a;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(current[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5679));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22806_3_lut_4_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29811));
    defparam i22806_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16447_3_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .I2(control_update), .I3(GND_net), .O(n30455));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16448_3_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .I2(control_update), .I3(GND_net), .O(n30456));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22768_3_lut_4_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29810));
    defparam i22768_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(current[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_5678));   // verilog/TinyFPGA_B.v(121[16:24])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22737_3_lut_4_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29809));
    defparam i22737_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16449_3_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .I2(control_update), .I3(GND_net), .O(n30457));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16449_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16450_3_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .I2(control_update), .I3(GND_net), .O(n30458));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15870_3_lut (.I0(\data_in_frame[1] [4]), .I1(rx_data[4]), .I2(n57044), 
            .I3(GND_net), .O(n29878));   // verilog/coms.v(130[12] 305[6])
    defparam i15870_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16451_3_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .I2(control_update), .I3(GND_net), .O(n30459));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16452_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .I2(control_update), .I3(GND_net), .O(n30460));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15873_3_lut (.I0(\data_in_frame[1] [5]), .I1(rx_data[5]), .I2(n57044), 
            .I3(GND_net), .O(n29881));   // verilog/coms.v(130[12] 305[6])
    defparam i15873_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16453_3_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .I2(control_update), .I3(GND_net), .O(n30461));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16453_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15800_3_lut_4_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29808));   // verilog/coms.v(130[12] 305[6])
    defparam i15800_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16454_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .I2(control_update), .I3(GND_net), .O(n30462));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16455_3_lut (.I0(\PID_CONTROLLER.integral [1]), .I1(\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .I2(control_update), .I3(GND_net), .O(n30463));   // verilog/motorControl.v(41[14] 62[8])
    defparam i16455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15799_3_lut_4_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29807));   // verilog/coms.v(130[12] 305[6])
    defparam i15799_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15798_3_lut_4_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29806));   // verilog/coms.v(130[12] 305[6])
    defparam i15798_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1239_3_lut (.I0(n1820), .I1(n1887), 
            .I2(n1851), .I3(GND_net), .O(n1919));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1239_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15797_3_lut_4_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29805));   // verilog/coms.v(130[12] 305[6])
    defparam i15797_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15796_3_lut_4_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29804));   // verilog/coms.v(130[12] 305[6])
    defparam i15796_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15795_3_lut_4_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29803));   // verilog/coms.v(130[12] 305[6])
    defparam i15795_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15794_3_lut_4_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29802));   // verilog/coms.v(130[12] 305[6])
    defparam i15794_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_4_lut_adj_2206 (.I0(control_mode[0]), .I1(n61854), 
            .I2(control_mode[5]), .I3(control_mode[7]), .O(n25398));   // verilog/TinyFPGA_B.v(287[5:22])
    defparam i1_2_lut_4_lut_adj_2206.LUT_INIT = 16'hfffe;
    SB_LUT4 i15793_3_lut_4_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29801));   // verilog/coms.v(130[12] 305[6])
    defparam i15793_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15655_3_lut (.I0(\data_in_frame[22] [1]), .I1(rx_data[1]), 
            .I2(n28428), .I3(GND_net), .O(n29663));   // verilog/coms.v(130[12] 305[6])
    defparam i15655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16480_4_lut (.I0(commutation_state_7__N_27[2]), .I1(commutation_state[1]), 
            .I2(n20890), .I3(n4_adj_5907), .O(n30488));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i16480_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i15792_3_lut_4_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29800));   // verilog/coms.v(130[12] 305[6])
    defparam i15792_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15791_3_lut_4_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29799));   // verilog/coms.v(130[12] 305[6])
    defparam i15791_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16484_4_lut (.I0(state_7__N_4124[3]), .I1(data_adj_5966[0]), 
            .I2(n10_adj_5844), .I3(n25540), .O(n30492));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16484_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16490_3_lut (.I0(n58000), .I1(r_Bit_Index[0]), .I2(n27966), 
            .I3(GND_net), .O(n30498));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16490_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i15789_3_lut_4_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29797));   // verilog/coms.v(130[12] 305[6])
    defparam i15789_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i4891_4_lut (.I0(n25422), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5816));
    defparam i4891_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut (.I0(n24_adj_5816), .I1(delay_counter[14]), .I2(delay_counter[12]), 
            .I3(delay_counter[13]), .O(n59675));
    defparam i2_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 i2_3_lut_adj_2207 (.I0(n59675), .I1(delay_counter[18]), .I2(n25424), 
            .I3(GND_net), .O(n59710));
    defparam i2_3_lut_adj_2207.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_1584_i6_3_lut (.I0(duty[8]), .I1(duty[5]), .I2(n260), 
            .I3(GND_net), .O(n12216));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i15788_3_lut_4_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29796));   // verilog/coms.v(130[12] 305[6])
    defparam i15788_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i2_4_lut_adj_2208 (.I0(n59710), .I1(delay_counter[23]), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7_adj_5898));
    defparam i2_4_lut_adj_2208.LUT_INIT = 16'heccc;
    SB_LUT4 i4_4_lut_adj_2209 (.I0(n7_adj_5898), .I1(delay_counter[21]), 
            .I2(delay_counter[22]), .I3(n25410), .O(n62));
    defparam i4_4_lut_adj_2209.LUT_INIT = 16'hfffe;
    SB_LUT4 i16494_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n60772), 
            .I3(n27_adj_5781), .O(n30502));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i16494_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15787_3_lut_4_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29795));   // verilog/coms.v(130[12] 305[6])
    defparam i15787_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i16498_4_lut (.I0(CS_MISO_c), .I1(data_adj_5974[0]), .I2(n11_adj_5734), 
            .I3(state_7__N_4317), .O(n30506));   // verilog/tli4970.v(35[10] 68[6])
    defparam i16498_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i28913_2_lut (.I0(n62), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_409));   // verilog/TinyFPGA_B.v(365[12:35])
    defparam i28913_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5_3_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n14_adj_5909));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_2210 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15_adj_5908));
    defparam i6_4_lut_adj_2210.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_2211 (.I0(n15_adj_5908), .I1(delay_counter[2]), 
            .I2(n14_adj_5909), .I3(delay_counter[6]), .O(n25422));
    defparam i8_4_lut_adj_2211.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_2212 (.I0(delay_counter[27]), .I1(delay_counter[29]), 
            .I2(delay_counter[24]), .I3(delay_counter[26]), .O(n12_adj_5890));
    defparam i5_4_lut_adj_2212.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_2213 (.I0(delay_counter[28]), .I1(n12_adj_5890), 
            .I2(delay_counter[25]), .I3(delay_counter[30]), .O(n25410));
    defparam i6_4_lut_adj_2213.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_2214 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n25424));
    defparam i2_3_lut_adj_2214.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_2215 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5893));
    defparam i1_2_lut_adj_2215.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_30__I_0_i1306_3_lut (.I0(n1919), .I1(n1986), 
            .I2(n1950), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1306_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_4_lut_adj_2216 (.I0(delay_counter[9]), .I1(n4_adj_5893), 
            .I2(delay_counter[10]), .I3(n25422), .O(n59575));
    defparam i2_4_lut_adj_2216.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_2217 (.I0(n59575), .I1(n25424), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n59282));
    defparam i2_4_lut_adj_2217.LUT_INIT = 16'hffec;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_5914));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut_adj_2218 (.I0(delay_counter[22]), .I1(n59282), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5915));
    defparam i2_4_lut_adj_2218.LUT_INIT = 16'ha8a0;
    SB_LUT4 i28918_4_lut (.I0(n7_adj_5915), .I1(delay_counter[31]), .I2(n25410), 
            .I3(n8_adj_5914), .O(n1319));   // verilog/TinyFPGA_B.v(379[14:38])
    defparam i28918_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i15786_3_lut_4_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29794));   // verilog/coms.v(130[12] 305[6])
    defparam i15786_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i30_4_lut (.I0(state_7__N_3916[0]), .I1(n25404), .I2(state_adj_5967[1]), 
            .I3(n4_adj_5842), .O(n12_adj_5912));   // verilog/eeprom.v(35[8] 81[4])
    defparam i30_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i29_4_lut (.I0(n12_adj_5912), .I1(n65486), .I2(state_adj_5967[0]), 
            .I3(state_adj_5967[2]), .O(n56203));   // verilog/eeprom.v(35[8] 81[4])
    defparam i29_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 i15785_3_lut_4_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29793));   // verilog/coms.v(130[12] 305[6])
    defparam i15785_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i584_2_lut (.I0(n1319), .I1(n42632), .I2(GND_net), .I3(GND_net), 
            .O(n2820));   // verilog/TinyFPGA_B.v(383[18] 385[12])
    defparam i584_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_245_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15_adj_5681), .I3(n15), .O(motor_state_23__N_91[17]));   // verilog/TinyFPGA_B.v(286[5] 288[10])
    defparam mux_245_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i49959_4_lut (.I0(data_ready), .I1(n6617), .I2(n24_adj_5895), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n65444));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i49959_4_lut.LUT_INIT = 16'hdccc;
    SB_LUT4 i50587_2_lut (.I0(n24_adj_5895), .I1(n6617), .I2(GND_net), 
            .I3(GND_net), .O(n65447));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i50587_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49_4_lut (.I0(n65447), .I1(n65444), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(n6_adj_5900), .O(n55331));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i49_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i15961_3_lut_4_lut (.I0(reset), .I1(n172), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n29969));
    defparam i15961_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15938_3_lut_4_lut (.I0(reset), .I1(n172), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n29946));
    defparam i15938_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1584_i7_3_lut (.I0(duty[9]), .I1(duty[6]), .I2(n260), 
            .I3(GND_net), .O(n12214));   // verilog/TinyFPGA_B.v(117[13] 128[7])
    defparam mux_1584_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i15784_3_lut_4_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29792));   // verilog/coms.v(130[12] 305[6])
    defparam i15784_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15941_3_lut_4_lut (.I0(reset), .I1(n172), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n29949));
    defparam i15941_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15945_3_lut_4_lut (.I0(reset), .I1(n172), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n29953));
    defparam i15945_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 encoder0_position_30__I_0_i1318_3_lut (.I0(n1931), .I1(n1998), 
            .I2(n1950), .I3(GND_net), .O(n2030));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i42186_3_lut (.I0(n5_adj_5709), .I1(n7453), .I2(n57811), .I3(GND_net), 
            .O(n57816));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1386_3_lut (.I0(n2031), .I1(n2098), 
            .I2(n2049), .I3(GND_net), .O(n2130));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i42187_3_lut (.I0(encoder0_position[27]), .I1(n57816), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1385_3_lut (.I0(n2030), .I1(n2097), 
            .I2(n2049), .I3(GND_net), .O(n2129));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i570_3_lut (.I0(n831), .I1(n898), 
            .I2(n861), .I3(GND_net), .O(n930));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15948_3_lut_4_lut (.I0(reset), .I1(n172), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n29956));
    defparam i15948_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15951_3_lut_4_lut (.I0(reset), .I1(n172), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n29959));
    defparam i15951_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15783_3_lut_4_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29791));   // verilog/coms.v(130[12] 305[6])
    defparam i15783_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1389_3_lut (.I0(n945), .I1(n2101), 
            .I2(n2049), .I3(GND_net), .O(n2133));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i637_3_lut (.I0(n930), .I1(n997), 
            .I2(n960), .I3(GND_net), .O(n1029));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i1388_3_lut (.I0(n2033), .I1(n2100), 
            .I2(n2049), .I3(GND_net), .O(n2132));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i704_3_lut (.I0(n1029), .I1(n1096), 
            .I2(n1059), .I3(GND_net), .O(n1128));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1387_3_lut (.I0(n2032), .I1(n2099), 
            .I2(n2049), .I3(GND_net), .O(n2131));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i771_3_lut (.I0(n1128), .I1(n1195), 
            .I2(n1158), .I3(GND_net), .O(n1227_adj_5795));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i771_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i12_3_lut (.I0(encoder0_position[11]), .I1(n21_adj_5693), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n946));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_2219 (.I0(ID[5]), .I1(ID[4]), .I2(ID[1]), .I3(ID[7]), 
            .O(n14_adj_5686));   // verilog/TinyFPGA_B.v(377[12:17])
    defparam i6_4_lut_adj_2219.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_30__I_0_i838_3_lut (.I0(n1227_adj_5795), .I1(n1294), 
            .I2(n1257), .I3(GND_net), .O(n1326));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1379_3_lut (.I0(n2024), .I1(n2091), 
            .I2(n2049), .I3(GND_net), .O(n2123));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5_4_lut_adj_2220 (.I0(ID[0]), .I1(ID[3]), .I2(ID[6]), .I3(ID[2]), 
            .O(n13_adj_5687));   // verilog/TinyFPGA_B.v(377[12:17])
    defparam i5_4_lut_adj_2220.LUT_INIT = 16'hfffe;
    SB_LUT4 i28730_4_lut (.I0(n13_adj_5687), .I1(baudrate[0]), .I2(n14_adj_5686), 
            .I3(n25530), .O(n42632));
    defparam i28730_4_lut.LUT_INIT = 16'hc8fa;
    SB_LUT4 encoder0_position_30__I_0_i905_3_lut (.I0(n1326), .I1(n1393), 
            .I2(n1356), .I3(GND_net), .O(n1425));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i905_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1378_3_lut (.I0(n2023), .I1(n2090), 
            .I2(n2049), .I3(GND_net), .O(n2122));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i972_3_lut (.I0(n1425), .I1(n1492), 
            .I2(n1455), .I3(GND_net), .O(n1524));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i972_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1039_3_lut (.I0(n1524), .I1(n1591), 
            .I2(n1554), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1377_3_lut (.I0(n2022), .I1(n2089), 
            .I2(n2049), .I3(GND_net), .O(n2121));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14877_4_lut (.I0(n27698), .I1(n1319), .I2(n65309), .I3(n42746), 
            .O(n28885));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i14877_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53603 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n69306));
    defparam byte_transmit_counter_0__bdd_4_lut_53603.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_30__I_0_i1106_3_lut (.I0(n1623), .I1(n1690), 
            .I2(n1653), .I3(GND_net), .O(n1722));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1173_3_lut (.I0(n1722), .I1(n1789), 
            .I2(n1752), .I3(GND_net), .O(n1821));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15782_3_lut_4_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29790));   // verilog/coms.v(130[12] 305[6])
    defparam i15782_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_adj_2221 (.I0(n2128), .I1(n2124), .I2(GND_net), .I3(GND_net), 
            .O(n61086));
    defparam i1_2_lut_adj_2221.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_30__I_0_i1441_3_lut (.I0(n2118), .I1(n2185), 
            .I2(n2148), .I3(GND_net), .O(n2217));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1240_3_lut (.I0(n1821), .I1(n1888), 
            .I2(n1851), .I3(GND_net), .O(n1920));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_2222 (.I0(n2126), .I1(n61086), .I2(n2127), .I3(n2125), 
            .O(n61090));
    defparam i1_4_lut_adj_2222.LUT_INIT = 16'hfffe;
    SB_LUT4 i42188_3_lut (.I0(n6_adj_5707), .I1(n7454), .I2(n57811), .I3(GND_net), 
            .O(n57818));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29679_4_lut (.I0(n946), .I1(n2131), .I2(n2132), .I3(n2133), 
            .O(n43588));
    defparam i29679_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i42189_3_lut (.I0(encoder0_position[26]), .I1(n57818), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n69306_bdd_4_lut (.I0(n69306), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n69309));
    defparam n69306_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15781_3_lut_4_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29789));   // verilog/coms.v(130[12] 305[6])
    defparam i15781_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15780_3_lut_4_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29788));   // verilog/coms.v(130[12] 305[6])
    defparam i15780_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_4_lut_adj_2223 (.I0(n2121), .I1(n2122), .I2(n61090), .I3(n2123), 
            .O(n61096));
    defparam i1_4_lut_adj_2223.LUT_INIT = 16'hfffe;
    SB_LUT4 i15779_3_lut_4_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29787));   // verilog/coms.v(130[12] 305[6])
    defparam i15779_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i571_3_lut (.I0(n832), .I1(n899), 
            .I2(n861), .I3(GND_net), .O(n931));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i638_3_lut (.I0(n931), .I1(n998), 
            .I2(n960), .I3(GND_net), .O(n1030));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15778_3_lut_4_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29786));   // verilog/coms.v(130[12] 305[6])
    defparam i15778_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15777_3_lut_4_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29785));   // verilog/coms.v(130[12] 305[6])
    defparam i15777_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i637_1_lut (.I0(reset), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2873));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i637_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i705_3_lut (.I0(n1030), .I1(n1097), 
            .I2(n1059), .I3(GND_net), .O(n1129));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i772_3_lut (.I0(n1129), .I1(n1196), 
            .I2(n1158), .I3(GND_net), .O(n1228_adj_5796));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2224 (.I0(n36759), .I1(Ki[1]), .I2(GND_net), 
            .I3(GND_net), .O(n125));
    defparam i1_2_lut_adj_2224.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_2225 (.I0(n36723), .I1(Ki[0]), .I2(GND_net), 
            .I3(GND_net), .O(n56));
    defparam i1_2_lut_adj_2225.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_i839_3_lut (.I0(n1228_adj_5796), .I1(n1295), 
            .I2(n1257), .I3(GND_net), .O(n1327));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16732_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [2]), 
            .O(n30740));   // verilog/coms.v(130[12] 305[6])
    defparam i16732_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_2226 (.I0(n2129), .I1(n61096), .I2(n43588), .I3(n2130), 
            .O(n61098));
    defparam i1_4_lut_adj_2226.LUT_INIT = 16'heccc;
    SB_LUT4 i15776_3_lut_4_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29784));   // verilog/coms.v(130[12] 305[6])
    defparam i15776_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_4_lut_adj_2227 (.I0(n2118), .I1(n2119), .I2(n2120), .I3(n61098), 
            .O(n61104));
    defparam i1_4_lut_adj_2227.LUT_INIT = 16'hfffe;
    SB_LUT4 i53149_4_lut (.I0(n2116), .I1(n2115), .I2(n2117), .I3(n61104), 
            .O(n2148));
    defparam i53149_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_30__I_0_i906_3_lut (.I0(n1327), .I1(n1394), 
            .I2(n1356), .I3(GND_net), .O(n1426));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i906_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15775_3_lut_4_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29783));   // verilog/coms.v(130[12] 305[6])
    defparam i15775_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i973_3_lut (.I0(n1426), .I1(n1493), 
            .I2(n1455), .I3(GND_net), .O(n1525));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i973_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1040_3_lut (.I0(n1525), .I1(n1592), 
            .I2(n1554), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15774_3_lut_4_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29782));   // verilog/coms.v(130[12] 305[6])
    defparam i15774_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15773_3_lut_4_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29781));   // verilog/coms.v(130[12] 305[6])
    defparam i15773_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15772_3_lut_4_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29780));   // verilog/coms.v(130[12] 305[6])
    defparam i15772_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i2_2_lut_adj_2228 (.I0(hall2), .I1(commutation_state_7__N_27[2]), 
            .I2(GND_net), .I3(GND_net), .O(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(166[7:32])
    defparam i2_2_lut_adj_2228.LUT_INIT = 16'h4444;
    SB_LUT4 i16577_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [0]), 
            .O(n30585));   // verilog/coms.v(130[12] 305[6])
    defparam i16577_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i42311_3_lut_4_lut (.I0(n8_adj_5760), .I1(n57917), .I2(n10_adj_5758), 
            .I3(reset), .O(n57948));
    defparam i42311_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i15771_3_lut_4_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29779));   // verilog/coms.v(130[12] 305[6])
    defparam i15771_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_3_lut_adj_2229 (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_208[0]));   // verilog/TinyFPGA_B.v(163[4] 165[7])
    defparam i1_3_lut_adj_2229.LUT_INIT = 16'h1414;
    SB_LUT4 i1_2_lut_3_lut_adj_2230 (.I0(hall1), .I1(hall2), .I2(n20890), 
            .I3(GND_net), .O(n4_adj_5907));   // verilog/TinyFPGA_B.v(151[7:22])
    defparam i1_2_lut_3_lut_adj_2230.LUT_INIT = 16'hf2f2;
    SB_LUT4 i53474_4_lut_4_lut_4_lut (.I0(hall3), .I1(hall1), .I2(commutation_state_7__N_27[2]), 
            .I3(hall2), .O(n7_adj_5916));
    defparam i53474_4_lut_4_lut_4_lut.LUT_INIT = 16'h77fc;
    SB_LUT4 i15770_3_lut_4_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29778));   // verilog/coms.v(130[12] 305[6])
    defparam i15770_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15769_3_lut_4_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29777));   // verilog/coms.v(130[12] 305[6])
    defparam i15769_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15767_3_lut_4_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29775));   // verilog/coms.v(130[12] 305[6])
    defparam i15767_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_4_lut_4_lut_adj_2231 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(read_N_409), .I3(n2820), .O(n25_adj_5897));   // verilog/TinyFPGA_B.v(376[7:11])
    defparam i1_4_lut_4_lut_adj_2231.LUT_INIT = 16'h5450;
    SB_LUT4 encoder0_position_30__I_0_i1107_3_lut (.I0(n1624), .I1(n1691), 
            .I2(n1653), .I3(GND_net), .O(n1723));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14864_2_lut (.I0(n27646), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n28878));   // verilog/TinyFPGA_B.v(143[9] 222[5])
    defparam i14864_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52635_4_lut (.I0(commutation_state[1]), .I1(n22849), .I2(dti), 
            .I3(commutation_state[2]), .O(n27646));
    defparam i52635_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 encoder0_position_30__I_0_i1373_3_lut (.I0(n2018), .I1(n2085), 
            .I2(n2049), .I3(GND_net), .O(n2117));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1174_3_lut (.I0(n1723), .I1(n1790_adj_5805), 
            .I2(n1752), .I3(GND_net), .O(n1822_adj_5809));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1440_3_lut (.I0(n2117), .I1(n2184), 
            .I2(n2148), .I3(GND_net), .O(n2216));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1241_3_lut (.I0(n1822_adj_5809), .I1(n1889), 
            .I2(n1851), .I3(GND_net), .O(n1921));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1241_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1308_3_lut (.I0(n1921), .I1(n1988), 
            .I2(n1950), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i26_3_lut (.I0(encoder0_position[25]), .I1(n7_adj_5706), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n518));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_2232 (.I0(n4_adj_5714), .I1(n5_adj_5709), .I2(n518), 
            .I3(n6_adj_5707), .O(n5_adj_5894));
    defparam i1_4_lut_adj_2232.LUT_INIT = 16'heeea;
    SB_LUT4 i1_3_lut_adj_2233 (.I0(n3), .I1(n2_adj_5715), .I2(n5_adj_5894), 
            .I3(GND_net), .O(n57811));
    defparam i1_3_lut_adj_2233.LUT_INIT = 16'h8080;
    SB_LUT4 i15738_3_lut_3_lut (.I0(\FRAME_MATCHER.rx_data_ready_prev ), .I1(rx_data_ready), 
            .I2(reset), .I3(GND_net), .O(n29746));   // verilog/coms.v(130[12] 305[6])
    defparam i15738_3_lut_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_3_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2513 ), 
            .I2(n33769), .I3(GND_net), .O(n22726));   // verilog/TinyFPGA_B.v(358[10] 388[6])
    defparam i1_3_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i42190_3_lut (.I0(n7_adj_5706), .I1(n7455), .I2(n57811), .I3(GND_net), 
            .O(n57820));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42191_3_lut (.I0(encoder0_position[25]), .I1(n57820), .I2(encoder0_position[30]), 
            .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam i42191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_2234 (.I0(commutation_state[0]), .I1(n4_adj_5684), 
            .I2(commutation_state_prev[0]), .I3(dti_N_404), .O(n27622));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_2_lut_4_lut_adj_2234.LUT_INIT = 16'hdeff;
    SB_LUT4 encoder0_position_30__I_0_i572_3_lut (.I0(n833), .I1(n900), 
            .I2(n861), .I3(GND_net), .O(n932));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i639_3_lut (.I0(n932), .I1(n999), 
            .I2(n960), .I3(GND_net), .O(n1031));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_2235 (.I0(commutation_state[0]), .I1(n4_adj_5684), 
            .I2(commutation_state_prev[0]), .I3(n42723), .O(n27780));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i1_2_lut_4_lut_adj_2235.LUT_INIT = 16'hffde;
    SB_LUT4 i15159_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5684), 
            .I2(commutation_state_prev[0]), .I3(n42723), .O(n29162));   // verilog/TinyFPGA_B.v(146[7:48])
    defparam i15159_2_lut_4_lut.LUT_INIT = 16'h00de;
    SB_LUT4 encoder0_position_30__I_0_i706_3_lut (.I0(n1031), .I1(n1098), 
            .I2(n1059), .I3(GND_net), .O(n1130));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i706_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i50284_2_lut (.I0(n111_adj_5814), .I1(n8_adj_5786), .I2(GND_net), 
            .I3(GND_net), .O(n65437));   // verilog/coms.v(94[13:20])
    defparam i50284_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_30__I_0_i773_3_lut (.I0(n1130), .I1(n1197), 
            .I2(n1158), .I3(GND_net), .O(n1229_adj_5797));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_1083_i6_3_lut_3_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), .O(n6_adj_5829));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1083_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i50495_3_lut_4_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count[2]), .O(n66181));   // verilog/uart_rx.v(119[17:57])
    defparam i50495_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i27070_4_lut (.I0(n65437), .I1(n65436), .I2(rx_data[0]), .I3(\data_in_frame[22] [0]), 
            .O(n41003));   // verilog/coms.v(94[13:20])
    defparam i27070_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 encoder0_position_30__I_0_i840_3_lut (.I0(n1229_adj_5797), .I1(n1296), 
            .I2(n1257), .I3(GND_net), .O(n1328));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i27071_3_lut (.I0(n41003), .I1(\data_in_frame[22] [0]), .I2(reset), 
            .I3(GND_net), .O(n29968));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i27071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_30__I_0_i907_3_lut (.I0(n1328), .I1(n1395), 
            .I2(n1356), .I3(GND_net), .O(n1427));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i974_3_lut (.I0(n1427), .I1(n1494), 
            .I2(n1455), .I3(GND_net), .O(n1526));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_15_inv_0_i24_1_lut (.I0(duty[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(119[24:29])
    defparam unary_minus_15_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1041_3_lut (.I0(n1526), .I1(n1593), 
            .I2(n1554), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1108_3_lut (.I0(n1625), .I1(n1692), 
            .I2(n1653), .I3(GND_net), .O(n1724));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15716_3_lut_4_lut (.I0(n1742), .I1(b_prev), .I2(a_new[1]), 
            .I3(position_31__N_3827), .O(n29724));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15716_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 encoder0_position_30__I_0_i1175_3_lut (.I0(n1724), .I1(n1791), 
            .I2(n1752), .I3(GND_net), .O(n1823));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1242_3_lut (.I0(n1823), .I1(n1890), 
            .I2(n1851), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1242_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1309_3_lut (.I0(n1922), .I1(n1989), 
            .I2(n1950), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1307_3_lut (.I0(n1920), .I1(n1987), 
            .I2(n1950), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1376_3_lut (.I0(n2021), .I1(n2088), 
            .I2(n2049), .I3(GND_net), .O(n2120));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1375_3_lut (.I0(n2020), .I1(n2087), 
            .I2(n2049), .I3(GND_net), .O(n2119));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_2236 (.I0(n36759), .I1(Ki[2]), .I2(GND_net), 
            .I3(GND_net), .O(n198));
    defparam i1_2_lut_adj_2236.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_i1374_3_lut (.I0(n2019), .I1(n2086), 
            .I2(n2049), .I3(GND_net), .O(n2118));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_4310_i25_3_lut (.I0(encoder0_position[24]), .I1(n8_adj_5705), 
            .I2(encoder0_position[30]), .I3(GND_net), .O(n519));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam mux_4310_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15592_3_lut_4_lut (.I0(reset), .I1(n28383), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n29600));
    defparam i15592_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21755_3_lut_4_lut (.I0(reset), .I1(n28383), .I2(\data_in_frame[20] [6]), 
            .I3(rx_data[6]), .O(n30155));
    defparam i21755_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i15586_3_lut_4_lut (.I0(reset), .I1(n28383), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n29594));
    defparam i15586_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15583_3_lut_4_lut (.I0(reset), .I1(n28383), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n29591));
    defparam i15583_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 encoder0_position_30__I_0_i573_3_lut (.I0(n519), .I1(n901), 
            .I2(n861), .I3(GND_net), .O(n933));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15580_3_lut_4_lut (.I0(reset), .I1(n28383), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n29588));
    defparam i15580_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15571_3_lut_4_lut (.I0(reset), .I1(n28383), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n29579));
    defparam i15571_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 encoder0_position_30__I_0_i640_3_lut (.I0(n933), .I1(n1000), 
            .I2(n960), .I3(GND_net), .O(n1032));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28821_2_lut (.I0(n22849), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n42723));
    defparam i28821_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_30__I_0_i707_3_lut (.I0(n1032), .I1(n1099), 
            .I2(n1059), .I3(GND_net), .O(n1131));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i774_3_lut (.I0(n1131), .I1(n1198), 
            .I2(n1158), .I3(GND_net), .O(n1230_adj_5798));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i841_3_lut (.I0(n1230_adj_5798), .I1(n1297), 
            .I2(n1257), .I3(GND_net), .O(n1329));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i908_3_lut (.I0(n1329), .I1(n1396), 
            .I2(n1356), .I3(GND_net), .O(n1428));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i975_3_lut (.I0(n1428), .I1(n1495), 
            .I2(n1455), .I3(GND_net), .O(n1527));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_30__I_0_i1042_3_lut (.I0(n1527), .I1(n1594), 
            .I2(n1554), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15696_3_lut_4_lut (.I0(n1784), .I1(b_prev_adj_5736), .I2(a_new_adj_5954[1]), 
            .I3(position_31__N_3827_adj_5737), .O(n29704));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15696_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 encoder0_position_30__I_0_i1109_3_lut (.I0(n1626), .I1(n1693), 
            .I2(n1653), .I3(GND_net), .O(n1725));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15653_4_lut_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5986[1]), 
            .I2(r_SM_Main_adj_5986[2]), .I3(n6_adj_5891), .O(n29661));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i15653_4_lut_4_lut.LUT_INIT = 16'ha3aa;
    SB_LUT4 i15636_3_lut_4_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29644));   // verilog/coms.v(130[12] 305[6])
    defparam i15636_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_3_lut_4_lut_adj_2237 (.I0(n51676), .I1(\data_out_frame[19] [7]), 
            .I2(\data_out_frame[19] [6]), .I3(n57131), .O(n6_adj_5824));
    defparam i1_3_lut_4_lut_adj_2237.LUT_INIT = 16'h9669;
    SB_LUT4 encoder0_position_30__I_0_i1176_3_lut (.I0(n1725), .I1(n1792_adj_5806), 
            .I2(n1752), .I3(GND_net), .O(n1824_adj_5810));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i50485_3_lut_4_lut (.I0(r_Clock_Count_adj_5987[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count_adj_5987[2]), .O(n66171));   // verilog/uart_tx.v(117[17:57])
    defparam i50485_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_1086_i6_3_lut_3_lut (.I0(r_Clock_Count_adj_5987[3]), 
            .I1(o_Rx_DV_N_3488[3]), .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), 
            .O(n6_adj_5833));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1086_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    motorControl control (.GND_net(GND_net), .control_update(control_update), 
            .duty({duty}), .clk16MHz(clk16MHz), .reset(reset), .\PID_CONTROLLER.integral ({\PID_CONTROLLER.integral }), 
            .PWMLimit({PWMLimit}), .n361(n361), .IntegralLimit({IntegralLimit}), 
            .n155(n155), .\PID_CONTROLLER.integral_23__N_3715[0] (\PID_CONTROLLER.integral_23__N_3715 [0]), 
            .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), .\Kp[1] (Kp[1]), 
            .\Kp[10] (Kp[10]), .\Kp[0] (Kp[0]), .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), 
            .n20194(n20194), .n6(n6_adj_5827), .n36723(n36723), .\Ki[4] (Ki[4]), 
            .\Kp[4] (Kp[4]), .\Ki[0] (Ki[0]), .\Kp[5] (Kp[5]), .\Ki[2] (Ki[2]), 
            .\PID_CONTROLLER.integral_23__N_3715[20] (\PID_CONTROLLER.integral_23__N_3715 [20]), 
            .n20222(n20222), .\Kp[11] (Kp[11]), .n212(n212), .n213(n213), 
            .\PID_CONTROLLER.integral_23__N_3715[22] (\PID_CONTROLLER.integral_23__N_3715 [22]), 
            .\PID_CONTROLLER.integral_23__N_3715[21] (\PID_CONTROLLER.integral_23__N_3715 [21]), 
            .\Ki[1] (Ki[1]), .\PID_CONTROLLER.integral_23__N_3715[23] (\PID_CONTROLLER.integral_23__N_3715 [23]), 
            .n36694(n36694), .\Ki[5] (Ki[5]), .\Kp[12] (Kp[12]), .\Ki[3] (Ki[3]), 
            .\Kp[13] (Kp[13]), .n6_adj_31(n6_adj_5882), .\Kp[6] (Kp[6]), 
            .\Kp[14] (Kp[14]), .\Kp[15] (Kp[15]), .deadband({deadband}), 
            .\PID_CONTROLLER.integral_23__N_3715[13] (\PID_CONTROLLER.integral_23__N_3715 [13]), 
            .\PID_CONTROLLER.integral_23__N_3715[12] (\PID_CONTROLLER.integral_23__N_3715 [12]), 
            .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), .\Ki[9] (Ki[9]), 
            .\Ki[10] (Ki[10]), .\Ki[11] (Ki[11]), .n219(n219), .\PID_CONTROLLER.integral_23__N_3715[11] (\PID_CONTROLLER.integral_23__N_3715 [11]), 
            .\Ki[12] (Ki[12]), .n53(n53), .\PID_CONTROLLER.integral_23__N_3715[10] (\PID_CONTROLLER.integral_23__N_3715 [10]), 
            .\Ki[13] (Ki[13]), .n4(n4_adj_5821), .\PID_CONTROLLER.integral_23__N_3715[9] (\PID_CONTROLLER.integral_23__N_3715 [9]), 
            .n11610(n11610), .n27692(n27692), .\Ki[14] (Ki[14]), .\PID_CONTROLLER.integral_23__N_3715[8] (\PID_CONTROLLER.integral_23__N_3715 [8]), 
            .setpoint({setpoint}), .\motor_state[23] (motor_state[23]), 
            .\motor_state[22] (motor_state[22]), .\motor_state[21] (motor_state[21]), 
            .\Ki[15] (Ki[15]), .\PID_CONTROLLER.integral_23__N_3715[7] (\PID_CONTROLLER.integral_23__N_3715 [7]), 
            .n38(n38), .n110(n110), .\PID_CONTROLLER.integral_23__N_3715[14] (\PID_CONTROLLER.integral_23__N_3715 [14]), 
            .\motor_state[20] (motor_state[20]), .\motor_state[19] (motor_state[19]), 
            .n490(n490), .n417(n417), .n20149(n20149), .n344(n344), 
            .n20150(n20150), .n271(n271), .\PID_CONTROLLER.integral_23__N_3715[6] (\PID_CONTROLLER.integral_23__N_3715 [6]), 
            .n29641(n29641), .n20151(n20151), .n198(n198), .VCC_net(VCC_net), 
            .n56(n56), .n125(n125), .n30463(n30463), .n30462(n30462), 
            .n30461(n30461), .n30460(n30460), .n30459(n30459), .n30458(n30458), 
            .n30457(n30457), .n30456(n30456), .n30455(n30455), .n30454(n30454), 
            .n30453(n30453), .n30452(n30452), .n30451(n30451), .n30450(n30450), 
            .n30449(n30449), .n30448(n30448), .n30447(n30447), .n30445(n30445), 
            .n30443(n30443), .n30442(n30442), .n30441(n30441), .n30440(n30440), 
            .n30439(n30439), .\motor_state[18] (motor_state[18]), .\PID_CONTROLLER.integral_23__N_3715[5] (\PID_CONTROLLER.integral_23__N_3715 [5]), 
            .n455(n455), .n456(n456), .\motor_state[17] (motor_state[17]), 
            .n20(n20_adj_5812), .\motor_state[15] (motor_state[15]), .\motor_state[14] (motor_state[14]), 
            .\motor_state[13] (motor_state[13]), .\motor_state[12] (motor_state[12]), 
            .n1(n1), .\motor_state[10] (motor_state[10]), .\motor_state[9] (motor_state[9]), 
            .\motor_state[8] (motor_state[8]), .n401(n401), .n43(n43_adj_5825), 
            .\motor_state[7] (motor_state[7]), .n41622(n41622), .\motor_state[5] (motor_state[5]), 
            .\motor_state[4] (motor_state[4]), .n42235(n42235), .\motor_state[2] (motor_state[2]), 
            .\motor_state[1] (motor_state[1]), .\motor_state[0] (motor_state[0]), 
            .n375(n375), .n376(n376), .\PID_CONTROLLER.integral_23__N_3715[4] (\PID_CONTROLLER.integral_23__N_3715 [4]), 
            .\PID_CONTROLLER.integral_23__N_3715[3] (\PID_CONTROLLER.integral_23__N_3715 [3]), 
            .\PID_CONTROLLER.integral_23__N_3715[15] (\PID_CONTROLLER.integral_23__N_3715 [15]), 
            .\PID_CONTROLLER.integral_23__N_3715[16] (\PID_CONTROLLER.integral_23__N_3715 [16]), 
            .\PID_CONTROLLER.integral_23__N_3715[2] (\PID_CONTROLLER.integral_23__N_3715 [2]), 
            .\PID_CONTROLLER.integral_23__N_3715[1] (\PID_CONTROLLER.integral_23__N_3715 [1]), 
            .n214(n214), .n131(n131), .n204(n204), .n4_adj_32(n4_adj_5883), 
            .n20195(n20195), .n43349(n43349), .n37189(n37189), .n4_adj_33(n4_adj_5818), 
            .n30(n30_adj_5819), .n32(n32_adj_5820), .n4_adj_34(n4_adj_5817), 
            .n20196(n20196)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(290[16] 302[4])
    SB_LUT4 encoder0_position_30__I_0_i1243_3_lut (.I0(n1824_adj_5810), .I1(n1891), 
            .I2(n1851), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1243_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15628_3_lut_4_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29636));   // verilog/coms.v(130[12] 305[6])
    defparam i15628_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i15627_3_lut_4_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29635));   // verilog/coms.v(130[12] 305[6])
    defparam i15627_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 encoder0_position_30__I_0_i1310_3_lut (.I0(n1923), .I1(n1990), 
            .I2(n1950), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15605_3_lut_4_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29613));   // verilog/coms.v(130[12] 305[6])
    defparam i15605_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    \quadrature_decoder(1)  quad_counter1 (.b_prev(b_prev_adj_5736), .GND_net(GND_net), 
            .a_new({a_new_adj_5954[1], Open_4}), .position_31__N_3827(position_31__N_3827_adj_5737), 
            .ENCODER1_B_N_keep(ENCODER1_B_N), .n1779(clk16MHz), .ENCODER1_A_N_keep(ENCODER1_A_N), 
            .n29704(n29704), .n1784(n1784), .n1824(n1824), .n1786(n1786), 
            .n1788(n1788), .n1790(n1790), .n1792(n1792), .n1794(n1794), 
            .n1796(n1796), .\encoder1_position[25] (encoder1_position[25]), 
            .\encoder1_position[24] (encoder1_position[24]), .\encoder1_position[23] (encoder1_position[23]), 
            .\encoder1_position[22] (encoder1_position[22]), .\encoder1_position[21] (encoder1_position[21]), 
            .\encoder1_position[20] (encoder1_position[20]), .\encoder1_position[19] (encoder1_position[19]), 
            .\encoder1_position[18] (encoder1_position[18]), .\encoder1_position[17] (encoder1_position[17]), 
            .\encoder1_position[16] (encoder1_position[16]), .\encoder1_position[15] (encoder1_position[15]), 
            .\encoder1_position[14] (encoder1_position[14]), .\encoder1_position[13] (encoder1_position[13]), 
            .\encoder1_position[12] (encoder1_position[12]), .\encoder1_position[11] (encoder1_position[11]), 
            .\encoder1_position[10] (encoder1_position[10]), .\encoder1_position[9] (encoder1_position[9]), 
            .\encoder1_position[8] (encoder1_position[8]), .\encoder1_position[7] (encoder1_position[7]), 
            .\encoder1_position[6] (encoder1_position[6]), .\encoder1_position[5] (encoder1_position[5]), 
            .\encoder1_position[4] (encoder1_position[4]), .\encoder1_position[3] (encoder1_position[3]), 
            .\encoder1_position[2] (encoder1_position[2]), .n1822(n1822), 
            .VCC_net(VCC_net)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(312[49] 318[6])
    coms neopxl_color_23__I_0 (.n29968(n29968), .\data_in_frame[22] ({\data_in_frame[22] }), 
         .clk16MHz(clk16MHz), .VCC_net(VCC_net), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .\FRAME_MATCHER.i_31__N_2509 (\FRAME_MATCHER.i_31__N_2509 ), .\data_out_frame[23] ({\data_out_frame[23] }), 
         .neopxl_color({neopxl_color}), .\data_out_frame[25] ({\data_out_frame[25] }), 
         .GND_net(GND_net), .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), 
         .\data_out_frame[22] ({\data_out_frame[22] }), .\current[7] (current[7]), 
         .n51598(n51598), .n3470(n3470), .\current[6] (current[6]), .\current[5] (current[5]), 
         .n2873(n2873), .\data_out_frame[8] ({\data_out_frame[8] }), .n56908(n56908), 
         .\current[4] (current[4]), .n56907(n56907), .\current[3] (current[3]), 
         .\current[2] (current[2]), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .\current[1] (current[1]), .\current[0] (current[0]), .\data_out_frame[21] ({\data_out_frame[21] }), 
         .\current[15] (current[15]), .n52657(n52657), .\current[11] (current[11]), 
         .n57377(n57377), .n57350(n57350), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .\current[10] (current[10]), .\data_out_frame[24] ({\data_out_frame[24] }), 
         .\current[9] (current[9]), .\current[8] (current[8]), .displacement({displacement}), 
         .n59466(n59466), .n57295(n57295), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .n51730(n51730), .n51640(n51640), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .n51676(n51676), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .n57232(n57232), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .n52803(n52803), .n59193(n59193), .n57398(n57398), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .n68335(n68335), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .n68339(n68339), .\data_out_frame[11] ({\data_out_frame[11] }), 
         .\data_out_frame[12] ({\data_out_frame[12] }), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .n29959(n29959), .n51654(n51654), .n29956(n29956), .n29953(n29953), 
         .n29663(n29663), .n29949(n29949), .n29946(n29946), .n57741(n57741), 
         .\data_in_frame[3][6] (\data_in_frame[3] [6]), .\data_in_frame[3][5] (\data_in_frame[3] [5]), 
         .n25810(n25810), .n65441(n65441), .n65487(n65487), .\data_in_frame[3][4] (\data_in_frame[3] [4]), 
         .n29669(n29669), .\data_in_frame[3][3] (\data_in_frame[3] [3]), 
         .\data_in_frame[3][2] (\data_in_frame[3] [2]), .\data_in_frame[3][1] (\data_in_frame[3] [1]), 
         .n57456(n57456), .\data_in_frame[3][0] (\data_in_frame[3] [0]), 
         .\data_in_frame[2] ({\data_in_frame[2] }), .n29674(n29674), .n57131(n57131), 
         .n22726(n22726), .\data_in_frame[11] ({\data_in_frame[11] }), .\data_in_frame[17] ({\data_in_frame[17] }), 
         .\data_in_frame[8] ({\data_in_frame[8] }), .\data_in_frame[9] ({\data_in_frame[9] }), 
         .\data_out_frame[10] ({\data_out_frame[10] }), .\data_in_frame[10] ({Open_5, 
         \data_in_frame[10] [6], Open_6, \data_in_frame[10] [4], Open_7, 
         Open_8, Open_9, Open_10}), .\data_in_frame[1] ({\data_in_frame[1] }), 
         .setpoint({setpoint}), .\data_in_frame[6][5] (\data_in_frame[6] [5]), 
         .\data_out_frame[5] ({\data_out_frame[5] }), .\data_out_frame[7] ({\data_out_frame[7] }), 
         .n56906(n56906), .n56905(n56905), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .n26524(n26524), .\data_out_frame[4] ({\data_out_frame[4] }), .n56952(n56952), 
         .\data_in_frame[6][4] (\data_in_frame[6] [4]), .Kp_23__N_1748(Kp_23__N_1748), 
         .reset(reset), .n59636(n59636), .\data_in_frame[20] ({\data_in_frame[20] }), 
         .n56031(n56031), .\data_in_frame[18] ({\data_in_frame[18] }), .\data_in_frame[21] ({\data_in_frame[21] }), 
         .rx_data_ready(rx_data_ready), .rx_data({rx_data}), .n57516(n57516), 
         .n56904(n56904), .n56773(n56773), .n56903(n56903), .pwm_setpoint({pwm_setpoint}), 
         .\data_in_frame[16] ({Open_11, \data_in_frame[16] [6:3], Open_12, 
         Open_13, Open_14}), .n56902(n56902), .n56901(n56901), .n56900(n56900), 
         .n56899(n56899), .n56898(n56898), .n56897(n56897), .n56896(n56896), 
         .n56895(n56895), .n56894(n56894), .n56893(n56893), .n56892(n56892), 
         .n56891(n56891), .n56890(n56890), .n56889(n56889), .n56888(n56888), 
         .n56887(n56887), .n56886(n56886), .n56885(n56885), .n56884(n56884), 
         .n56883(n56883), .n56882(n56882), .n56881(n56881), .n56880(n56880), 
         .n56879(n56879), .n56878(n56878), .n56877(n56877), .n56876(n56876), 
         .n56875(n56875), .n56874(n56874), .n56873(n56873), .n30569(n30569), 
         .n29046(n29046), .n56872(n56872), .\data_in_frame[12] ({\data_in_frame[12] }), 
         .n26482(n26482), .n56871(n56871), .n56870(n56870), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .\FRAME_MATCHER.rx_data_ready_prev (\FRAME_MATCHER.rx_data_ready_prev ), 
         .n57917(n57917), .\data_in_frame[19] ({Open_15, \data_in_frame[19] [6], 
         Open_16, Open_17, Open_18, Open_19, Open_20, Open_21}), 
         .n56869(n56869), .n56868(n56868), .n56867(n56867), .n28417(n28417), 
         .n29684(n29684), .n8(n8_adj_5731), .n161(n161), .n10(n10_adj_5683), 
         .n10_adj_11(n10_adj_5758), .encoder0_position_scaled({encoder0_position_scaled}), 
         .\data_out_frame[26][2] (\data_out_frame[26] [2]), .\byte_transmit_counter[2] (byte_transmit_counter[2]), 
         .n29889(n29889), .n29687(n29687), .\byte_transmit_counter[1] (byte_transmit_counter[1]), 
         .encoder1_position_scaled({encoder1_position_scaled}), .n29885(n29885), 
         .n29881(n29881), .n29878(n29878), .n56866(n56866), .n56865(n56865), 
         .n56864(n56864), .\data_in_frame[15][6] (\data_in_frame[15] [6]), 
         .\data_out_frame[27][2] (\data_out_frame[27] [2]), .n56027(n56027), 
         .n56863(n56863), .n29874(n29874), .n56862(n56862), .n56861(n56861), 
         .n56860(n56860), .n59242(n59242), .n56859(n56859), .n56858(n56858), 
         .n30585(n30585), .n29030(n29030), .n56857(n56857), .n56856(n56856), 
         .n56855(n56855), .n29870(n29870), .n29867(n29867), .n28387(n28387), 
         .\FRAME_MATCHER.i[5] (\FRAME_MATCHER.i [5]), .\FRAME_MATCHER.i[3] (\FRAME_MATCHER.i [3]), 
         .\byte_transmit_counter[0] (byte_transmit_counter[0]), .n376(n376), 
         .n456(n456), .n11610(n11610), .n27692(n27692), .n29853(n29853), 
         .deadband({deadband}), .n29849(n29849), .n29848(n29848), .n29847(n29847), 
         .n29846(n29846), .n29845(n29845), .n29844(n29844), .n29843(n29843), 
         .n29842(n29842), .n29841(n29841), .n29840(n29840), .n29839(n29839), 
         .n29837(n29837), .n29836(n29836), .n29835(n29835), .n29834(n29834), 
         .n29833(n29833), .n29832(n29832), .n29831(n29831), .n29830(n29830), 
         .n29829(n29829), .n29828(n29828), .n29827(n29827), .IntegralLimit({IntegralLimit}), 
         .n29826(n29826), .n29825(n29825), .n29824(n29824), .n29823(n29823), 
         .n29822(n29822), .n29821(n29821), .n29820(n29820), .n29819(n29819), 
         .n29818(n29818), .n29817(n29817), .n29816(n29816), .n29815(n29815), 
         .n29814(n29814), .n29813(n29813), .n29812(n29812), .n29811(n29811), 
         .n29810(n29810), .n29809(n29809), .n29808(n29808), .n29807(n29807), 
         .n29806(n29806), .n29805(n29805), .n29804(n29804), .\Kp[1] (Kp[1]), 
         .n29803(n29803), .\Kp[2] (Kp[2]), .n29802(n29802), .\Kp[3] (Kp[3]), 
         .\pwm_counter[22] (pwm_counter[22]), .n45(n45), .\pwm_counter[21] (pwm_counter[21]), 
         .n43(n43), .n29801(n29801), .\Kp[4] (Kp[4]), .n29800(n29800), 
         .\Kp[5] (Kp[5]), .n29799(n29799), .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), 
         .n29797(n29797), .\Kp[8] (Kp[8]), .n29796(n29796), .\Kp[9] (Kp[9]), 
         .n29795(n29795), .\Kp[10] (Kp[10]), .n29794(n29794), .\Kp[11] (Kp[11]), 
         .n29793(n29793), .\Kp[12] (Kp[12]), .n29792(n29792), .\Kp[13] (Kp[13]), 
         .n29791(n29791), .\Kp[14] (Kp[14]), .n29790(n29790), .\Kp[15] (Kp[15]), 
         .n29789(n29789), .\Ki[1] (Ki[1]), .n29788(n29788), .\Ki[2] (Ki[2]), 
         .n29787(n29787), .\Ki[3] (Ki[3]), .n29786(n29786), .\Ki[4] (Ki[4]), 
         .n29785(n29785), .\Ki[5] (Ki[5]), .n29784(n29784), .\Ki[6] (Ki[6]), 
         .n29783(n29783), .\Ki[7] (Ki[7]), .n29782(n29782), .\Ki[8] (Ki[8]), 
         .n29781(n29781), .\Ki[9] (Ki[9]), .n29780(n29780), .\Ki[10] (Ki[10]), 
         .n29779(n29779), .\Ki[11] (Ki[11]), .n29778(n29778), .\Ki[12] (Ki[12]), 
         .n29777(n29777), .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), .n29775(n29775), 
         .\Ki[15] (Ki[15]), .n56854(n56854), .n56853(n56853), .n56852(n56852), 
         .n56851(n56851), .n56850(n56850), .n56849(n56849), .n56775(n56775), 
         .n56777(n56777), .n57044(n57044), .n56778(n56778), .n56779(n56779), 
         .n56780(n56780), .n56781(n56781), .n56783(n56783), .n56784(n56784), 
         .n56785(n56785), .n56786(n56786), .n56787(n56787), .n56788(n56788), 
         .n29746(n29746), .n56789(n56789), .n56790(n56790), .n56791(n56791), 
         .n56792(n56792), .n29736(n29736), .n56793(n56793), .n56774(n56774), 
         .n56794(n56794), .n56795(n56795), .n56796(n56796), .n29735(n29735), 
         .current_limit({current_limit}), .n29734(n29734), .control_mode({control_mode}), 
         .n29733(n29733), .n29732(n29732), .n29731(n29731), .n56797(n56797), 
         .n56798(n56798), .n29727(n29727), .n29726(n29726), .n29725(n29725), 
         .n29723(n29723), .n29722(n29722), .n29721(n29721), .n29720(n29720), 
         .n29719(n29719), .n29718(n29718), .n29717(n29717), .n56799(n56799), 
         .n56800(n56800), .n29716(n29716), .n29712(n29712), .n29711(n29711), 
         .n56801(n56801), .n56802(n56802), .n29708(n29708), .n29707(n29707), 
         .n56803(n56803), .n29706(n29706), .n29705(n29705), .n29703(n29703), 
         .n29702(n29702), .n29698(n29698), .n29694(n29694), .n40973(n40973), 
         .n28438(n28438), .n29691(n29691), .Kp_23__N_1301(Kp_23__N_1301), 
         .n57039(n57039), .\data_in_frame[15][7] (\data_in_frame[15] [7]), 
         .\data_in_frame[15][4] (\data_in_frame[15] [4]), .n57780(n57780), 
         .n29673(n29673), .n29672(n29672), .n29662(n29662), .n29644(n29644), 
         .PWMLimit({PWMLimit}), .n29639(n29639), .n29638(n29638), .n29637(n29637), 
         .n29636(n29636), .\Ki[0] (Ki[0]), .n29635(n29635), .\Kp[0] (Kp[0]), 
         .n29613(n29613), .n56804(n56804), .n56805(n56805), .n56806(n56806), 
         .n30647(n30647), .n28989(n28989), .n56807(n56807), .n30649(n30649), 
         .n28987(n28987), .n56808(n56808), .n56809(n56809), .n56810(n56810), 
         .n56811(n56811), .n56812(n56812), .n30655(n30655), .n28981(n28981), 
         .n56813(n56813), .n56814(n56814), .n56815(n56815), .n56816(n56816), 
         .n56817(n56817), .n56818(n56818), .n56819(n56819), .n56820(n56820), 
         .n56821(n56821), .n56822(n56822), .n56823(n56823), .n56824(n56824), 
         .n56825(n56825), .n8_adj_12(n8_adj_5760), .n56826(n56826), .n56827(n56827), 
         .n56828(n56828), .n56829(n56829), .n56830(n56830), .n56831(n56831), 
         .\data_out_frame[0][2] (\data_out_frame[0] [2]), .n56951(n56951), 
         .\data_out_frame[0][3] (\data_out_frame[0] [3]), .n56950(n56950), 
         .\data_out_frame[0][4] (\data_out_frame[0] [4]), .n56949(n56949), 
         .\data_out_frame[1][0] (\data_out_frame[1] [0]), .n56948(n56948), 
         .\data_in_frame[16][7] (\data_in_frame[16] [7]), .\data_in_frame[19][3] (\data_in_frame[19] [3]), 
         .n57717(n57717), .\data_out_frame[1][1] (\data_out_frame[1] [1]), 
         .n56947(n56947), .\data_out_frame[1][3] (\data_out_frame[1] [3]), 
         .n56946(n56946), .\data_out_frame[1][5] (\data_out_frame[1] [5]), 
         .n56945(n56945), .\data_in_frame[15][1] (\data_in_frame[15] [1]), 
         .\data_in_frame[14] ({\data_in_frame[14] }), .n25864(n25864), .n57720(n57720), 
         .\data_out_frame[1][6] (\data_out_frame[1] [6]), .n56944(n56944), 
         .\data_in_frame[19][4] (\data_in_frame[19] [4]), .\data_out_frame[1][7] (\data_out_frame[1] [7]), 
         .n56943(n56943), .\data_out_frame[3][1] (\data_out_frame[3] [1]), 
         .n56942(n56942), .\data_in_frame[15][3] (\data_in_frame[15] [3]), 
         .n30519(n30519), .n30518(n30518), .n30517(n30517), .n30515(n30515), 
         .n30514(n30514), .n30513(n30513), .n30512(n30512), .\data_in_frame[15][0] (\data_in_frame[15] [0]), 
         .\data_in_frame[15][2] (\data_in_frame[15] [2]), .n30470(n30470), 
         .n30468(n30468), .n30467(n30467), .n30466(n30466), .n30465(n30465), 
         .n30464(n30464), .n30444(n30444), .n30398(n30398), .n30396(n30396), 
         .n30395(n30395), .n30384(n30384), .n30375(n30375), .\data_out_frame[3][3] (\data_out_frame[3] [3]), 
         .n56941(n56941), .n25952(n25952), .\data_out_frame[3][4] (\data_out_frame[3] [4]), 
         .n56940(n56940), .n30350(n30350), .n30349(n30349), .n30348(n30348), 
         .n30347(n30347), .n29973(n29973), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .n29976(n29976), .n30343(n30343), .n29979(n29979), .n29982(n29982), 
         .n56201(n56201), .\data_in_frame[16][1] (\data_in_frame[16] [1]), 
         .n30339(n30339), .n56199(n56199), .\data_in_frame[16][2] (\data_in_frame[16] [2]), 
         .n29490(n29490), .n29493(n29493), .n29496(n29496), .n29499(n29499), 
         .n56249(n56249), .n56107(n56107), .n56103(n56103), .n56101(n56101), 
         .n56099(n56099), .n56095(n56095), .n56091(n56091), .\data_out_frame[3][6] (\data_out_frame[3] [6]), 
         .n56771(n56771), .n29986(n29986), .n29989(n29989), .n29992(n29992), 
         .n56087(n56087), .n56083(n56083), .n56079(n56079), .n30305(n30305), 
         .n29995(n29995), .\data_in_frame[6][0] (\data_in_frame[6] [0]), 
         .\data_in_frame[6][1] (\data_in_frame[6] [1]), .\data_in_frame[6][2] (\data_in_frame[6] [2]), 
         .\data_in_frame[6][3] (\data_in_frame[6] [3]), .n30299(n30299), 
         .\data_out_frame[3][7] (\data_out_frame[3] [7]), .n56939(n56939), 
         .n30047(n30047), .n30050(n30050), .n30054(n30054), .n30057(n30057), 
         .n30282(n30282), .n30281(n30281), .n30280(n30280), .n30063(n30063), 
         .n30066(n30066), .n30069(n30069), .n30072(n30072), .n30075(n30075), 
         .n30079(n30079), .n30082(n30082), .n30085(n30085), .n30089(n30089), 
         .n30092(n30092), .n30095(n30095), .\data_in_frame[10][1] (\data_in_frame[10] [1]), 
         .\data_in_frame[10][2] (\data_in_frame[10] [2]), .\data_in_frame[10][3] (\data_in_frame[10] [3]), 
         .\data_in_frame[10][5] (\data_in_frame[10] [5]), .\data_in_frame[10][7] (\data_in_frame[10] [7]), 
         .n30149(n30149), .n30152(n30152), .n30250(n30250), .n30156(n30156), 
         .n56303(n56303), .n56343(n56343), .n30166(n30166), .n30169(n30169), 
         .n30172(n30172), .n30176(n30176), .n30179(n30179), .n30182(n30182), 
         .n30186(n30186), .n30189(n30189), .n30192(n30192), .n30196(n30196), 
         .n56075(n56075), .n56071(n56071), .n30232(n30232), .n29540(n29540), 
         .n29543(n29543), .n29546(n29546), .n56065(n56065), .n56061(n56061), 
         .n56057(n56057), .\data_in_frame[19][0] (\data_in_frame[19] [0]), 
         .n56053(n56053), .\data_in_frame[19][1] (\data_in_frame[19] [1]), 
         .n56049(n56049), .\data_in_frame[19][2] (\data_in_frame[19] [2]), 
         .n30207(n30207), .n56045(n56045), .n56041(n56041), .\data_in_frame[19][5] (\data_in_frame[19] [5]), 
         .n56037(n56037), .n29579(n29579), .n29588(n29588), .n29591(n29591), 
         .n29594(n29594), .n30155(n30155), .n57701(n57701), .n29600(n29600), 
         .n57361(n57361), .n57467(n57467), .n56938(n56938), .n172(n172), 
         .n33761(n33761), .n30739(n30739), .n29117(n29117), .n30740(n30740), 
         .n29116(n29116), .n30741(n30741), .n29115(n29115), .n56937(n56937), 
         .n59574(n59574), .n29509(n29509), .n10_adj_13(n10_adj_5903), 
         .n56936(n56936), .n56935(n56935), .n57473(n57473), .\FRAME_MATCHER.i_31__N_2513 (\FRAME_MATCHER.i_31__N_2513 ), 
         .n56934(n56934), .n56933(n56933), .n56932(n56932), .n56931(n56931), 
         .n56930(n56930), .n56929(n56929), .n56928(n56928), .n56927(n56927), 
         .n56926(n56926), .n56925(n56925), .n56924(n56924), .n56923(n56923), 
         .n56922(n56922), .n56921(n56921), .n56920(n56920), .n56919(n56919), 
         .n29480(n29480), .n57125(n57125), .n57680(n57680), .n29478(n29478), 
         .n56832(n56832), .n56833(n56833), .n56834(n56834), .n56835(n56835), 
         .n56836(n56836), .n56837(n56837), .n56838(n56838), .n56839(n56839), 
         .n56840(n56840), .n56772(n56772), .n56782(n56782), .n56841(n56841), 
         .n56842(n56842), .n56843(n56843), .n56844(n56844), .n56918(n56918), 
         .n56917(n56917), .n56916(n56916), .n56915(n56915), .n56845(n56845), 
         .n56846(n56846), .n56847(n56847), .n56848(n56848), .n56776(n56776), 
         .LED_c(LED_c), .n56914(n56914), .DE_c(DE_c), .n56913(n56913), 
         .n56912(n56912), .n56911(n56911), .n56910(n56910), .n29969(n29969), 
         .n56909(n56909), .n92(n92), .ID({ID}), .n33769(n33769), .n27696(n27696), 
         .n28383(n28383), .n28379(n28379), .n28434(n28434), .n26(n26), 
         .n21(n21_adj_5850), .tx_active(tx_active), .n57921(n57921), .n260(n260), 
         .n8_adj_14(n8_adj_5786), .n130(n130), .n65436(n65436), .n28428(n28428), 
         .n59230(n59230), .n375(n375), .n455(n455), .n37189(n37189), 
         .n15(n15_adj_5681), .n15_adj_15(n15), .n19(n19_adj_5811), .n28375(n28375), 
         .n56988(n56988), .n8_adj_16(n8_adj_5741), .n28381(n28381), .n69525(n69525), 
         .n4(n4_adj_5818), .n4_adj_17(n4_adj_5821), .n30(n30_adj_5819), 
         .n361(n361), .n32(n32_adj_5820), .n69309(n69309), .n25(n25_adj_5803), 
         .n134(n134), .n20(n20_adj_5848), .n43_adj_18(n43_adj_5825), .n401(n401), 
         .n4_adj_19(n4_adj_5817), .n65432(n65432), .n69489(n69489), .n62711(n62711), 
         .n62712(n62712), .n62859(n62859), .n62858(n62858), .n52677(n52677), 
         .r_SM_Main({r_SM_Main_adj_5986}), .n57935(n57935), .n6(n6_adj_5891), 
         .tx_o(tx_o), .n29661(n29661), .r_Clock_Count({r_Clock_Count_adj_5987}), 
         .n4940(n4940), .n27(n27_adj_5781), .tx_enable(tx_enable), .\r_Bit_Index[0] (r_Bit_Index[0]), 
         .n4937(n4937), .\o_Rx_DV_N_3488[8] (o_Rx_DV_N_3488[8]), .n60724(n60724), 
         .baudrate({baudrate}), .\r_SM_Main[2]_adj_20 (r_SM_Main[2]), .n25530(n25530), 
         .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), .\r_SM_Main[1]_adj_21 (r_SM_Main[1]), 
         .n27966(n27966), .n56959(n56959), .n60740(n60740), .n29884(n29884), 
         .n60788(n60788), .n60756(n60756), .n29866(n29866), .\o_Rx_DV_N_3488[7] (o_Rx_DV_N_3488[7]), 
         .\o_Rx_DV_N_3488[6] (o_Rx_DV_N_3488[6]), .\o_Rx_DV_N_3488[5] (o_Rx_DV_N_3488[5]), 
         .\o_Rx_DV_N_3488[4] (o_Rx_DV_N_3488[4]), .\o_Rx_DV_N_3488[3] (o_Rx_DV_N_3488[3]), 
         .\o_Rx_DV_N_3488[2] (o_Rx_DV_N_3488[2]), .\o_Rx_DV_N_3488[1] (o_Rx_DV_N_3488[1]), 
         .\o_Rx_DV_N_3488[0] (o_Rx_DV_N_3488[0]), .n29774(n29774), .n29773(n29773), 
         .n29772(n29772), .r_Clock_Count_adj_30({r_Clock_Count}), .n58000(n58000), 
         .n30502(n30502), .n52851(n52851), .n30498(n30498), .n30201(n30201), 
         .n30200(n30200), .n60708(n60708), .n60692(n60692), .n60804(n60804), 
         .n27724(n27724), .n60772(n60772)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(255[22] 280[4])
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[23] [1]), .I1(\data_out_frame[18] [5]), 
            .I2(\data_out_frame[16] [1]), .I3(GND_net), .O(n10_adj_5823));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i16647_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [1]), 
            .O(n30655));   // verilog/coms.v(130[12] 305[6])
    defparam i16647_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_30__I_0_i1104_3_lut (.I0(n1621), .I1(n1688), 
            .I2(n1653), .I3(GND_net), .O(n1720));   // verilog/TinyFPGA_B.v(321[33:59])
    defparam encoder0_position_30__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16641_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [3]), 
            .O(n30649));   // verilog/coms.v(130[12] 305[6])
    defparam i16641_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    pwm PWM (.n2873(n2873), .pwm_out(pwm_out), .clk32MHz(clk32MHz), .pwm_setpoint({pwm_setpoint}), 
        .GND_net(GND_net), .n45(n45), .n43(n43), .reset(reset), .\pwm_counter[22] (pwm_counter[22]), 
        .\pwm_counter[21] (pwm_counter[21]), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(97[6] 102[3])
    SB_LUT4 i16639_2_lut_2_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [1]), 
            .O(n30647));   // verilog/coms.v(130[12] 305[6])
    defparam i16639_2_lut_2_lut_4_lut.LUT_INIT = 16'h5555;
    TLI4970 tli (.\state[1] (state_adj_5976[1]), .\state[0] (state_adj_5976[0]), 
            .GND_net(GND_net), .n6(n6_adj_5732), .n5(n5_adj_5784), .n6_adj_8(n6_adj_5730), 
            .n42774(n42774), .state_7__N_4317(state_7__N_4317), .n42779(n42779), 
            .\data[15] (data_adj_5974[15]), .n27706(n27706), .clk16MHz(clk16MHz), 
            .n11(n11_adj_5734), .n9(n9_adj_5910), .clk_out(clk_out), .n29648(n29648), 
            .CS_c(CS_c), .n29646(n29646), .\current[0] (current[0]), .n29643(n29643), 
            .n29628(n29628), .\data[12] (data_adj_5974[12]), .n29627(n29627), 
            .\data[11] (data_adj_5974[11]), .n29626(n29626), .\data[10] (data_adj_5974[10]), 
            .n29625(n29625), .\data[9] (data_adj_5974[9]), .n29624(n29624), 
            .\data[8] (data_adj_5974[8]), .n29617(n29617), .\data[7] (data_adj_5974[7]), 
            .n29612(n29612), .\data[6] (data_adj_5974[6]), .n29608(n29608), 
            .\data[5] (data_adj_5974[5]), .n29607(n29607), .\data[4] (data_adj_5974[4]), 
            .n29606(n29606), .\data[3] (data_adj_5974[3]), .n29605(n29605), 
            .\data[2] (data_adj_5974[2]), .n29604(n29604), .\data[1] (data_adj_5974[1]), 
            .VCC_net(VCC_net), .n30506(n30506), .\data[0] (data_adj_5974[0]), 
            .n30394(n30394), .\current[1] (current[1]), .n30393(n30393), 
            .\current[2] (current[2]), .n30392(n30392), .\current[3] (current[3]), 
            .n30391(n30391), .\current[4] (current[4]), .n30390(n30390), 
            .\current[5] (current[5]), .n30389(n30389), .\current[6] (current[6]), 
            .n30388(n30388), .\current[7] (current[7]), .n30387(n30387), 
            .\current[8] (current[8]), .n30386(n30386), .\current[9] (current[9]), 
            .n30385(n30385), .\current[10] (current[10]), .n30383(n30383), 
            .\current[11] (current[11]), .\current[15] (current[15]), .CS_CLK_c(CS_CLK_c), 
            .n6_adj_9(n6), .n5_adj_10(n5_adj_5708), .n15(n15_adj_5733), 
            .n25532(n25532), .n25571(n25571), .n25523(n25523), .n25519(n25519), 
            .n4(n4_adj_5783), .n25527(n25527)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(404[11] 410[4])
    EEPROM eeprom (.\state[1] (state_adj_5967[1]), .\state[0] (state_adj_5967[0]), 
           .n3(n3_adj_5845), .\state[2] (state_adj_5967[2]), .GND_net(GND_net), 
           .enable_slow_N_4211(enable_slow_N_4211), .ready_prev(ready_prev), 
           .n42699(n42699), .n57012(n57012), .n25516(n25516), .data({data_adj_5966}), 
           .ID({ID}), .clk16MHz(clk16MHz), .n5773({n5774}), .n25404(n25404), 
           .n27997(n27997), .n29647(n29647), .rw(rw), .n56425(n56425), 
           .data_ready(data_ready), .n55999(n55999), .n56203(n56203), 
           .baudrate({baudrate}), .n30406(n30406), .n30405(n30405), .n30404(n30404), 
           .n30403(n30403), .n30402(n30402), .n30401(n30401), .n30400(n30400), 
           .n30399(n30399), .\state_7__N_3916[0] (state_7__N_3916[0]), .\state[0]_adj_4 (state_adj_5997[0]), 
           .n4(n4_adj_5842), .scl_enable(scl_enable), .n6428(n6428), .\state_7__N_4108[0] (state_7__N_4108[0]), 
           .scl(scl), .sda_enable(sda_enable), .sda_out(sda_out), .n29654(n29654), 
           .\saved_addr[0] (saved_addr[0]), .VCC_net(VCC_net), .n30492(n30492), 
           .n8(n8_adj_5911), .n30216(n30216), .n30215(n30215), .n30214(n30214), 
           .n30213(n30213), .n30212(n30212), .n30211(n30211), .n30210(n30210), 
           .n4_adj_5(n4_adj_5727), .n4_adj_6(n4_adj_5728), .n65481(n65481), 
           .n42804(n42804), .n10(n10_adj_5729), .n25540(n25540), .n25535(n25535), 
           .\state_7__N_4124[3] (state_7__N_4124[3]), .n10_adj_7(n10_adj_5844)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(390[10] 402[6])
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (timer, GND_net, clk16MHz, 
            state, n25, VCC_net, bit_ctr, neopxl_color, n111, \neo_pixel_transmitter.t0 , 
            n29677, n27920, n30323, n30322, n30321, n30320, n30319, 
            n30318, n30317, n30316, n30315, n30308, n30221, n5, 
            NEOPXL_c, LED_c, n43462, n23) /* synthesis syn_module_defined=1 */ ;
    output [10:0]timer;
    input GND_net;
    input clk16MHz;
    output [1:0]state;
    output n25;
    input VCC_net;
    output [4:0]bit_ctr;
    input [23:0]neopxl_color;
    output n111;
    output [10:0]\neo_pixel_transmitter.t0 ;
    input n29677;
    output n27920;
    input n30323;
    input n30322;
    input n30321;
    input n30320;
    input n30319;
    input n30318;
    input n30317;
    input n30316;
    input n30315;
    input n30308;
    input n30221;
    input n5;
    output NEOPXL_c;
    input LED_c;
    output n43462;
    output n23;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [10:0]one_wire_N_479;
    wire [10:0]n13;
    
    wire n49187, \neo_pixel_transmitter.done_N_516 , n60204, \neo_pixel_transmitter.done , 
        start_N_507, n7, start, n112, n59, n33, n57929, n49188, 
        n49186, n49185, n58002, n4, n69162;
    wire [4:0]bit_ctr_c;   // verilog/neopixel.v(17[11:18])
    wire [31:0]n137;
    
    wire n69492, n58018, n57931, n51273, n115, n41, n62468, n65451, 
        n40745, n7_adj_5650, n8;
    wire [10:0]n49;
    
    wire n29169, n50403, n50402, n50401, n50400, n50399, n50398, 
        n50397, n50396, n50395, n50394, n1, n27910, n28881;
    wire [1:0]state_1__N_440;
    
    wire n27924, n29173, \neo_pixel_transmitter.done_N_524 , n27677, 
        n60211, n49194, n49193, n49192, n49191, n49190, n6_adj_5654, 
        n49189, n62792, n62793, n62796, n62795, n62852, n62853, 
        n62865, n62864, n57801, n43356, n51740;
    wire [5:0]color_bit_N_502;
    
    wire n6897, n25492, n25491, n69327, n65478, n69273, n67521, 
        n67668, n65449, n69324, n58040, n48, n54_adj_5657, n69165, 
        n69495, n69270, n41_adj_5658;
    
    SB_LUT4 sub_67_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n13[3]), 
            .I3(n49187), .O(one_wire_N_479[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFE \neo_pixel_transmitter.done_96  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk16MHz), .E(n60204), .D(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFE start_95 (.Q(start), .C(clk16MHz), .E(n7), .D(start_N_507));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 i1_4_lut (.I0(n112), .I1(n59), .I2(state[0]), .I3(\neo_pixel_transmitter.done ), 
            .O(n33));
    defparam i1_4_lut.LUT_INIT = 16'hdccd;
    SB_LUT4 i1_4_lut_adj_1807 (.I0(state[1]), .I1(n33), .I2(n57929), .I3(start), 
            .O(n25));
    defparam i1_4_lut_adj_1807.LUT_INIT = 16'haaae;
    SB_CARRY sub_67_add_2_5 (.CI(n49187), .I0(timer[3]), .I1(n13[3]), 
            .CO(n49188));
    SB_LUT4 sub_67_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n13[2]), 
            .I3(n49186), .O(one_wire_N_479[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n13[0]), 
            .CO(n49185));
    SB_CARRY sub_67_add_2_4 (.CI(n49186), .I0(timer[2]), .I1(n13[2]), 
            .CO(n49187));
    SB_LUT4 sub_67_add_2_3_lut (.I0(n4), .I1(timer[1]), .I2(n13[1]), .I3(n49185), 
            .O(n58002)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 bit_ctr_0__bdd_4_lut_53746_4_lut_4_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), 
            .I2(neopxl_color[13]), .I3(neopxl_color[12]), .O(n69162));   // verilog/neopixel.v(18[6:15])
    defparam bit_ctr_0__bdd_4_lut_53746_4_lut_4_lut.LUT_INIT = 16'hd5c4;
    SB_LUT4 i2094_2_lut_3_lut (.I0(bit_ctr_c[2]), .I1(bit_ctr[1]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n137[2]));   // verilog/neopixel.v(68[23:32])
    defparam i2094_2_lut_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 bit_ctr_0__bdd_4_lut_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n69492));
    defparam bit_ctr_0__bdd_4_lut_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 i42380_2_lut_3_lut (.I0(state[1]), .I1(start), .I2(n57929), 
            .I3(GND_net), .O(n58018));
    defparam i42380_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut (.I0(n58002), .I1(\neo_pixel_transmitter.done ), .I2(state[0]), 
            .I3(GND_net), .O(n59));
    defparam i1_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i42276_2_lut (.I0(one_wire_N_479[3]), .I1(one_wire_N_479[2]), 
            .I2(GND_net), .I3(GND_net), .O(n112));
    defparam i42276_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i42294_2_lut (.I0(state[1]), .I1(start), .I2(GND_net), .I3(GND_net), 
            .O(n57931));
    defparam i42294_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY sub_67_add_2_3 (.CI(n49185), .I0(timer[1]), .I1(n13[1]), 
            .CO(n49186));
    SB_LUT4 i1_4_lut_adj_1808 (.I0(n58002), .I1(n57929), .I2(n112), .I3(state[0]), 
            .O(n51273));   // verilog/neopixel.v(16[11:16])
    defparam i1_4_lut_adj_1808.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_2_lut (.I0(one_wire_N_479[10]), .I1(n115), .I2(GND_net), 
            .I3(GND_net), .O(n41));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i53453_4_lut (.I0(n62468), .I1(n112), .I2(one_wire_N_479[7]), 
            .I3(n59), .O(n60204));
    defparam i53453_4_lut.LUT_INIT = 16'hfafe;
    SB_LUT4 i15_4_lut (.I0(n65451), .I1(n40745), .I2(state[1]), .I3(state[0]), 
            .O(n7));
    defparam i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i50584_2_lut_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(n51273), 
            .I2(start), .I3(GND_net), .O(n65451));   // verilog/neopixel.v(16[11:16])
    defparam i50584_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i1_2_lut_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(n51273), 
            .I2(start), .I3(GND_net), .O(n111));   // verilog/neopixel.v(16[11:16])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i53221_2_lut (.I0(start), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(start_N_507));   // verilog/neopixel.v(35[4] 115[11])
    defparam i53221_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i46791_2_lut_3_lut (.I0(n7_adj_5650), .I1(n8), .I2(n57931), 
            .I3(GND_net), .O(n62468));   // verilog/neopixel.v(101[14:24])
    defparam i46791_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i42292_2_lut_3_lut (.I0(n7_adj_5650), .I1(n8), .I2(one_wire_N_479[7]), 
            .I3(GND_net), .O(n57929));   // verilog/neopixel.v(101[14:24])
    defparam i42292_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i26815_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[1]), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(16[11:16])
    defparam i26815_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 i1_2_lut_adj_1809 (.I0(one_wire_N_479[2]), .I1(one_wire_N_479[3]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/neopixel.v(101[14:24])
    defparam i1_2_lut_adj_1809.LUT_INIT = 16'h8888;
    SB_LUT4 sub_67_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[1]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_DFF timer_1938__i0 (.Q(timer[0]), .C(clk16MHz), .D(n49[0]));   // verilog/neopixel.v(12[12:21])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk16MHz), .D(n29677));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR bit_ctr_i2 (.Q(bit_ctr_c[2]), .C(clk16MHz), .E(n27920), 
            .D(n137[2]), .R(n29169));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR bit_ctr_i3 (.Q(bit_ctr_c[3]), .C(clk16MHz), .E(n27920), 
            .D(n137[3]), .R(n29169));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR bit_ctr_i4 (.Q(bit_ctr_c[4]), .C(clk16MHz), .E(n27920), 
            .D(n137[4]), .R(n29169));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF timer_1938__i10 (.Q(timer[10]), .C(clk16MHz), .D(n49[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1938__i9 (.Q(timer[9]), .C(clk16MHz), .D(n49[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1938__i8 (.Q(timer[8]), .C(clk16MHz), .D(n49[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1938__i7 (.Q(timer[7]), .C(clk16MHz), .D(n49[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1938__i6 (.Q(timer[6]), .C(clk16MHz), .D(n49[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1938__i5 (.Q(timer[5]), .C(clk16MHz), .D(n49[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1938__i4 (.Q(timer[4]), .C(clk16MHz), .D(n49[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1938__i3 (.Q(timer[3]), .C(clk16MHz), .D(n49[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1938__i2 (.Q(timer[2]), .C(clk16MHz), .D(n49[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1938__i1 (.Q(timer[1]), .C(clk16MHz), .D(n49[1]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 timer_1938_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n50403), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1938_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n50402), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_11 (.CI(n50402), .I0(GND_net), .I1(timer[9]), 
            .CO(n50403));
    SB_LUT4 timer_1938_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n50401), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_10 (.CI(n50401), .I0(GND_net), .I1(timer[8]), 
            .CO(n50402));
    SB_LUT4 timer_1938_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n50400), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_9 (.CI(n50400), .I0(GND_net), .I1(timer[7]), 
            .CO(n50401));
    SB_LUT4 timer_1938_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n50399), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_8 (.CI(n50399), .I0(GND_net), .I1(timer[6]), 
            .CO(n50400));
    SB_LUT4 timer_1938_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n50398), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_7 (.CI(n50398), .I0(GND_net), .I1(timer[5]), 
            .CO(n50399));
    SB_LUT4 timer_1938_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n50397), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_6 (.CI(n50397), .I0(GND_net), .I1(timer[4]), 
            .CO(n50398));
    SB_LUT4 timer_1938_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n50396), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_5 (.CI(n50396), .I0(GND_net), .I1(timer[3]), 
            .CO(n50397));
    SB_LUT4 timer_1938_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n50395), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_4 (.CI(n50395), .I0(GND_net), .I1(timer[2]), 
            .CO(n50396));
    SB_LUT4 timer_1938_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n50394), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_3 (.CI(n50394), .I0(GND_net), .I1(timer[1]), 
            .CO(n50395));
    SB_LUT4 timer_1938_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1938_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1938_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n50394));
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk16MHz), .D(n30323));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk16MHz), .D(n30322));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk16MHz), .D(n30321));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk16MHz), .D(n30320));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk16MHz), .D(n30319));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk16MHz), .D(n30318));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk16MHz), .D(n30317));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk16MHz), .D(n30316));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk16MHz), .D(n30315));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk16MHz), .D(n30308));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFF bit_ctr_i1 (.Q(bit_ctr[1]), .C(clk16MHz), .D(n30221));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(VCC_net), .D(n5));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR bit_ctr_i0 (.Q(bit_ctr[0]), .C(clk16MHz), .E(n27910), .D(n1), 
            .R(n28881));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESS state_i0 (.Q(state[0]), .C(clk16MHz), .E(n27924), .D(state_1__N_440[0]), 
            .S(n29173));   // verilog/neopixel.v(34[12] 116[6])
    SB_DFFESR one_wire_99 (.Q(NEOPXL_c), .C(clk16MHz), .E(n27677), .D(\neo_pixel_transmitter.done_N_524 ), 
            .R(n60211));   // verilog/neopixel.v(34[12] 116[6])
    SB_LUT4 sub_67_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[3]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n13[10]), 
            .I3(n49194), .O(one_wire_N_479[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_67_add_2_11_lut (.I0(one_wire_N_479[8]), .I1(timer[9]), 
            .I2(n13[9]), .I3(n49193), .O(n115)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_11_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_67_add_2_11 (.CI(n49193), .I0(timer[9]), .I1(n13[9]), 
            .CO(n49194));
    SB_LUT4 sub_67_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n13[8]), 
            .I3(n49192), .O(one_wire_N_479[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_10 (.CI(n49192), .I0(timer[8]), .I1(n13[8]), 
            .CO(n49193));
    SB_LUT4 sub_67_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n13[7]), 
            .I3(n49191), .O(one_wire_N_479[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_67_add_2_9 (.CI(n49191), .I0(timer[7]), .I1(n13[7]), 
            .CO(n49192));
    SB_LUT4 sub_67_add_2_8_lut (.I0(one_wire_N_479[10]), .I1(timer[6]), 
            .I2(n13[6]), .I3(n49190), .O(n7_adj_5650)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_67_add_2_8 (.CI(n49190), .I0(timer[6]), .I1(n13[6]), 
            .CO(n49191));
    SB_LUT4 sub_67_add_2_7_lut (.I0(n115), .I1(timer[5]), .I2(n13[5]), 
            .I3(n49189), .O(n6_adj_5654)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_7_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_67_add_2_7 (.CI(n49189), .I0(timer[5]), .I1(n13[5]), 
            .CO(n49190));
    SB_LUT4 sub_67_add_2_6_lut (.I0(n6_adj_5654), .I1(timer[4]), .I2(n13[4]), 
            .I3(n49188), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_67_add_2_6_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_67_add_2_6 (.CI(n49188), .I0(timer[4]), .I1(n13[4]), 
            .CO(n49189));
    SB_LUT4 i47106_3_lut (.I0(neopxl_color[0]), .I1(neopxl_color[1]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n62792));
    defparam i47106_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47107_3_lut (.I0(neopxl_color[2]), .I1(neopxl_color[3]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n62793));
    defparam i47107_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47110_3_lut (.I0(neopxl_color[6]), .I1(neopxl_color[7]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n62796));
    defparam i47110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47109_3_lut (.I0(neopxl_color[4]), .I1(neopxl_color[5]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n62795));
    defparam i47109_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47166_3_lut (.I0(neopxl_color[16]), .I1(neopxl_color[17]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n62852));
    defparam i47166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47167_3_lut (.I0(neopxl_color[18]), .I1(neopxl_color[19]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n62853));
    defparam i47167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47179_3_lut (.I0(neopxl_color[22]), .I1(neopxl_color[23]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n62865));
    defparam i47179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47178_3_lut (.I0(neopxl_color[20]), .I1(neopxl_color[21]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n62864));
    defparam i47178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_4_lut (.I0(n111), .I1(state[1]), .I2(n40745), .I3(state[0]), 
            .O(n27924));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'heee2;
    SB_LUT4 i1_2_lut_3_lut_adj_1810 (.I0(n111), .I1(state[1]), .I2(n27910), 
            .I3(GND_net), .O(n27920));
    defparam i1_2_lut_3_lut_adj_1810.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[0]), .I1(LED_c), .I2(n57801), .I3(state[1]), 
            .O(n27910));   // verilog/neopixel.v(34[12] 116[6])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h80ff;
    SB_LUT4 i14873_2_lut_4_lut (.I0(state[0]), .I1(LED_c), .I2(n57801), 
            .I3(state[1]), .O(n28881));   // verilog/neopixel.v(34[12] 116[6])
    defparam i14873_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i29554_2_lut_3_lut (.I0(bit_ctr_c[3]), .I1(n43356), .I2(bit_ctr_c[4]), 
            .I3(GND_net), .O(n43462));
    defparam i29554_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1811 (.I0(bit_ctr_c[3]), .I1(n43356), .I2(bit_ctr_c[4]), 
            .I3(GND_net), .O(n51740));
    defparam i1_2_lut_3_lut_adj_1811.LUT_INIT = 16'h7878;
    SB_LUT4 sub_67_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[4]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_adj_1812 (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr_c[2]), 
            .I3(GND_net), .O(color_bit_N_502[2]));
    defparam i1_2_lut_3_lut_adj_1812.LUT_INIT = 16'h1e1e;
    SB_LUT4 i1_2_lut_adj_1813 (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(color_bit_N_502[1]));
    defparam i1_2_lut_adj_1813.LUT_INIT = 16'h6666;
    SB_LUT4 i29451_2_lut_3_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr_c[2]), 
            .I3(GND_net), .O(n43356));
    defparam i29451_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 sub_67_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[5]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2108_3_lut_4_lut (.I0(bit_ctr_c[2]), .I1(n6897), .I2(bit_ctr_c[3]), 
            .I3(bit_ctr_c[4]), .O(n137[4]));   // verilog/neopixel.v(68[23:32])
    defparam i2108_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 sub_67_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[6]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_4_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(n57929), .I3(n112), .O(n25492));   // verilog/neopixel.v(34[12] 116[6])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hbbbf;
    SB_LUT4 i1_3_lut_4_lut_adj_1814 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(n57929), .I3(n58002), .O(n25491));   // verilog/neopixel.v(34[12] 116[6])
    defparam i1_3_lut_4_lut_adj_1814.LUT_INIT = 16'hbbbf;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(n41), .I3(\neo_pixel_transmitter.done_N_524 ), 
            .O(n60211));   // verilog/neopixel.v(34[12] 116[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 sub_67_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[7]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i50125_2_lut_3_lut (.I0(bit_ctr_c[3]), .I1(n43356), .I2(n69327), 
            .I3(GND_net), .O(n65478));
    defparam i50125_2_lut_3_lut.LUT_INIT = 16'h6060;
    SB_LUT4 i51982_3_lut_4_lut (.I0(bit_ctr_c[3]), .I1(n43356), .I2(n69273), 
            .I3(n67521), .O(n67668));
    defparam i51982_3_lut_4_lut.LUT_INIT = 16'hf960;
    SB_LUT4 sub_67_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[8]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[9]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[10]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i50335_2_lut_3_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(one_wire_N_479[10]), 
            .I3(n115), .O(n65449));   // verilog/neopixel.v(34[12] 116[6])
    defparam i50335_2_lut_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i2101_2_lut_3_lut_4_lut (.I0(bit_ctr_c[2]), .I1(bit_ctr[1]), 
            .I2(bit_ctr[0]), .I3(bit_ctr_c[3]), .O(n137[3]));   // verilog/neopixel.v(68[23:32])
    defparam i2101_2_lut_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 sub_67_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[0]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_67_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13[2]));   // verilog/neopixel.v(101[14:24])
    defparam sub_67_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 color_bit_N_502_1__bdd_4_lut (.I0(color_bit_N_502[1]), .I1(n62864), 
            .I2(n62865), .I3(color_bit_N_502[2]), .O(n69324));
    defparam color_bit_N_502_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n69324_bdd_4_lut (.I0(n69324), .I1(n62853), .I2(n62852), .I3(color_bit_N_502[2]), 
            .O(n69327));
    defparam n69324_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1815 (.I0(\neo_pixel_transmitter.done ), .I1(one_wire_N_479[10]), 
            .I2(n115), .I3(GND_net), .O(n40745));   // verilog/neopixel.v(34[12] 116[6])
    defparam i1_2_lut_3_lut_adj_1815.LUT_INIT = 16'h4040;
    SB_LUT4 i42402_2_lut (.I0(n58002), .I1(n58018), .I2(GND_net), .I3(GND_net), 
            .O(n58040));
    defparam i42402_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i71_4_lut (.I0(n41), .I1(n58040), .I2(\neo_pixel_transmitter.done ), 
            .I3(state[1]), .O(n48));
    defparam i71_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i1_4_lut_adj_1816 (.I0(n112), .I1(\neo_pixel_transmitter.done_N_524 ), 
            .I2(n58002), .I3(state[0]), .O(n54_adj_5657));
    defparam i1_4_lut_adj_1816.LUT_INIT = 16'h5d55;
    SB_LUT4 i1_4_lut_adj_1817 (.I0(state[0]), .I1(n54_adj_5657), .I2(n48), 
            .I3(n58018), .O(n27677));
    defparam i1_4_lut_adj_1817.LUT_INIT = 16'h50dc;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(\neo_pixel_transmitter.done_N_524 ));   // verilog/neopixel.v(34[12] 116[6])
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut (.I0(n65449), .I1(n57931), .I2(\neo_pixel_transmitter.done ), 
            .I3(n51273), .O(n29173));   // verilog/neopixel.v(34[12] 116[6])
    defparam i14_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i51835_3_lut (.I0(n69165), .I1(n69495), .I2(color_bit_N_502[2]), 
            .I3(GND_net), .O(n67521));
    defparam i51835_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28732_4_lut (.I0(n65478), .I1(n57801), .I2(n67668), .I3(n51740), 
            .O(state_1__N_440[0]));   // verilog/neopixel.v(39[18] 44[12])
    defparam i28732_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 color_bit_N_502_1__bdd_4_lut_53608 (.I0(color_bit_N_502[1]), .I1(n62795), 
            .I2(n62796), .I3(color_bit_N_502[2]), .O(n69270));
    defparam color_bit_N_502_1__bdd_4_lut_53608.LUT_INIT = 16'he4aa;
    SB_LUT4 n69270_bdd_4_lut (.I0(n69270), .I1(n62793), .I2(n62792), .I3(color_bit_N_502[2]), 
            .O(n69273));
    defparam n69270_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 state_1__I_0_102_Mux_0_i1_4_lut (.I0(n25491), .I1(n25492), .I2(state[0]), 
            .I3(bit_ctr[0]), .O(n1));   // verilog/neopixel.v(35[4] 115[11])
    defparam state_1__I_0_102_Mux_0_i1_4_lut.LUT_INIT = 16'hca35;
    SB_LUT4 n69492_bdd_4_lut (.I0(n69492), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(color_bit_N_502[1]), .O(n69495));
    defparam n69492_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i52_3_lut (.I0(bit_ctr_c[2]), .I1(bit_ctr_c[3]), .I2(bit_ctr[1]), 
            .I3(GND_net), .O(n41_adj_5658));
    defparam i52_3_lut.LUT_INIT = 16'h2424;
    SB_LUT4 i3_4_lut (.I0(n51740), .I1(n41_adj_5658), .I2(bit_ctr[1]), 
            .I3(bit_ctr[0]), .O(n23));
    defparam i3_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i42173_2_lut (.I0(n23), .I1(n43462), .I2(GND_net), .I3(GND_net), 
            .O(n57801));
    defparam i42173_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2089_2_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6897));   // verilog/neopixel.v(68[23:32])
    defparam i2089_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15161_2_lut (.I0(n27920), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n29169));   // verilog/neopixel.v(34[12] 116[6])
    defparam i15161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n69162_bdd_4_lut_4_lut (.I0(color_bit_N_502[1]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(n69162), .O(n69165));   // verilog/neopixel.v(18[6:15])
    defparam n69162_bdd_4_lut_4_lut.LUT_INIT = 16'hf588;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1)_U0 
//

module \quadrature_decoder(1)_U0  (b_prev, GND_net, a_new, position_31__N_3827, 
            ENCODER0_B_N_keep, n1779, ENCODER0_A_N_keep, n29724, n1742, 
            n1744, \encoder0_position[30] , \encoder0_position[29] , \encoder0_position[28] , 
            \encoder0_position[27] , \encoder0_position[26] , \encoder0_position[25] , 
            \encoder0_position[24] , \encoder0_position[23] , \encoder0_position[22] , 
            \encoder0_position[21] , \encoder0_position[20] , \encoder0_position[19] , 
            \encoder0_position[18] , \encoder0_position[17] , \encoder0_position[16] , 
            \encoder0_position[15] , \encoder0_position[14] , \encoder0_position[13] , 
            \encoder0_position[12] , \encoder0_position[11] , \encoder0_position[10] , 
            \encoder0_position[9] , \encoder0_position[8] , \encoder0_position[7] , 
            \encoder0_position[6] , \encoder0_position[5] , \encoder0_position[4] , 
            \encoder0_position[3] , \encoder0_position[2] , \encoder0_position[1] , 
            \encoder0_position[0] , VCC_net) /* synthesis lattice_noprune=1 */ ;
    output b_prev;
    input GND_net;
    output [1:0]a_new;
    output position_31__N_3827;
    input ENCODER0_B_N_keep;
    input n1779;
    input ENCODER0_A_N_keep;
    input n29724;
    output n1742;
    output n1744;
    output \encoder0_position[30] ;
    output \encoder0_position[29] ;
    output \encoder0_position[28] ;
    output \encoder0_position[27] ;
    output \encoder0_position[26] ;
    output \encoder0_position[25] ;
    output \encoder0_position[24] ;
    output \encoder0_position[23] ;
    output \encoder0_position[22] ;
    output \encoder0_position[21] ;
    output \encoder0_position[20] ;
    output \encoder0_position[19] ;
    output \encoder0_position[18] ;
    output \encoder0_position[17] ;
    output \encoder0_position[16] ;
    output \encoder0_position[15] ;
    output \encoder0_position[14] ;
    output \encoder0_position[13] ;
    output \encoder0_position[12] ;
    output \encoder0_position[11] ;
    output \encoder0_position[10] ;
    output \encoder0_position[9] ;
    output \encoder0_position[8] ;
    output \encoder0_position[7] ;
    output \encoder0_position[6] ;
    output \encoder0_position[5] ;
    output \encoder0_position[4] ;
    output \encoder0_position[3] ;
    output \encoder0_position[2] ;
    output \encoder0_position[1] ;
    output \encoder0_position[0] ;
    input VCC_net;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire position_31__N_3830, debounce_cnt, a_prev, direction_N_3832;
    wire [1:0]a_new_c;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire a_prev_N_3835, n29751, n29750;
    wire [31:0]n133;
    
    wire n50590, n50589, n50588, n50587, n50586, n50585, n50584, 
        n50583, n50582, n50581, n50580, n50579, n50578, n50577, 
        n50576, n50575, n50574, n50573, n50572, n50571, n50570, 
        n50569, n50568, n50567, n50566, n50565, n50564, n50563, 
        n50562, n50561, n50560;
    
    SB_LUT4 b_prev_I_0_43_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(position_31__N_3830));   // vhdl/quadrature_decoder.vhd(63[37:56])
    defparam b_prev_I_0_43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(position_31__N_3830), 
            .I3(a_new[1]), .O(position_31__N_3827));   // vhdl/quadrature_decoder.vhd(62[7] 63[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 b_prev_I_0_45_2_lut (.I0(b_prev), .I1(a_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3832));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_45_2_lut.LUT_INIT = 16'h9999;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1779), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new_c[0]), .C(n1779), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 i52690_4_lut (.I0(a_new_c[0]), .I1(b_new[0]), .I2(a_new[1]), 
            .I3(b_new[1]), .O(a_prev_N_3835));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i52690_4_lut.LUT_INIT = 16'h8421;
    SB_DFF debounce_cnt_37 (.Q(debounce_cnt), .C(n1779), .D(a_prev_N_3835));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_prev_38 (.Q(a_prev), .C(n1779), .D(n29751));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_39 (.Q(b_prev), .C(n1779), .D(n29750));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_40 (.Q(n1742), .C(n1779), .D(n29724));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_1956_add_4_33_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1744), .I3(n50590), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_1956_add_4_32_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[30] ), .I3(n50589), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_32 (.CI(n50589), .I0(direction_N_3832), 
            .I1(\encoder0_position[30] ), .CO(n50590));
    SB_LUT4 position_1956_add_4_31_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[29] ), .I3(n50588), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_31 (.CI(n50588), .I0(direction_N_3832), 
            .I1(\encoder0_position[29] ), .CO(n50589));
    SB_LUT4 position_1956_add_4_30_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[28] ), .I3(n50587), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_30 (.CI(n50587), .I0(direction_N_3832), 
            .I1(\encoder0_position[28] ), .CO(n50588));
    SB_LUT4 position_1956_add_4_29_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[27] ), .I3(n50586), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_29 (.CI(n50586), .I0(direction_N_3832), 
            .I1(\encoder0_position[27] ), .CO(n50587));
    SB_LUT4 position_1956_add_4_28_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[26] ), .I3(n50585), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_28 (.CI(n50585), .I0(direction_N_3832), 
            .I1(\encoder0_position[26] ), .CO(n50586));
    SB_LUT4 position_1956_add_4_27_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[25] ), .I3(n50584), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_27 (.CI(n50584), .I0(direction_N_3832), 
            .I1(\encoder0_position[25] ), .CO(n50585));
    SB_LUT4 position_1956_add_4_26_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[24] ), .I3(n50583), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_26 (.CI(n50583), .I0(direction_N_3832), 
            .I1(\encoder0_position[24] ), .CO(n50584));
    SB_LUT4 position_1956_add_4_25_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[23] ), .I3(n50582), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_25 (.CI(n50582), .I0(direction_N_3832), 
            .I1(\encoder0_position[23] ), .CO(n50583));
    SB_LUT4 position_1956_add_4_24_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[22] ), .I3(n50581), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_24 (.CI(n50581), .I0(direction_N_3832), 
            .I1(\encoder0_position[22] ), .CO(n50582));
    SB_LUT4 position_1956_add_4_23_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[21] ), .I3(n50580), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_23 (.CI(n50580), .I0(direction_N_3832), 
            .I1(\encoder0_position[21] ), .CO(n50581));
    SB_LUT4 position_1956_add_4_22_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[20] ), .I3(n50579), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_22 (.CI(n50579), .I0(direction_N_3832), 
            .I1(\encoder0_position[20] ), .CO(n50580));
    SB_LUT4 position_1956_add_4_21_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[19] ), .I3(n50578), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_21 (.CI(n50578), .I0(direction_N_3832), 
            .I1(\encoder0_position[19] ), .CO(n50579));
    SB_LUT4 position_1956_add_4_20_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[18] ), .I3(n50577), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_20 (.CI(n50577), .I0(direction_N_3832), 
            .I1(\encoder0_position[18] ), .CO(n50578));
    SB_LUT4 position_1956_add_4_19_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[17] ), .I3(n50576), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_19 (.CI(n50576), .I0(direction_N_3832), 
            .I1(\encoder0_position[17] ), .CO(n50577));
    SB_LUT4 position_1956_add_4_18_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[16] ), .I3(n50575), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_18 (.CI(n50575), .I0(direction_N_3832), 
            .I1(\encoder0_position[16] ), .CO(n50576));
    SB_LUT4 position_1956_add_4_17_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[15] ), .I3(n50574), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_17 (.CI(n50574), .I0(direction_N_3832), 
            .I1(\encoder0_position[15] ), .CO(n50575));
    SB_LUT4 position_1956_add_4_16_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[14] ), .I3(n50573), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_16 (.CI(n50573), .I0(direction_N_3832), 
            .I1(\encoder0_position[14] ), .CO(n50574));
    SB_LUT4 position_1956_add_4_15_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[13] ), .I3(n50572), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_15 (.CI(n50572), .I0(direction_N_3832), 
            .I1(\encoder0_position[13] ), .CO(n50573));
    SB_LUT4 position_1956_add_4_14_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[12] ), .I3(n50571), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_14 (.CI(n50571), .I0(direction_N_3832), 
            .I1(\encoder0_position[12] ), .CO(n50572));
    SB_LUT4 position_1956_add_4_13_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[11] ), .I3(n50570), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_13 (.CI(n50570), .I0(direction_N_3832), 
            .I1(\encoder0_position[11] ), .CO(n50571));
    SB_LUT4 position_1956_add_4_12_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[10] ), .I3(n50569), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_12 (.CI(n50569), .I0(direction_N_3832), 
            .I1(\encoder0_position[10] ), .CO(n50570));
    SB_LUT4 position_1956_add_4_11_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[9] ), .I3(n50568), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_11 (.CI(n50568), .I0(direction_N_3832), 
            .I1(\encoder0_position[9] ), .CO(n50569));
    SB_LUT4 position_1956_add_4_10_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[8] ), .I3(n50567), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_10 (.CI(n50567), .I0(direction_N_3832), 
            .I1(\encoder0_position[8] ), .CO(n50568));
    SB_LUT4 position_1956_add_4_9_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[7] ), .I3(n50566), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_9 (.CI(n50566), .I0(direction_N_3832), 
            .I1(\encoder0_position[7] ), .CO(n50567));
    SB_LUT4 position_1956_add_4_8_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[6] ), .I3(n50565), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_8 (.CI(n50565), .I0(direction_N_3832), 
            .I1(\encoder0_position[6] ), .CO(n50566));
    SB_LUT4 position_1956_add_4_7_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[5] ), .I3(n50564), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_7 (.CI(n50564), .I0(direction_N_3832), 
            .I1(\encoder0_position[5] ), .CO(n50565));
    SB_LUT4 position_1956_add_4_6_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[4] ), .I3(n50563), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFE position_1956__i31 (.Q(n1744), .C(n1779), .E(position_31__N_3827), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_CARRY position_1956_add_4_6 (.CI(n50563), .I0(direction_N_3832), 
            .I1(\encoder0_position[4] ), .CO(n50564));
    SB_LUT4 position_1956_add_4_5_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[3] ), .I3(n50562), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_5 (.CI(n50562), .I0(direction_N_3832), 
            .I1(\encoder0_position[3] ), .CO(n50563));
    SB_LUT4 position_1956_add_4_4_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[2] ), .I3(n50561), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_4 (.CI(n50561), .I0(direction_N_3832), 
            .I1(\encoder0_position[2] ), .CO(n50562));
    SB_LUT4 position_1956_add_4_3_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder0_position[1] ), .I3(n50560), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_3 (.CI(n50560), .I0(direction_N_3832), 
            .I1(\encoder0_position[1] ), .CO(n50561));
    SB_LUT4 position_1956_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\encoder0_position[0] ), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1956_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1956_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\encoder0_position[0] ), 
            .CO(n50560));
    SB_DFFE position_1956__i30 (.Q(\encoder0_position[30] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i29 (.Q(\encoder0_position[29] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i28 (.Q(\encoder0_position[28] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i27 (.Q(\encoder0_position[27] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i26 (.Q(\encoder0_position[26] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i25 (.Q(\encoder0_position[25] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i24 (.Q(\encoder0_position[24] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i23 (.Q(\encoder0_position[23] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i22 (.Q(\encoder0_position[22] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i21 (.Q(\encoder0_position[21] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i20 (.Q(\encoder0_position[20] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i19 (.Q(\encoder0_position[19] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i18 (.Q(\encoder0_position[18] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i17 (.Q(\encoder0_position[17] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i16 (.Q(\encoder0_position[16] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i15 (.Q(\encoder0_position[15] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i14 (.Q(\encoder0_position[14] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i13 (.Q(\encoder0_position[13] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i12 (.Q(\encoder0_position[12] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i11 (.Q(\encoder0_position[11] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i10 (.Q(\encoder0_position[10] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i9 (.Q(\encoder0_position[9] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i8 (.Q(\encoder0_position[8] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i7 (.Q(\encoder0_position[7] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i6 (.Q(\encoder0_position[6] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i5 (.Q(\encoder0_position[5] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i4 (.Q(\encoder0_position[4] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i3 (.Q(\encoder0_position[3] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i2 (.Q(\encoder0_position[2] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i1 (.Q(\encoder0_position[1] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1956__i0 (.Q(\encoder0_position[0] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF a_new_i1 (.Q(a_new[1]), .C(n1779), .D(a_new_c[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1779), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 i15743_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3835), .I2(a_new[1]), 
            .I3(a_prev), .O(n29751));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15743_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15742_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3835), .I2(b_new[1]), 
            .I3(b_prev), .O(n29750));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15742_3_lut_4_lut.LUT_INIT = 16'hf780;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, clk16MHz, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk16MHz;
    input VCC_net;
    output clk32MHz;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(clk16MHz), .PLLOUTCORE(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=38 */ ;   // verilog/TinyFPGA_B.v(34[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, control_update, duty, clk16MHz, reset, 
            \PID_CONTROLLER.integral , PWMLimit, n361, IntegralLimit, 
            n155, \PID_CONTROLLER.integral_23__N_3715[0] , \Kp[7] , \Kp[8] , 
            \Kp[9] , \Kp[1] , \Kp[10] , \Kp[0] , \Kp[2] , \Kp[3] , 
            n20194, n6, n36723, \Ki[4] , \Kp[4] , \Ki[0] , \Kp[5] , 
            \Ki[2] , \PID_CONTROLLER.integral_23__N_3715[20] , n20222, 
            \Kp[11] , n212, n213, \PID_CONTROLLER.integral_23__N_3715[22] , 
            \PID_CONTROLLER.integral_23__N_3715[21] , \Ki[1] , \PID_CONTROLLER.integral_23__N_3715[23] , 
            n36694, \Ki[5] , \Kp[12] , \Ki[3] , \Kp[13] , n6_adj_31, 
            \Kp[6] , \Kp[14] , \Kp[15] , deadband, \PID_CONTROLLER.integral_23__N_3715[13] , 
            \PID_CONTROLLER.integral_23__N_3715[12] , \Ki[6] , \Ki[7] , 
            \Ki[8] , \Ki[9] , \Ki[10] , \Ki[11] , n219, \PID_CONTROLLER.integral_23__N_3715[11] , 
            \Ki[12] , n53, \PID_CONTROLLER.integral_23__N_3715[10] , \Ki[13] , 
            n4, \PID_CONTROLLER.integral_23__N_3715[9] , n11610, n27692, 
            \Ki[14] , \PID_CONTROLLER.integral_23__N_3715[8] , setpoint, 
            \motor_state[23] , \motor_state[22] , \motor_state[21] , \Ki[15] , 
            \PID_CONTROLLER.integral_23__N_3715[7] , n38, n110, \PID_CONTROLLER.integral_23__N_3715[14] , 
            \motor_state[20] , \motor_state[19] , n490, n417, n20149, 
            n344, n20150, n271, \PID_CONTROLLER.integral_23__N_3715[6] , 
            n29641, n20151, n198, VCC_net, n56, n125, n30463, 
            n30462, n30461, n30460, n30459, n30458, n30457, n30456, 
            n30455, n30454, n30453, n30452, n30451, n30450, n30449, 
            n30448, n30447, n30445, n30443, n30442, n30441, n30440, 
            n30439, \motor_state[18] , \PID_CONTROLLER.integral_23__N_3715[5] , 
            n455, n456, \motor_state[17] , n20, \motor_state[15] , 
            \motor_state[14] , \motor_state[13] , \motor_state[12] , n1, 
            \motor_state[10] , \motor_state[9] , \motor_state[8] , n401, 
            n43, \motor_state[7] , n41622, \motor_state[5] , \motor_state[4] , 
            n42235, \motor_state[2] , \motor_state[1] , \motor_state[0] , 
            n375, n376, \PID_CONTROLLER.integral_23__N_3715[4] , \PID_CONTROLLER.integral_23__N_3715[3] , 
            \PID_CONTROLLER.integral_23__N_3715[15] , \PID_CONTROLLER.integral_23__N_3715[16] , 
            \PID_CONTROLLER.integral_23__N_3715[2] , \PID_CONTROLLER.integral_23__N_3715[1] , 
            n214, n131, n204, n4_adj_32, n20195, n43349, n37189, 
            n4_adj_33, n30, n32, n4_adj_34, n20196) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output control_update;
    output [23:0]duty;
    input clk16MHz;
    input reset;
    output [23:0]\PID_CONTROLLER.integral ;
    input [23:0]PWMLimit;
    output n361;
    input [23:0]IntegralLimit;
    output n155;
    output \PID_CONTROLLER.integral_23__N_3715[0] ;
    input \Kp[7] ;
    input \Kp[8] ;
    input \Kp[9] ;
    input \Kp[1] ;
    input \Kp[10] ;
    input \Kp[0] ;
    input \Kp[2] ;
    input \Kp[3] ;
    input n20194;
    input n6;
    input n36723;
    input \Ki[4] ;
    input \Kp[4] ;
    input \Ki[0] ;
    input \Kp[5] ;
    input \Ki[2] ;
    output \PID_CONTROLLER.integral_23__N_3715[20] ;
    output n20222;
    input \Kp[11] ;
    output n212;
    output n213;
    output \PID_CONTROLLER.integral_23__N_3715[22] ;
    output \PID_CONTROLLER.integral_23__N_3715[21] ;
    input \Ki[1] ;
    output \PID_CONTROLLER.integral_23__N_3715[23] ;
    input n36694;
    input \Ki[5] ;
    input \Kp[12] ;
    input \Ki[3] ;
    input \Kp[13] ;
    input n6_adj_31;
    input \Kp[6] ;
    input \Kp[14] ;
    input \Kp[15] ;
    input [23:0]deadband;
    output \PID_CONTROLLER.integral_23__N_3715[13] ;
    input \PID_CONTROLLER.integral_23__N_3715[12] ;
    input \Ki[6] ;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Ki[9] ;
    input \Ki[10] ;
    input \Ki[11] ;
    output n219;
    output \PID_CONTROLLER.integral_23__N_3715[11] ;
    input \Ki[12] ;
    input n53;
    output \PID_CONTROLLER.integral_23__N_3715[10] ;
    input \Ki[13] ;
    input n4;
    output \PID_CONTROLLER.integral_23__N_3715[9] ;
    output n11610;
    input n27692;
    input \Ki[14] ;
    output \PID_CONTROLLER.integral_23__N_3715[8] ;
    input [23:0]setpoint;
    input \motor_state[23] ;
    input \motor_state[22] ;
    input \motor_state[21] ;
    input \Ki[15] ;
    output \PID_CONTROLLER.integral_23__N_3715[7] ;
    input n38;
    input n110;
    output \PID_CONTROLLER.integral_23__N_3715[14] ;
    input \motor_state[20] ;
    input \motor_state[19] ;
    input n490;
    input n417;
    input n20149;
    input n344;
    input n20150;
    input n271;
    output \PID_CONTROLLER.integral_23__N_3715[6] ;
    input n29641;
    input n20151;
    input n198;
    input VCC_net;
    input n56;
    input n125;
    input n30463;
    input n30462;
    input n30461;
    input n30460;
    input n30459;
    input n30458;
    input n30457;
    input n30456;
    input n30455;
    input n30454;
    input n30453;
    input n30452;
    input n30451;
    input n30450;
    input n30449;
    input n30448;
    input n30447;
    input n30445;
    input n30443;
    input n30442;
    input n30441;
    input n30440;
    input n30439;
    input \motor_state[18] ;
    output \PID_CONTROLLER.integral_23__N_3715[5] ;
    output n455;
    output n456;
    input \motor_state[17] ;
    input n20;
    input \motor_state[15] ;
    input \motor_state[14] ;
    input \motor_state[13] ;
    input \motor_state[12] ;
    input n1;
    input \motor_state[10] ;
    input \motor_state[9] ;
    input \motor_state[8] ;
    output n401;
    output n43;
    input \motor_state[7] ;
    input n41622;
    input \motor_state[5] ;
    input \motor_state[4] ;
    input n42235;
    input \motor_state[2] ;
    input \motor_state[1] ;
    input \motor_state[0] ;
    output n375;
    output n376;
    output \PID_CONTROLLER.integral_23__N_3715[4] ;
    output \PID_CONTROLLER.integral_23__N_3715[3] ;
    output \PID_CONTROLLER.integral_23__N_3715[15] ;
    output \PID_CONTROLLER.integral_23__N_3715[16] ;
    output \PID_CONTROLLER.integral_23__N_3715[2] ;
    output \PID_CONTROLLER.integral_23__N_3715[1] ;
    output n214;
    input n131;
    input n204;
    output n4_adj_32;
    output n20195;
    output n43349;
    input n37189;
    input n4_adj_33;
    output n30;
    input n32;
    input n4_adj_34;
    output n20196;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [43:0]n257;
    wire [47:0]n49;
    
    wire n49241;
    wire [23:0]n352;
    wire [23:0]n432;
    
    wire n45, n43_c;
    wire [23:0]n51;
    wire [23:0]n130;
    wire [23:0]n55;
    
    wire n49240;
    wire [23:0]n57;
    
    wire n37, n23, n25;
    wire [23:0]n182;
    
    wire n6_c, n68212, n39, n68136, n43_adj_5119, n41, n68111, 
        n66419, n67615, n67291, n45_adj_5120, n66415, n67920, n65576, 
        n66577, n29, n31, n35, n33, n68121, n181;
    wire [23:0]n207;
    
    wire n9, n533, n606, n679, n80, n752, n11, n153, n226;
    wire [4:0]n20146;
    
    wire n299, n372_adj_5122;
    wire [1:0]n20229;
    
    wire n49059, n17, n19, n825, n62;
    wire [16:0]n16376;
    wire [15:0]n16987;
    
    wire n49597, n61832, n61836, n898, n61834, n971, n49008, n61842, 
        n4_c, n8, n59684, n49596, n49239, n1114, n49595, n1041, 
        n49594, n968, n49593, n21_adj_5124, n11_adj_5125, counter_31__N_3714, 
        n895, n49592, n13, n445_adj_5126, n15, n49238, n518, n822, 
        n49591, n27, n66219, n749, n49590, n49237, n591, n66211, 
        n12, n664, n676, n49589, n737, n49236, n101, n32_c, 
        n603, n49588, n810, n530, n49587, n457, n49586, n384, 
        n49585, n10, n1044, n1117, n311, n49584, n30_c, n49235, 
        n238, n49583, n165, n49582, n174, n883, n23_adj_5128, 
        n92, n956, n49234, n49233, n1029, n247, n1102, n66229, 
        n67099, n49232, n320, n66382, n125_c, n49231, n66398, 
        n56_c;
    wire [14:0]n17530;
    
    wire n49569, n49568, n49567, n49230, n49566, n198_c, n67661, 
        n11608, n49565, n393, n886, n66260, n66266, n271_c, n48904, 
        n61894, n67095, n68033, n344_c;
    wire [2:0]n20198;
    
    wire n4_adj_5131;
    wire [4:0]n20100;
    
    wire n49564, n466, n539, n417_c, n347, n6_adj_5132, n57286, 
        n959, n49563, n49562, n49229, n49561, n61890, n49560, 
        n49228, n62_adj_5133, n48918, n60074, n490_c, n61880, n69804, 
        n61884, n8_adj_5134, n6_adj_5135, n59192, n41_adj_5136, n1032, 
        n183_adj_5137, n256, n329, n402;
    wire [0:0]n12226;
    wire [21:0]n12733;
    
    wire n50874, n475, n67493, n460, n49559, n548, n621, n694, 
        n767, n840, n68148, n107_adj_5139, n50873, n50872, n387, 
        n49558, n50871, n50870, n50869, n314, n49557, n50868;
    wire [0:0]n11650;
    wire [21:0]n12109;
    
    wire n49831, n50867, n1096, n50866, n1023, n50865, n950, n50864, 
        n241, n49556, n168, n49555, n877, n50863, n49830, n26, 
        n95, n180, n804, n50862, n731, n50861, n658, n50860, 
        n253, n6_adj_5141, n67656, n612, n49829, n585, n50859, 
        n49828, n512, n50858;
    wire [6:0]n19984;
    wire [5:0]n20078;
    
    wire n560, n49554, n487, n49553, n49827, n326, n49826, n399, 
        n414, n49552, n49825, n16_adj_5142, n49824, n1096_adj_5143, 
        n49823, n1023_adj_5144, n49822, n950_adj_5145, n49821, n472, 
        n439_adj_5147, n50857, n545, n618, n691, n764, n877_adj_5148, 
        n49820, n341_adj_5149, n49551, n366_adj_5150, n50856, n293, 
        n50855, n268, n49550, n804_adj_5151, n49819, n220, n50854, 
        n837, n910, n731_adj_5153, n49818, n122_adj_5154, n53_c, 
        n195, n147, n50853, n658_adj_5155, n49817, n585_adj_5157, 
        n49816, n49227, n195_adj_5158, n49549, n5, n74, n512_adj_5159, 
        n49815, n8_adj_5160;
    wire [20:0]n13698;
    
    wire n50852, n24, n268_adj_5161, n50851, n341_adj_5162, n50850, 
        n67657, n414_adj_5163, n50849, n50848, n50847, n50846, n122_adj_5165, 
        n1099, n50845, n1026, n50844, n685, n66185, n953, n50843, 
        n439_adj_5166, n49814, n880, n50842, n487_adj_5167, n560_adj_5168, 
        n807, n50841, n734, n50840, n661, n50839, n588, n50838, 
        n104, n35_adj_5171, n66183, n67299, n177, n250, n323, 
        n515, n50837, n396, n366_adj_5172, n49813, n469, n542, 
        n66606, n615, n688, n442_adj_5173, n50836, n293_adj_5174, 
        n49812, n761, n369_adj_5175, n50835, n296_adj_5176, n50834, 
        n834, n907, n980, n223, n50833, n67654, n150, n50832, 
        n8_adj_5178, n77;
    wire [19:0]n14576;
    
    wire n50831, n50830, n50829, n1105, n50828, n67655, n101_adj_5179, 
        n32_adj_5180, n174_adj_5181, n49226, n50827, n66205, n50826, 
        n247_adj_5182, n320_adj_5183, n758, n1102_adj_5184, n50825, 
        n1029_adj_5185, n50824, n956_adj_5186, n50823, n883_adj_5187, 
        n50822, n810_adj_5188, n50821, n737_adj_5189, n50820, n664_adj_5190, 
        n50819, n591_adj_5191, n50818, n220_adj_5192, n49811, n147_adj_5194, 
        n49810, n65738, n518_adj_5195, n50817, n5_adj_5196, n74_adj_5197, 
        n445_adj_5198, n50816, n372_adj_5199, n50815, n299_adj_5200, 
        n50814, n226_adj_5201, n50813, n153_adj_5202, n50812, n66203, 
        n68071, n49225, n11_adj_5203, n80_adj_5204;
    wire [10:0]n19102;
    wire [9:0]n19365;
    
    wire n840_adj_5205, n50811, n767_adj_5206, n50810;
    wire [13:0]n18009;
    
    wire n1120, n49537, n694_adj_5207, n50809, n1047, n49536, n621_adj_5208, 
        n50808, n548_adj_5209, n50807, n974, n49535, n475_adj_5210, 
        n50806, n402_adj_5211, n50805, n329_adj_5212, n50804, n256_adj_5213, 
        n50803, n183_adj_5215, n50802, n393_adj_5216, n41_adj_5217, 
        n110_adj_5218, n466_adj_5219, n49224;
    wire [18:0]n15372;
    
    wire n50801, n50800, n831, n50799, n50798, n50797, n1105_adj_5221, 
        n50796, n1032_adj_5222, n50795, n959_adj_5223, n50794, n886_adj_5224, 
        n50793, n813, n50792, n740, n50791, n66608, n68247, n68248, 
        n39_adj_5225, n68202, n41_adj_5226, n66187, n67928, n66614, 
        n68125, n68126, n405, n60219, n667, n50790, n594, n50789, 
        n539_adj_5227, n521, n50788, n448_adj_5228, n50787, n375_c, 
        n50786, n302, n50785, n229, n50784, n156, n50783;
    wire [9:0]n19506;
    wire [8:0]n19702;
    
    wire n770, n49791, n49223, n14_adj_5229, n83;
    wire [17:0]n16090;
    
    wire n50782, n50781, n50780, n50779, n612_adj_5230, n904, n1108, 
        n50778, n1035, n50777, n962, n50776, n889, n50775, n697, 
        n49790, n816, n50774, n743, n50773, n624, n49789, n670, 
        n50772, n597, n50771, n524, n50770, n451_adj_5231, n50769, 
        n378, n50768, n305, n50767, n232, n50766, n159, n50765, 
        n17_adj_5232, n86;
    wire [8:0]n19584;
    
    wire n770_adj_5233, n50764, n551, n49788, n697_adj_5234, n50763, 
        n901, n49534, n624_adj_5235, n50762, n478, n49787, n551_adj_5236, 
        n50761, n478_adj_5237, n50760, n6_adj_5238, n977, n685_adj_5239, 
        n405_adj_5240, n50759, n332_adj_5241, n50758, n259, n50757, 
        n186_adj_5242, n50756, n44, n113_adj_5243;
    wire [16:0]n16734;
    
    wire n50755, n50754, n50753, n828, n49533, n1111, n50752, 
        n1038, n50751, n965, n50750, n49222, n892, n50749, n819, 
        n50748, n746, n50747, n673, n50746, n600, n50745, n527, 
        n50744, n454, n50743, n381, n50742, n308, n50741, n235, 
        n50740, n162, n50739, n20_adj_5244, n89;
    wire [15:0]n17308;
    
    wire n50738, n50737, n1114_adj_5245, n50736, n1041_adj_5246, n50735, 
        n968_adj_5247, n50734, n895_adj_5248, n50733, n822_adj_5249, 
        n50732, n749_adj_5250, n50731, n405_adj_5251, n49786, n676_adj_5252, 
        n50730, n603_adj_5253, n50729, n77_adj_5254, n755, n49532, 
        n530_adj_5255, n50728, n682, n49531, n457_adj_5256, n50727, 
        n384_adj_5257, n50726, n311_adj_5258, n50725, n238_adj_5259, 
        n50724, n332_adj_5260, n49785, n165_adj_5261, n50723, n609, 
        n49530, n49221, n23_adj_5263, n92_adj_5264, n8_adj_5265;
    wire [7:0]n19763;
    
    wire n700, n50722, n536, n49529, n627, n50721, n259_adj_5266, 
        n49784, n463, n49528, n554, n50720, n758_adj_5267, n481, 
        n50719, n408, n50718, n335_adj_5268, n50717, n390, n49527, 
        n262, n50716, n186_adj_5269, n49783, n189, n50715, n831_adj_5270, 
        n47, n116_adj_5271, n317, n49526;
    wire [14:0]n17816;
    
    wire n50714, n1117_adj_5272, n50713, n1044_adj_5273, n50712, n971_adj_5274, 
        n50711, n150_adj_5275, n898_adj_5276, n50710, n825_adj_5277, 
        n50709, n752_adj_5278, n50708, n679_adj_5279, n50707, n44_adj_5280, 
        n113_adj_5281, n606_adj_5283, n50706, n244, n49525, n533_adj_5284, 
        n50705, n904_adj_5285, n171, n49524, n460_adj_5286, n50704, 
        n1050, n387_adj_5287, n50703, n314_adj_5288, n50702, n241_adj_5289, 
        n50701;
    wire [20:0]n13171;
    
    wire n49782, n977_adj_5290, n29_adj_5291, n98, n49220, n49781, 
        n168_adj_5292, n50700, n49379, n49780, n26_adj_5293, n95_adj_5294, 
        n1050_adj_5296, n49378, n119_adj_5298;
    wire [13:0]n18262;
    
    wire n1120_adj_5299, n50699, n50, n1047_adj_5300, n50698, n223_adj_5301, 
        n974_adj_5302, n50697, n49779, n49778, n901_adj_5303, n50696, 
        n49777, n828_adj_5304, n50695, n755_adj_5305, n50694, n49377, 
        n49776, n682_adj_5307, n50693, n49376, n296_adj_5309, n192, 
        n1099_adj_5310, n49775, n609_adj_5311, n50692, n265, n49375, 
        n1026_adj_5313, n49774, n953_adj_5314, n49773, n49374, n536_adj_5315, 
        n50691, n880_adj_5317, n49772, n338_adj_5318, n807_adj_5319, 
        n49771, n463_adj_5320, n50690, n369_adj_5321, n442_adj_5322, 
        n734_adj_5323, n49770, n661_adj_5324, n49769, n390_adj_5325, 
        n50689, n317_adj_5326, n50688, n244_adj_5327, n50687, n411, 
        n484, n515_adj_5328, n557, n588_adj_5329, n49768, n171_adj_5330, 
        n50686, n630, n49373, n29_adj_5332, n98_adj_5333;
    wire [6:0]n19906;
    
    wire n50685, n50684, n49767, n50683, n50682, n49766, n49765, 
        n50681, n49372, n50680, n49219, n50679, n49764, n49763, 
        n49371;
    wire [12:0]n18650;
    
    wire n50678, n49370, n50677;
    wire [12:0]n18428;
    
    wire n49513, n49218, n50676, n49762, n50675, n41_adj_5335, n50674, 
        n50673, n49512, n49511, n50672, n50671, n49510, n50670, 
        n50669, n49369, n49217, n49509, n50668, n50667, n39_adj_5336, 
        n50666, n49216;
    wire [11:0]n18984;
    
    wire n50665, n50664, n50663, n50662, n50661, n50660, n50659, 
        n50658, n50657, n50656, n50655, n50654, n45_adj_5337;
    wire [5:0]n20017;
    
    wire n50653, n50652, n49215, n49508, n50651, n43_adj_5338, n50650, 
        n50649, n50648;
    wire [10:0]n19268;
    
    wire n50647, n50646, n50645, n50644, n50643, n50642, n50641, 
        n50640, n50639, n49507, n50638, n50637;
    wire [19:0]n14095;
    
    wire n49744, n50636, n50635, n37_adj_5341, n50634, n50633, n50632, 
        n50631, n49368, n50630, n49743, n50629, n50628, n50627, 
        n50626, n49742, n50625, n49506, n49505, n50624, n49367, 
        n50623, n49504, n49366, n23_adj_5343, n50622, n25_adj_5344, 
        n49214, n49741, n49503, n49365, n49740, n49739, n49364, 
        n35_adj_5346, n29_adj_5347, n49738, n49502, n49363, n49737, 
        n31_adj_5348, n49736, n49735, n49501, n49362, n49734, n49733, 
        n49732, n49213, n49731, n49730, n49729, n49500, n49728, 
        n49727, n33_adj_5350, n49499, n49726, n49725, n11_adj_5352, 
        n49361, n49498, n49360, n13_adj_5354, n49497, n15_adj_5356, 
        n49359, n27_adj_5357, n9_adj_5358, n17_adj_5359, n19_adj_5360, 
        n21_adj_5361, n65702, n65676, n12_adj_5362;
    wire [31:0]n59;
    wire [31:0]counter;   // verilog/motorControl.v(21[11:18])
    
    wire n50495, n50494, n50493, n50492, n50491, n50490, n50489, 
        n50488, n50487, n50486, n50485, n50484, n50483, n50482, 
        n50481, n50480, n50479, n50478, n50477, n50476, n50475, 
        n50474, n50473, n50472, n50471, n50470, n49496, n50469, 
        n10_adj_5391, n50468, n50467, n50466, n50465, n30_adj_5392, 
        n49212, n66411, n49358, n66641, n66631, n67912, n67281, 
        n68115, n16_adj_5404, n67910, n67911, n8_adj_5405, n24_adj_5406, 
        n65599, n65581, n67289, n67607, n4_adj_5407, n67859, n67860, 
        n65664, n65657, n68152, n67609, n68287, n68288, n68250, 
        n65614, n67612, n40_adj_5408, n67918;
    wire [18:0]n14934;
    
    wire n49708, n49707, n37_adj_5409, n49706, n49357, n49705, n49704, 
        n29_adj_5411, n49703, n49702, n31_adj_5412, n49701, n49700, 
        n23_adj_5413;
    wire [11:0]n18791;
    
    wire n980_adj_5414, n49486, n813_adj_5415, n49699, n907_adj_5416, 
        n49485, n47_adj_5417;
    wire [23:0]n61;
    
    wire n49356, n740_adj_5419, n49698, n667_adj_5420, n49697, n594_adj_5421, 
        n49696, n521_adj_5422, n49695;
    wire [23:0]n63;
    
    wire n49355, n834_adj_5424, n49484, n448_adj_5425, n49694, n375_adj_5426, 
        n49693, n49211, n761_adj_5427, n49483, n49354, n302_adj_5430, 
        n49692, n688_adj_5431, n49482, n229_adj_5432, n49691, n156_adj_5433, 
        n49690, n49353, n14_adj_5435, n83_adj_5436, n615_adj_5437, 
        n49481, n49352, n542_adj_5439, n49480, n469_adj_5440, n49479, 
        n396_adj_5441, n49478, n49351;
    wire [7:0]n19860;
    
    wire n700_adj_5444, n49689, n49210, n627_adj_5446, n49688, n49350, 
        n25_adj_5448, n554_adj_5449, n49687, n49209, n49208, n481_adj_5450, 
        n49686, n408_adj_5451, n49685, n49349, n335_adj_5453, n49684, 
        n262_adj_5454, n49683, n323_adj_5455, n49477, n189_adj_5456, 
        n49682, n49207, n250_adj_5457, n49476, n47_adj_5458, n116_adj_5459, 
        n49348, n49206, n177_adj_5462, n49475, n49205, n49347, n49346, 
        n35_adj_5465, n104_adj_5466, n49204, n49345, n49344, n49343, 
        n49342, n49341, n49203, n49263;
    wire [17:0]n15693;
    
    wire n49666, n49340, n49665, n49664, n49339, n49663, n49262, 
        n1108_adj_5477, n49662, n1035_adj_5478, n49661, n49338, n962_adj_5480, 
        n49660, n889_adj_5481, n49659, n49261, n816_adj_5482, n49658, 
        n49337, n49336, n743_adj_5486, n49657, n49202, n670_adj_5487, 
        n49656, n49260, n49335, n597_adj_5489, n49655, n49334, n524_adj_5491, 
        n49654, n451_adj_5492, n49653, n378_adj_5493, n49652, n49259, 
        n305_adj_5494, n49651, n232_adj_5495, n49650, n159_adj_5496, 
        n49649, n37174, n17_adj_5499, n86_adj_5500, n49258;
    wire [23:0]n65;
    
    wire n49333, n49332, n49257, n49256, n49201, n49200, n49199, 
        n49331, n49330, n49329, n49255, n49634, n49633, n49254, 
        n49198, n49632, n49328, n49327, n1111_adj_5509, n49631, 
        n1038_adj_5510, n49630, n965_adj_5511, n49629, n49197, n49253, 
        n49196, n49326, n892_adj_5513, n49628, n910_adj_5514, n49448, 
        n837_adj_5515, n49447, n49195, n49325, n49252, n764_adj_5517, 
        n49446, n819_adj_5518, n49627, n49251, n49324, n691_adj_5520, 
        n49445, n618_adj_5521, n49444, n746_adj_5522, n49626, n49250, 
        n673_adj_5523, n49625, n600_adj_5524, n49624, n545_adj_5525, 
        n49443, n49249, n49323, n472_adj_5527, n49442, n399_adj_5528, 
        n49441, n49322, n49248, n326_adj_5530, n49440, n527_adj_5531, 
        n49623, n49321, n454_adj_5533, n49622, n381_adj_5534, n49621, 
        n49247, n253_adj_5535, n49439, n308_adj_5536, n49620, n49320, 
        n180_adj_5538, n49438, n49246, n235_adj_5539, n49619, n162_adj_5540, 
        n49618, n38_adj_5541, n107_adj_5542, n20_adj_5543, n89_adj_5544, 
        n49245, n630_adj_5545, n49617, n557_adj_5546, n49616, n49319, 
        n49318, n49317, n484_adj_5550, n49615, n411_adj_5551, n49614, 
        n49244, n35_adj_5552, n33_adj_5553, n11_adj_5554, n49316, 
        n338_adj_5556, n49613, n49315, n265_adj_5558, n49612, n49243, 
        n192_adj_5559, n49611, n13_adj_5560, n15_adj_5561, n27_adj_5562, 
        n9_adj_5563, n50_adj_5564, n119_adj_5565, n17_adj_5566, n49314, 
        n49313, n49242, n19_adj_5569, n49312, n49311, n21_adj_5574, 
        n11_adj_5575, n13_adj_5576, n9_adj_5577, n17_adj_5578, n7_adj_5579, 
        n19_adj_5580, n21_adj_5581, n65530, n23_adj_5582, n15_adj_5583, 
        n25_adj_5584, n65522, n12_adj_5586, n10_adj_5587, n30_adj_5588, 
        n66454, n66448, n67867, n65513, n67219;
    wire [2:0]n20220;
    
    wire n14_adj_5590, n15_adj_5591, n8_adj_5592, n12_adj_5593, n16_adj_5594, 
        n10_adj_5595, n59568, n59846, n16_adj_5596, n15_adj_5597, 
        n17_adj_5598, n16_adj_5599, n67855, n67856, n8_adj_5600, n24_adj_5604, 
        n4_adj_5605, n67853, n67854, n27892, n65515, n68061, n27887, 
        n27882, n28_adj_5606, n27877, n68211, n27872, n27867, n27862, 
        n27857, n33_adj_5607, n31_adj_5608, n37_adj_5609, n35_adj_5610, 
        n25_adj_5611, n27_adj_5612, n29_adj_5613, n21_adj_5614, n23_adj_5615, 
        n13_adj_5616, n15_adj_5617, n17_adj_5618, n9_adj_5619, n11_adj_5620, 
        n19_adj_5621, n43_adj_5622, n27852, n41_adj_5623, n37_adj_5624, 
        n39_adj_5625, n5_adj_5626, n66268, n66264, n10_adj_5627, n27847, 
        n27842, n12_adj_5628, n8_adj_5629, n27837, n27832, n6_adj_5630, 
        n27827, n16_adj_5631, n68069, n68070, n67949, n67799, n27822, 
        n67847, n66601, n68075, n68076, n27817, n27812, n27807, 
        n27802, n67662, n67663, n27797, n27792, n66246, n67111, 
        n34_adj_5635, n67622, n66603, n67660, n66356, n67171, n69591, 
        n67159, n69585, n12_adj_5636, n66320, n69610, n10_adj_5637, 
        n30_adj_5638, n66352, n67167, n69604, n67165, n69599, n16_adj_5639, 
        n66278, n8_adj_5640, n24_adj_5641, n66361, n69630, n66358, 
        n69623, n67531, n69626, n67169, n67805, n66337, n69589, 
        n67525, n69615, n68067, n69580, n68260, n69577, n10_adj_5642, 
        n67205, n67545, n67543, n66391, n65316, n6_adj_5643, n67680, 
        n14_adj_5644, n12_adj_5645, n32_adj_5646, n66388, n67681, 
        n66384, n68063, n66581, n6_adj_5647, n67676, n67677, n67670, 
        n67671, n66322, n68065, n66591, n68245, n68246, n68208, 
        n66282, n69574, n67295, n66589, n66289, n67924, n66597, 
        n8_adj_5649, n67682, n67683, n67195, n67293, n66579, n67811, 
        n68243, n67851, n68307, n68308, n68154, n68077, n68078, 
        n68123, n61858, n27787;
    
    SB_CARRY add_18_2 (.CI(GND_net), .I0(n257[0]), .I1(n49[0]), .CO(n49241));
    SB_LUT4 LessThan_25_i45_2_lut (.I0(n352[22]), .I1(n432[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i43_2_lut (.I0(n352[21]), .I1(n432[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_c));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i43_2_lut.LUT_INIT = 16'h6666;
    SB_DFFER result__i0 (.Q(duty[0]), .C(clk16MHz), .E(control_update), 
            .D(n51[0]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_LUT4 add_9_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n55[23]), .I3(n49240), .O(n130[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[3]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_25_i37_2_lut (.I0(n352[18]), .I1(n432[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i23_2_lut (.I0(n352[11]), .I1(n432[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i25_2_lut (.I0(n352[12]), .I1(n432[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i6_3_lut_3_lut (.I0(n130[3]), .I1(n182[3]), .I2(n182[2]), 
            .I3(GND_net), .O(n6_c));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i52450_3_lut (.I0(n68212), .I1(n182[19]), .I2(n39), .I3(GND_net), 
            .O(n68136));   // verilog/motorControl.v(48[21:44])
    defparam i52450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50733_4_lut (.I0(n43_adj_5119), .I1(n41), .I2(n39), .I3(n68111), 
            .O(n66419));
    defparam i50733_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52234_4_lut (.I0(n67615), .I1(n67291), .I2(n45_adj_5120), 
            .I3(n66415), .O(n67920));   // verilog/motorControl.v(48[21:44])
    defparam i52234_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49890_3_lut_4_lut (.I0(n130[3]), .I1(n182[3]), .I2(n182[2]), 
            .I3(n130[2]), .O(n65576));   // verilog/motorControl.v(48[21:44])
    defparam i49890_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i50891_3_lut (.I0(n68136), .I1(n182[20]), .I2(n41), .I3(GND_net), 
            .O(n66577));   // verilog/motorControl.v(48[21:44])
    defparam i50891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i29_2_lut (.I0(n352[14]), .I1(n432[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i31_2_lut (.I0(n361), .I1(n432[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i35_2_lut (.I0(n352[17]), .I1(n432[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i33_2_lut (.I0(n352[16]), .I1(n432[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52435_4_lut (.I0(n66577), .I1(n67920), .I2(n45_adj_5120), 
            .I3(n66419), .O(n68121));   // verilog/motorControl.v(48[21:44])
    defparam i52435_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52436_3_lut (.I0(n68121), .I1(n130[23]), .I2(n182[23]), .I3(GND_net), 
            .O(n181));   // verilog/motorControl.v(48[21:44])
    defparam i52436_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_14_i1_3_lut (.I0(n130[0]), .I1(n182[0]), .I2(n181), .I3(GND_net), 
            .O(n207[0]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i1_3_lut (.I0(n207[0]), .I1(IntegralLimit[0]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[0] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_25_i9_2_lut (.I0(n352[4]), .I1(n432[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i359_2_lut (.I0(\Kp[7] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i408_2_lut (.I0(\Kp[8] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[4]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_26_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[5]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i457_2_lut (.I0(\Kp[9] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n679));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i55_2_lut (.I0(\Kp[1] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n80));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i506_2_lut (.I0(\Kp[10] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i8_2_lut (.I0(\Kp[0] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i104_2_lut (.I0(\Kp[2] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n153));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i153_2_lut (.I0(\Kp[3] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n226));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(n20194), .I1(n6), .I2(n36723), .I3(\Ki[4] ), 
            .O(n20146[3]));   // verilog/motorControl.v(51[27:38])
    defparam i1_4_lut.LUT_INIT = 16'h9666;
    SB_LUT4 mult_16_i202_2_lut (.I0(\Kp[4] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n299));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n49[0]));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i251_2_lut (.I0(\Kp[5] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_5122));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1789 (.I0(n20229[0]), .I1(n49059), .I2(\Ki[2] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3715[20] ), .O(n20222));   // verilog/motorControl.v(51[27:38])
    defparam i1_4_lut_adj_1789.LUT_INIT = 16'h9666;
    SB_LUT4 LessThan_25_i17_2_lut (.I0(n352[8]), .I1(n432[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i19_2_lut (.I0(n352[9]), .I1(n432[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i555_2_lut (.I0(\Kp[11] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i42_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i21_3_lut (.I0(n130[20]), .I1(n182[20]), .I2(n181), 
            .I3(GND_net), .O(n207[20]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i21_3_lut (.I0(n207[20]), .I1(IntegralLimit[20]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[20] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i20_3_lut (.I0(n130[19]), .I1(n182[19]), .I2(n181), 
            .I3(GND_net), .O(n212));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i19_3_lut (.I0(n130[18]), .I1(n182[18]), .I2(n181), 
            .I3(GND_net), .O(n213));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i23_3_lut (.I0(n130[22]), .I1(n182[22]), .I2(n181), 
            .I3(GND_net), .O(n207[22]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6272_18_lut (.I0(GND_net), .I1(n16987[15]), .I2(GND_net), 
            .I3(n49597), .O(n16376[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i23_3_lut (.I0(n207[22]), .I1(IntegralLimit[22]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[22] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i22_3_lut (.I0(n130[21]), .I1(n182[21]), .I2(n181), 
            .I3(GND_net), .O(n207[21]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i22_3_lut (.I0(n207[21]), .I1(IntegralLimit[21]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[21] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1790 (.I0(\Ki[1] ), .I1(\Ki[0] ), .I2(\PID_CONTROLLER.integral_23__N_3715[22] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3715[23] ), .O(n61832));   // verilog/motorControl.v(51[27:38])
    defparam i1_4_lut_adj_1790.LUT_INIT = 16'h93a0;
    SB_LUT4 i1_4_lut_adj_1791 (.I0(n36723), .I1(n36694), .I2(\Ki[5] ), 
            .I3(\Ki[4] ), .O(n61836));   // verilog/motorControl.v(51[27:38])
    defparam i1_4_lut_adj_1791.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_16_i604_2_lut (.I0(\Kp[12] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1792 (.I0(\Ki[3] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3715[20] ), 
            .I3(\PID_CONTROLLER.integral_23__N_3715[21] ), .O(n61834));   // verilog/motorControl.v(51[27:38])
    defparam i1_4_lut_adj_1792.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_16_i653_2_lut (.I0(\Kp[13] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1793 (.I0(n61834), .I1(n49008), .I2(n61836), 
            .I3(n61832), .O(n61842));   // verilog/motorControl.v(51[27:38])
    defparam i1_4_lut_adj_1793.LUT_INIT = 16'h6996;
    SB_LUT4 i35183_4_lut (.I0(n20229[0]), .I1(\Ki[2] ), .I2(n49059), .I3(\PID_CONTROLLER.integral_23__N_3715[20] ), 
            .O(n4_c));   // verilog/motorControl.v(51[27:38])
    defparam i35183_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i35015_4_lut (.I0(n20194), .I1(n36723), .I2(n6), .I3(\Ki[4] ), 
            .O(n8));   // verilog/motorControl.v(51[27:38])
    defparam i35015_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_1794 (.I0(n6_adj_31), .I1(n8), .I2(n4_c), .I3(n61842), 
            .O(n59684));   // verilog/motorControl.v(51[27:38])
    defparam i1_4_lut_adj_1794.LUT_INIT = 16'h6996;
    SB_LUT4 add_6272_17_lut (.I0(GND_net), .I1(n16987[14]), .I2(GND_net), 
            .I3(n49596), .O(n16376[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_17 (.CI(n49596), .I0(n16987[14]), .I1(GND_net), 
            .CO(n49597));
    SB_LUT4 add_9_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n55[23]), .I3(n49239), .O(n130[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6272_16_lut (.I0(GND_net), .I1(n16987[13]), .I2(n1114), 
            .I3(n49595), .O(n16376[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i2_2_lut (.I0(\Kp[0] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n257[0]));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i2_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6272_16 (.CI(n49595), .I0(n16987[13]), .I1(n1114), .CO(n49596));
    SB_LUT4 add_6272_15_lut (.I0(GND_net), .I1(n16987[12]), .I2(n1041), 
            .I3(n49594), .O(n16376[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_15 (.CI(n49594), .I0(n16987[12]), .I1(n1041), .CO(n49595));
    SB_LUT4 add_6272_14_lut (.I0(GND_net), .I1(n16987[11]), .I2(n968), 
            .I3(n49593), .O(n16376[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_14 (.CI(n49593), .I0(n16987[11]), .I1(n968), .CO(n49594));
    SB_LUT4 LessThan_25_i21_2_lut (.I0(n352[10]), .I1(n432[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5124));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i11_2_lut (.I0(n352[5]), .I1(n432[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5125));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i11_2_lut.LUT_INIT = 16'h6666;
    SB_DFF control_update_37 (.Q(control_update), .C(clk16MHz), .D(counter_31__N_3714));   // verilog/motorControl.v(23[10] 30[6])
    SB_LUT4 add_6272_13_lut (.I0(GND_net), .I1(n16987[10]), .I2(n895), 
            .I3(n49592), .O(n16376[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_13 (.CI(n49592), .I0(n16987[10]), .I1(n895), .CO(n49593));
    SB_LUT4 LessThan_25_i13_2_lut (.I0(n352[6]), .I1(n432[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_9_24 (.CI(n49239), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n55[23]), .CO(n49240));
    SB_LUT4 mult_16_i300_2_lut (.I0(\Kp[6] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_5126));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_25_i15_2_lut (.I0(n352[7]), .I1(n432[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_9_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n55[23]), .I3(n49238), .O(n130[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i349_2_lut (.I0(\Kp[7] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6272_12_lut (.I0(GND_net), .I1(n16987[9]), .I2(n822), 
            .I3(n49591), .O(n16376[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_23 (.CI(n49238), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n55[23]), .CO(n49239));
    SB_LUT4 LessThan_25_i27_2_lut (.I0(n352[13]), .I1(n432[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i27_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6272_12 (.CI(n49591), .I0(n16987[9]), .I1(n822), .CO(n49592));
    SB_LUT4 i50533_4_lut (.I0(n21_adj_5124), .I1(n19), .I2(n17), .I3(n9), 
            .O(n66219));
    defparam i50533_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_6272_11_lut (.I0(GND_net), .I1(n16987[8]), .I2(n749), 
            .I3(n49590), .O(n16376[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n55[23]), .I3(n49237), .O(n130[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i398_2_lut (.I0(\Kp[8] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50525_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11_adj_5125), 
            .O(n66211));
    defparam i50525_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_6272_11 (.CI(n49590), .I0(n16987[8]), .I1(n749), .CO(n49591));
    SB_LUT4 LessThan_25_i12_3_lut (.I0(n432[7]), .I1(n432[16]), .I2(n33), 
            .I3(GND_net), .O(n12));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i447_2_lut (.I0(\Kp[9] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i447_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_9_22 (.CI(n49237), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n55[23]), .CO(n49238));
    SB_LUT4 add_6272_10_lut (.I0(GND_net), .I1(n16987[7]), .I2(n676), 
            .I3(n49589), .O(n16376[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_10 (.CI(n49589), .I0(n16987[7]), .I1(n676), .CO(n49590));
    SB_LUT4 mult_16_i496_2_lut (.I0(\Kp[10] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n55[23]), .I3(n49236), .O(n130[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_21 (.CI(n49236), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n55[23]), .CO(n49237));
    SB_LUT4 mult_16_i69_2_lut (.I0(\Kp[1] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i22_2_lut (.I0(\Kp[0] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n32_c));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6272_9_lut (.I0(GND_net), .I1(n16987[6]), .I2(n603), .I3(n49588), 
            .O(n16376[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_9 (.CI(n49588), .I0(n16987[6]), .I1(n603), .CO(n49589));
    SB_LUT4 mult_16_i545_2_lut (.I0(\Kp[11] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6272_8_lut (.I0(GND_net), .I1(n16987[5]), .I2(n530), .I3(n49587), 
            .O(n16376[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_8 (.CI(n49587), .I0(n16987[5]), .I1(n530), .CO(n49588));
    SB_LUT4 add_6272_7_lut (.I0(GND_net), .I1(n16987[4]), .I2(n457), .I3(n49586), 
            .O(n16376[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_7 (.CI(n49586), .I0(n16987[4]), .I1(n457), .CO(n49587));
    SB_LUT4 add_6272_6_lut (.I0(GND_net), .I1(n16987[3]), .I2(n384), .I3(n49585), 
            .O(n16376[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_25_i10_3_lut (.I0(n432[5]), .I1(n432[6]), .I2(n13), 
            .I3(GND_net), .O(n10));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i702_2_lut (.I0(\Kp[14] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i702_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6272_6 (.CI(n49585), .I0(n16987[3]), .I1(n384), .CO(n49586));
    SB_LUT4 mult_16_i751_2_lut (.I0(\Kp[15] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6272_5_lut (.I0(GND_net), .I1(n16987[2]), .I2(n311), .I3(n49584), 
            .O(n16376[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_25_i30_3_lut (.I0(n12), .I1(n432[17]), .I2(n35), 
            .I3(GND_net), .O(n30_c));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6272_5 (.CI(n49584), .I0(n16987[2]), .I1(n311), .CO(n49585));
    SB_LUT4 add_9_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n55[22]), .I3(n49235), .O(n130[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_20 (.CI(n49235), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n55[22]), .CO(n49236));
    SB_LUT4 unary_minus_26_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[6]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6272_4_lut (.I0(GND_net), .I1(n16987[1]), .I2(n238), .I3(n49583), 
            .O(n16376[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6272_4 (.CI(n49583), .I0(n16987[1]), .I1(n238), .CO(n49584));
    SB_LUT4 add_6272_3_lut (.I0(GND_net), .I1(n16987[0]), .I2(n165), .I3(n49582), 
            .O(n16376[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i118_2_lut (.I0(\Kp[2] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i594_2_lut (.I0(\Kp[12] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i594_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6272_3 (.CI(n49582), .I0(n16987[0]), .I1(n165), .CO(n49583));
    SB_LUT4 add_6272_2_lut (.I0(GND_net), .I1(n23_adj_5128), .I2(n92), 
            .I3(GND_net), .O(n16376[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6272_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i643_2_lut (.I0(\Kp[13] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i643_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6272_2 (.CI(GND_net), .I0(n23_adj_5128), .I1(n92), .CO(n49582));
    SB_LUT4 add_9_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n55[21]), .I3(n49234), .O(n130[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_19 (.CI(n49234), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n55[21]), .CO(n49235));
    SB_LUT4 add_9_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n55[20]), .I3(n49233), .O(n130[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i692_2_lut (.I0(\Kp[14] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[7]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i167_2_lut (.I0(\Kp[3] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n247));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i741_2_lut (.I0(\Kp[15] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[8]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51413_4_lut (.I0(n13), .I1(n11_adj_5125), .I2(n9), .I3(n66229), 
            .O(n67099));
    defparam i51413_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_9_18 (.CI(n49233), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n55[20]), .CO(n49234));
    SB_LUT4 add_9_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n55[19]), .I3(n49232), .O(n130[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[9]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i216_2_lut (.I0(\Kp[4] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n320));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50696_2_lut_4_lut (.I0(deadband[17]), .I1(n352[17]), .I2(deadband[8]), 
            .I3(n352[8]), .O(n66382));
    defparam i50696_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_9_17 (.CI(n49232), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n55[19]), .CO(n49233));
    SB_LUT4 mult_16_i85_2_lut (.I0(\Kp[1] ), .I1(n55[21]), .I2(GND_net), 
            .I3(GND_net), .O(n125_c));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n55[18]), .I3(n49231), .O(n130[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_16 (.CI(n49231), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n55[18]), .CO(n49232));
    SB_LUT4 i50712_2_lut_4_lut (.I0(deadband[9]), .I1(n352[9]), .I2(deadband[5]), 
            .I3(n352[5]), .O(n66398));
    defparam i50712_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i38_2_lut (.I0(\Kp[0] ), .I1(n55[22]), .I2(GND_net), 
            .I3(GND_net), .O(n56_c));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6305_17_lut (.I0(GND_net), .I1(n17530[14]), .I2(GND_net), 
            .I3(n49569), .O(n16987[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6305_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6305_16_lut (.I0(GND_net), .I1(n17530[13]), .I2(n1117), 
            .I3(n49568), .O(n16987[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6305_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6305_16 (.CI(n49568), .I0(n17530[13]), .I1(n1117), .CO(n49569));
    SB_LUT4 add_6305_15_lut (.I0(GND_net), .I1(n17530[12]), .I2(n1044), 
            .I3(n49567), .O(n16987[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6305_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6305_15 (.CI(n49567), .I0(n17530[12]), .I1(n1044), .CO(n49568));
    SB_LUT4 add_9_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n55[17]), .I3(n49230), .O(n130[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6305_14_lut (.I0(GND_net), .I1(n17530[11]), .I2(n971), 
            .I3(n49566), .O(n16987[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6305_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6305_14 (.CI(n49566), .I0(n17530[11]), .I1(n971), .CO(n49567));
    SB_LUT4 mult_16_i134_2_lut (.I0(\Kp[2] ), .I1(n55[21]), .I2(GND_net), 
            .I3(GND_net), .O(n198_c));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5967_2_lut_4_lut (.I0(control_update), .I1(n67661), .I2(PWMLimit[23]), 
            .I3(n352[23]), .O(n11608));
    defparam i5967_2_lut_4_lut.LUT_INIT = 16'h2a02;
    SB_LUT4 unary_minus_26_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[10]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6305_13_lut (.I0(GND_net), .I1(n17530[10]), .I2(n898), 
            .I3(n49565), .O(n16987[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6305_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i265_2_lut (.I0(\Kp[5] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i596_2_lut (.I0(\Kp[12] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50574_2_lut_4_lut (.I0(PWMLimit[8]), .I1(n352[8]), .I2(PWMLimit[4]), 
            .I3(n352[4]), .O(n66260));
    defparam i50574_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i50580_2_lut_4_lut (.I0(PWMLimit[6]), .I1(n352[6]), .I2(PWMLimit[5]), 
            .I3(n352[5]), .O(n66266));
    defparam i50580_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i183_2_lut (.I0(\Kp[3] ), .I1(n55[21]), .I2(GND_net), 
            .I3(GND_net), .O(n271_c));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1795 (.I0(n55[23]), .I1(\Kp[2] ), .I2(n48904), 
            .I3(n55[22]), .O(n61894));   // verilog/motorControl.v(51[18:24])
    defparam i1_4_lut_adj_1795.LUT_INIT = 16'h6ca0;
    SB_LUT4 unary_minus_26_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[11]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51409_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n67099), 
            .O(n67095));
    defparam i51409_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52347_4_lut (.I0(n25), .I1(n23), .I2(n21_adj_5124), .I3(n67095), 
            .O(n68033));
    defparam i52347_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_16_i232_2_lut (.I0(\Kp[4] ), .I1(n55[21]), .I2(GND_net), 
            .I3(GND_net), .O(n344_c));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1796 (.I0(n55[22]), .I1(n20198[1]), .I2(n4_adj_5131), 
            .I3(\Kp[3] ), .O(n20100[2]));   // verilog/motorControl.v(51[18:24])
    defparam i1_4_lut_adj_1796.LUT_INIT = 16'hc66c;
    SB_CARRY add_6305_13 (.CI(n49565), .I0(n17530[10]), .I1(n898), .CO(n49566));
    SB_LUT4 add_6305_12_lut (.I0(GND_net), .I1(n17530[9]), .I2(n825), 
            .I3(n49564), .O(n16987[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6305_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i314_2_lut (.I0(\Kp[6] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n466));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i363_2_lut (.I0(\Kp[7] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n539));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i281_2_lut (.I0(\Kp[5] ), .I1(n55[21]), .I2(GND_net), 
            .I3(GND_net), .O(n417_c));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i234_2_lut (.I0(\Kp[4] ), .I1(n55[22]), .I2(GND_net), 
            .I3(GND_net), .O(n347));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i234_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1797 (.I0(n20198[1]), .I1(n6_adj_5132), .I2(n347), 
            .I3(n57286), .O(n20100[3]));   // verilog/motorControl.v(51[18:24])
    defparam i1_4_lut_adj_1797.LUT_INIT = 16'h6996;
    SB_LUT4 mult_16_i645_2_lut (.I0(\Kp[13] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i645_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6305_12 (.CI(n49564), .I0(n17530[9]), .I1(n825), .CO(n49565));
    SB_LUT4 add_6305_11_lut (.I0(GND_net), .I1(n17530[8]), .I2(n752), 
            .I3(n49563), .O(n16987[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6305_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6305_11 (.CI(n49563), .I0(n17530[8]), .I1(n752), .CO(n49564));
    SB_LUT4 add_6305_10_lut (.I0(GND_net), .I1(n17530[7]), .I2(n679), 
            .I3(n49562), .O(n16987[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6305_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_15 (.CI(n49230), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n55[17]), .CO(n49231));
    SB_LUT4 add_9_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n55[16]), .I3(n49229), .O(n130[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6305_10 (.CI(n49562), .I0(n17530[7]), .I1(n679), .CO(n49563));
    SB_LUT4 i35041_2_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n48904));   // verilog/motorControl.v(51[18:24])
    defparam i35041_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6305_9_lut (.I0(GND_net), .I1(n17530[6]), .I2(n606), .I3(n49561), 
            .O(n16987[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6305_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut (.I0(n61890), .I1(n55[23]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_5131));   // verilog/motorControl.v(51[18:24])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35102_4_lut (.I0(n20198[1]), .I1(\Kp[3] ), .I2(n4_adj_5131), 
            .I3(n55[22]), .O(n6_adj_5132));   // verilog/motorControl.v(51[18:24])
    defparam i35102_4_lut.LUT_INIT = 16'he800;
    SB_CARRY add_6305_9 (.CI(n49561), .I0(n17530[6]), .I1(n606), .CO(n49562));
    SB_CARRY add_9_14 (.CI(n49229), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n55[16]), .CO(n49230));
    SB_LUT4 i1_3_lut (.I0(\Kp[0] ), .I1(\Kp[2] ), .I2(\Kp[1] ), .I3(GND_net), 
            .O(n61890));   // verilog/motorControl.v(51[18:24])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 add_6305_8_lut (.I0(GND_net), .I1(n17530[5]), .I2(n533), .I3(n49560), 
            .O(n16987[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6305_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n55[15]), .I3(n49228), .O(n130[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i40_2_lut (.I0(\Kp[0] ), .I1(n55[23]), .I2(GND_net), 
            .I3(GND_net), .O(n62_adj_5133));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i40_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46701_3_lut (.I0(n55[23]), .I1(n61890), .I2(\Kp[3] ), .I3(GND_net), 
            .O(n57286));   // verilog/motorControl.v(51[18:24])
    defparam i46701_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 i35233_3_lut (.I0(n55[23]), .I1(n48918), .I2(n60074), .I3(GND_net), 
            .O(n20198[1]));   // verilog/motorControl.v(51[18:24])
    defparam i35233_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_16_i330_2_lut (.I0(\Kp[6] ), .I1(n55[21]), .I2(GND_net), 
            .I3(GND_net), .O(n490_c));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1798 (.I0(n55[23]), .I1(\Kp[5] ), .I2(n60074), 
            .I3(n55[22]), .O(n61880));   // verilog/motorControl.v(51[18:24])
    defparam i1_4_lut_adj_1798.LUT_INIT = 16'hc60a;
    SB_CARRY add_6305_8 (.CI(n49560), .I0(n17530[5]), .I1(n533), .CO(n49561));
    SB_LUT4 i1_rep_294_2_lut (.I0(n20198[1]), .I1(n57286), .I2(GND_net), 
            .I3(GND_net), .O(n69804));   // verilog/motorControl.v(51[18:24])
    defparam i1_rep_294_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1799 (.I0(n48918), .I1(n61880), .I2(\Kp[4] ), 
            .I3(n55[23]), .O(n61884));   // verilog/motorControl.v(51[18:24])
    defparam i1_4_lut_adj_1799.LUT_INIT = 16'h9666;
    SB_LUT4 i35110_4_lut (.I0(n69804), .I1(\Kp[4] ), .I2(n6_adj_5132), 
            .I3(n55[22]), .O(n8_adj_5134));   // verilog/motorControl.v(51[18:24])
    defparam i35110_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i35063_4_lut (.I0(n20198[1]), .I1(\Kp[3] ), .I2(n61890), .I3(n55[23]), 
            .O(n6_adj_5135));   // verilog/motorControl.v(51[18:24])
    defparam i35063_4_lut.LUT_INIT = 16'he800;
    SB_LUT4 i1_4_lut_adj_1800 (.I0(n6_adj_5135), .I1(n8_adj_5134), .I2(n61884), 
            .I3(n57286), .O(n59192));   // verilog/motorControl.v(51[18:24])
    defparam i1_4_lut_adj_1800.LUT_INIT = 16'h6996;
    SB_LUT4 mult_17_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5136));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i694_2_lut (.I0(\Kp[14] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_5137));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n256));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3715[23] ), 
            .I1(n12733[21]), .I2(GND_net), .I3(n50874), .O(n12226[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_26_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[12]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51807_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n68033), 
            .O(n67493));
    defparam i51807_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 add_6305_7_lut (.I0(GND_net), .I1(n17530[4]), .I2(n460), .I3(n49559), 
            .O(n16987[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6305_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n621));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n694));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n767));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i13_3_lut (.I0(n130[12]), .I1(n182[12]), .I2(n181), 
            .I3(GND_net), .O(n219));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52462_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n67493), 
            .O(n68148));
    defparam i52462_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_17_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_5139));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i73_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6305_7 (.CI(n49559), .I0(n17530[4]), .I1(n460), .CO(n49560));
    SB_LUT4 mult_17_add_1225_23_lut (.I0(GND_net), .I1(n12733[20]), .I2(GND_net), 
            .I3(n50873), .O(n49[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_23 (.CI(n50873), .I0(n12733[20]), .I1(GND_net), 
            .CO(n50874));
    SB_LUT4 mult_17_add_1225_22_lut (.I0(GND_net), .I1(n12733[19]), .I2(GND_net), 
            .I3(n50872), .O(n49[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6305_6_lut (.I0(GND_net), .I1(n17530[3]), .I2(n387), .I3(n49558), 
            .O(n16987[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6305_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_22 (.CI(n50872), .I0(n12733[19]), .I1(GND_net), 
            .CO(n50873));
    SB_LUT4 mult_17_add_1225_21_lut (.I0(GND_net), .I1(n12733[18]), .I2(GND_net), 
            .I3(n50871), .O(n49[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_21 (.CI(n50871), .I0(n12733[18]), .I1(GND_net), 
            .CO(n50872));
    SB_LUT4 mult_17_add_1225_20_lut (.I0(GND_net), .I1(n12733[17]), .I2(GND_net), 
            .I3(n50870), .O(n49[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_20 (.CI(n50870), .I0(n12733[17]), .I1(GND_net), 
            .CO(n50871));
    SB_LUT4 mult_17_add_1225_19_lut (.I0(GND_net), .I1(n12733[16]), .I2(GND_net), 
            .I3(n50869), .O(n49[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6305_6 (.CI(n49558), .I0(n17530[3]), .I1(n387), .CO(n49559));
    SB_LUT4 add_6305_5_lut (.I0(GND_net), .I1(n17530[2]), .I2(n314), .I3(n49557), 
            .O(n16987[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6305_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_19 (.CI(n50869), .I0(n12733[16]), .I1(GND_net), 
            .CO(n50870));
    SB_LUT4 mult_17_add_1225_18_lut (.I0(GND_net), .I1(n12733[15]), .I2(GND_net), 
            .I3(n50868), .O(n49[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_18 (.CI(n50868), .I0(n12733[15]), .I1(GND_net), 
            .CO(n50869));
    SB_LUT4 mult_16_add_1221_24_lut (.I0(n55[23]), .I1(n12109[21]), .I2(GND_net), 
            .I3(n49831), .O(n11650[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_17_add_1225_17_lut (.I0(GND_net), .I1(n12733[14]), .I2(GND_net), 
            .I3(n50867), .O(n49[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_17 (.CI(n50867), .I0(n12733[14]), .I1(GND_net), 
            .CO(n50868));
    SB_LUT4 mult_17_add_1225_16_lut (.I0(GND_net), .I1(n12733[13]), .I2(n1096), 
            .I3(n50866), .O(n49[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_16 (.CI(n50866), .I0(n12733[13]), .I1(n1096), 
            .CO(n50867));
    SB_CARRY add_6305_5 (.CI(n49557), .I0(n17530[2]), .I1(n314), .CO(n49558));
    SB_LUT4 mult_17_add_1225_15_lut (.I0(GND_net), .I1(n12733[12]), .I2(n1023), 
            .I3(n50865), .O(n49[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_15 (.CI(n50865), .I0(n12733[12]), .I1(n1023), 
            .CO(n50866));
    SB_LUT4 mult_17_add_1225_14_lut (.I0(GND_net), .I1(n12733[11]), .I2(n950), 
            .I3(n50864), .O(n49[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6305_4_lut (.I0(GND_net), .I1(n17530[1]), .I2(n241), .I3(n49556), 
            .O(n16987[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6305_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6305_4 (.CI(n49556), .I0(n17530[1]), .I1(n241), .CO(n49557));
    SB_CARRY mult_17_add_1225_14 (.CI(n50864), .I0(n12733[11]), .I1(n950), 
            .CO(n50865));
    SB_LUT4 add_6305_3_lut (.I0(GND_net), .I1(n17530[0]), .I2(n168), .I3(n49555), 
            .O(n16987[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6305_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_13_lut (.I0(GND_net), .I1(n12733[10]), .I2(n877), 
            .I3(n50863), .O(n49[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_13 (.CI(n50863), .I0(n12733[10]), .I1(n877), 
            .CO(n50864));
    SB_LUT4 mult_16_add_1221_23_lut (.I0(GND_net), .I1(n12109[20]), .I2(GND_net), 
            .I3(n49830), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6305_3 (.CI(n49555), .I0(n17530[0]), .I1(n168), .CO(n49556));
    SB_LUT4 add_6305_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n16987[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6305_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1225_12_lut (.I0(GND_net), .I1(n12733[9]), .I2(n804), 
            .I3(n50862), .O(n49[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_12 (.CI(n50862), .I0(n12733[9]), .I1(n804), 
            .CO(n50863));
    SB_LUT4 mult_17_add_1225_11_lut (.I0(GND_net), .I1(n12733[8]), .I2(n731), 
            .I3(n50861), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_11 (.CI(n50861), .I0(n12733[8]), .I1(n731), 
            .CO(n50862));
    SB_LUT4 mult_17_add_1225_10_lut (.I0(GND_net), .I1(n12733[7]), .I2(n658), 
            .I3(n50860), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6305_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n49555));
    SB_LUT4 mult_17_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51970_3_lut (.I0(n6_adj_5141), .I1(n432[10]), .I2(n21_adj_5124), 
            .I3(GND_net), .O(n67656));   // verilog/motorControl.v(55[23:39])
    defparam i51970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i412_2_lut (.I0(\Kp[8] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n612));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i412_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_17_add_1225_10 (.CI(n50860), .I0(n12733[7]), .I1(n658), 
            .CO(n50861));
    SB_CARRY mult_16_add_1221_23 (.CI(n49830), .I0(n12109[20]), .I1(GND_net), 
            .CO(n49831));
    SB_LUT4 mult_16_add_1221_22_lut (.I0(GND_net), .I1(n12109[19]), .I2(GND_net), 
            .I3(n49829), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_22 (.CI(n49829), .I0(n12109[19]), .I1(GND_net), 
            .CO(n49830));
    SB_LUT4 mult_17_add_1225_9_lut (.I0(GND_net), .I1(n12733[6]), .I2(n585), 
            .I3(n50859), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1221_21_lut (.I0(GND_net), .I1(n12109[18]), .I2(GND_net), 
            .I3(n49828), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_21 (.CI(n49828), .I0(n12109[18]), .I1(GND_net), 
            .CO(n49829));
    SB_CARRY mult_17_add_1225_9 (.CI(n50859), .I0(n12733[6]), .I1(n585), 
            .CO(n50860));
    SB_LUT4 mult_17_add_1225_8_lut (.I0(GND_net), .I1(n12733[5]), .I2(n512), 
            .I3(n50858), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6521_8_lut (.I0(GND_net), .I1(n20078[5]), .I2(n560), .I3(n49554), 
            .O(n19984[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6521_7_lut (.I0(GND_net), .I1(n20078[4]), .I2(n487), .I3(n49553), 
            .O(n19984[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_7 (.CI(n49553), .I0(n20078[4]), .I1(n487), .CO(n49554));
    SB_LUT4 mult_16_add_1221_20_lut (.I0(GND_net), .I1(n12109[17]), .I2(GND_net), 
            .I3(n49827), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i220_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1221_20 (.CI(n49827), .I0(n12109[17]), .I1(GND_net), 
            .CO(n49828));
    SB_LUT4 mult_16_add_1221_19_lut (.I0(GND_net), .I1(n12109[16]), .I2(GND_net), 
            .I3(n49826), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6521_6_lut (.I0(GND_net), .I1(n20078[3]), .I2(n414), .I3(n49552), 
            .O(n19984[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_19 (.CI(n49826), .I0(n12109[16]), .I1(GND_net), 
            .CO(n49827));
    SB_LUT4 mult_16_add_1221_18_lut (.I0(GND_net), .I1(n12109[15]), .I2(GND_net), 
            .I3(n49825), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_18 (.CI(n49825), .I0(n12109[15]), .I1(GND_net), 
            .CO(n49826));
    SB_LUT4 LessThan_25_i16_3_lut (.I0(n432[9]), .I1(n432[21]), .I2(n43_c), 
            .I3(GND_net), .O(n16_adj_5142));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_add_1221_17_lut (.I0(GND_net), .I1(n12109[14]), .I2(GND_net), 
            .I3(n49824), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_17 (.CI(n49824), .I0(n12109[14]), .I1(GND_net), 
            .CO(n49825));
    SB_CARRY mult_17_add_1225_8 (.CI(n50858), .I0(n12733[5]), .I1(n512), 
            .CO(n50859));
    SB_LUT4 mult_16_add_1221_16_lut (.I0(GND_net), .I1(n12109[13]), .I2(n1096_adj_5143), 
            .I3(n49823), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_16 (.CI(n49823), .I0(n12109[13]), .I1(n1096_adj_5143), 
            .CO(n49824));
    SB_LUT4 mult_16_add_1221_15_lut (.I0(GND_net), .I1(n12109[12]), .I2(n1023_adj_5144), 
            .I3(n49822), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_15 (.CI(n49822), .I0(n12109[12]), .I1(n1023_adj_5144), 
            .CO(n49823));
    SB_LUT4 mult_16_add_1221_14_lut (.I0(GND_net), .I1(n12109[11]), .I2(n950_adj_5145), 
            .I3(n49821), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_6 (.CI(n49552), .I0(n20078[3]), .I1(n414), .CO(n49553));
    SB_LUT4 mult_17_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_add_1225_7_lut (.I0(GND_net), .I1(n12733[4]), .I2(n439_adj_5147), 
            .I3(n50857), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i367_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1221_14 (.CI(n49821), .I0(n12109[11]), .I1(n950_adj_5145), 
            .CO(n49822));
    SB_CARRY mult_17_add_1225_7 (.CI(n50857), .I0(n12733[4]), .I1(n439_adj_5147), 
            .CO(n50858));
    SB_LUT4 mult_17_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_add_1221_13_lut (.I0(GND_net), .I1(n12109[10]), .I2(n877_adj_5148), 
            .I3(n49820), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6521_5_lut (.I0(GND_net), .I1(n20078[2]), .I2(n341_adj_5149), 
            .I3(n49551), .O(n19984[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_add_1225_6_lut (.I0(GND_net), .I1(n12733[3]), .I2(n366_adj_5150), 
            .I3(n50856), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_6 (.CI(n50856), .I0(n12733[3]), .I1(n366_adj_5150), 
            .CO(n50857));
    SB_LUT4 mult_17_add_1225_5_lut (.I0(GND_net), .I1(n12733[2]), .I2(n293), 
            .I3(n50855), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_5 (.CI(n49551), .I0(n20078[2]), .I1(n341_adj_5149), 
            .CO(n49552));
    SB_LUT4 add_6521_4_lut (.I0(GND_net), .I1(n20078[1]), .I2(n268), .I3(n49550), 
            .O(n19984[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_13 (.CI(n49820), .I0(n12109[10]), .I1(n877_adj_5148), 
            .CO(n49821));
    SB_CARRY add_6521_4 (.CI(n49550), .I0(n20078[1]), .I1(n268), .CO(n49551));
    SB_LUT4 mult_16_add_1221_12_lut (.I0(GND_net), .I1(n12109[9]), .I2(n804_adj_5151), 
            .I3(n49819), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_17_add_1225_5 (.CI(n50855), .I0(n12733[2]), .I1(n293), 
            .CO(n50856));
    SB_LUT4 mult_17_add_1225_4_lut (.I0(GND_net), .I1(n12733[1]), .I2(n220), 
            .I3(n50854), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_12 (.CI(n49819), .I0(n12109[9]), .I1(n804_adj_5151), 
            .CO(n49820));
    SB_CARRY mult_17_add_1225_4 (.CI(n50854), .I0(n12733[1]), .I1(n220), 
            .CO(n50855));
    SB_LUT4 mult_17_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_add_1221_11_lut (.I0(GND_net), .I1(n12109[8]), .I2(n731_adj_5153), 
            .I3(n49818), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i83_2_lut (.I0(\Kp[1] ), .I1(n55[20]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_5154));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i36_2_lut (.I0(\Kp[0] ), .I1(n55[21]), .I2(GND_net), 
            .I3(GND_net), .O(n53_c));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i132_2_lut (.I0(\Kp[2] ), .I1(n55[20]), .I2(GND_net), 
            .I3(GND_net), .O(n195));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i132_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1221_11 (.CI(n49818), .I0(n12109[8]), .I1(n731_adj_5153), 
            .CO(n49819));
    SB_LUT4 mult_17_add_1225_3_lut (.I0(GND_net), .I1(n12733[0]), .I2(n147), 
            .I3(n50853), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1221_10_lut (.I0(GND_net), .I1(n12109[7]), .I2(n658_adj_5155), 
            .I3(n49817), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_10 (.CI(n49817), .I0(n12109[7]), .I1(n658_adj_5155), 
            .CO(n49818));
    SB_LUT4 mult_16_add_1221_9_lut (.I0(GND_net), .I1(n12109[6]), .I2(n585_adj_5157), 
            .I3(n49816), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_13 (.CI(n49228), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n55[15]), .CO(n49229));
    SB_CARRY mult_16_add_1221_9 (.CI(n49816), .I0(n12109[6]), .I1(n585_adj_5157), 
            .CO(n49817));
    SB_CARRY mult_17_add_1225_3 (.CI(n50853), .I0(n12733[0]), .I1(n147), 
            .CO(n50854));
    SB_LUT4 add_9_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n55[14]), .I3(n49227), .O(n130[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6521_3_lut (.I0(GND_net), .I1(n20078[0]), .I2(n195_adj_5158), 
            .I3(n49549), .O(n19984[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_12 (.CI(n49227), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n55[14]), .CO(n49228));
    SB_LUT4 mult_17_add_1225_2_lut (.I0(GND_net), .I1(n5), .I2(n74), .I3(GND_net), 
            .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_17_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1221_8_lut (.I0(GND_net), .I1(n12109[5]), .I2(n512_adj_5159), 
            .I3(n49815), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_8 (.CI(n49815), .I0(n12109[5]), .I1(n512_adj_5159), 
            .CO(n49816));
    SB_LUT4 LessThan_25_i8_3_lut (.I0(n432[4]), .I1(n432[8]), .I2(n17), 
            .I3(GND_net), .O(n8_adj_5160));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_17_add_1225_2 (.CI(GND_net), .I0(n5), .I1(n74), .CO(n50853));
    SB_LUT4 add_6100_23_lut (.I0(GND_net), .I1(n13698[20]), .I2(GND_net), 
            .I3(n50852), .O(n12733[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_25_i24_3_lut (.I0(n16_adj_5142), .I1(n432[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i181_2_lut (.I0(\Kp[3] ), .I1(n55[20]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_5161));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6100_22_lut (.I0(GND_net), .I1(n13698[19]), .I2(GND_net), 
            .I3(n50851), .O(n12733[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_22 (.CI(n50851), .I0(n13698[19]), .I1(GND_net), 
            .CO(n50852));
    SB_LUT4 mult_16_i230_2_lut (.I0(\Kp[4] ), .I1(n55[20]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_5162));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6100_21_lut (.I0(GND_net), .I1(n13698[18]), .I2(GND_net), 
            .I3(n50850), .O(n12733[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_21 (.CI(n50850), .I0(n13698[18]), .I1(GND_net), 
            .CO(n50851));
    SB_LUT4 i51971_3_lut (.I0(n67656), .I1(n432[11]), .I2(n23), .I3(GND_net), 
            .O(n67657));   // verilog/motorControl.v(55[23:39])
    defparam i51971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i279_2_lut (.I0(\Kp[5] ), .I1(n55[20]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_5163));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6100_20_lut (.I0(GND_net), .I1(n13698[17]), .I2(GND_net), 
            .I3(n50849), .O(n12733[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_20 (.CI(n50849), .I0(n13698[17]), .I1(GND_net), 
            .CO(n50850));
    SB_LUT4 add_6100_19_lut (.I0(GND_net), .I1(n13698[16]), .I2(GND_net), 
            .I3(n50848), .O(n12733[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_19 (.CI(n50848), .I0(n13698[16]), .I1(GND_net), 
            .CO(n50849));
    SB_LUT4 add_6100_18_lut (.I0(GND_net), .I1(n13698[15]), .I2(GND_net), 
            .I3(n50847), .O(n12733[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_18 (.CI(n50847), .I0(n13698[15]), .I1(GND_net), 
            .CO(n50848));
    SB_LUT4 add_6100_17_lut (.I0(GND_net), .I1(n13698[14]), .I2(GND_net), 
            .I3(n50846), .O(n12733[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_3 (.CI(n49549), .I0(n20078[0]), .I1(n195_adj_5158), 
            .CO(n49550));
    SB_LUT4 add_6521_2_lut (.I0(GND_net), .I1(n53), .I2(n122_adj_5165), 
            .I3(GND_net), .O(n19984[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_17 (.CI(n50846), .I0(n13698[14]), .I1(GND_net), 
            .CO(n50847));
    SB_LUT4 add_6100_16_lut (.I0(GND_net), .I1(n13698[13]), .I2(n1099), 
            .I3(n50845), .O(n12733[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_16 (.CI(n50845), .I0(n13698[13]), .I1(n1099), .CO(n50846));
    SB_LUT4 add_6100_15_lut (.I0(GND_net), .I1(n13698[12]), .I2(n1026), 
            .I3(n50844), .O(n12733[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i461_2_lut (.I0(\Kp[9] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i461_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6100_15 (.CI(n50844), .I0(n13698[12]), .I1(n1026), .CO(n50845));
    SB_CARRY add_6521_2 (.CI(GND_net), .I0(n53), .I1(n122_adj_5165), .CO(n49549));
    SB_LUT4 i50499_4_lut (.I0(n43_c), .I1(n25), .I2(n23), .I3(n66219), 
            .O(n66185));
    defparam i50499_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_6100_14_lut (.I0(GND_net), .I1(n13698[11]), .I2(n953), 
            .I3(n50843), .O(n12733[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_14 (.CI(n50843), .I0(n13698[11]), .I1(n953), .CO(n50844));
    SB_LUT4 mult_16_add_1221_7_lut (.I0(GND_net), .I1(n12109[4]), .I2(n439_adj_5166), 
            .I3(n49814), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6100_13_lut (.I0(GND_net), .I1(n13698[10]), .I2(n880), 
            .I3(n50842), .O(n12733[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_13 (.CI(n50842), .I0(n13698[10]), .I1(n880), .CO(n50843));
    SB_LUT4 mult_16_i328_2_lut (.I0(\Kp[6] ), .I1(n55[20]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_5167));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i377_2_lut (.I0(\Kp[7] ), .I1(n55[20]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_5168));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i377_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_16_add_1221_7 (.CI(n49814), .I0(n12109[4]), .I1(n439_adj_5166), 
            .CO(n49815));
    SB_LUT4 add_6100_12_lut (.I0(GND_net), .I1(n13698[9]), .I2(n807), 
            .I3(n50841), .O(n12733[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i12_3_lut (.I0(n130[11]), .I1(n182[11]), .I2(n181), 
            .I3(GND_net), .O(n207[11]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6100_12 (.CI(n50841), .I0(n13698[9]), .I1(n807), .CO(n50842));
    SB_LUT4 add_6100_11_lut (.I0(GND_net), .I1(n13698[8]), .I2(n734), 
            .I3(n50840), .O(n12733[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_11 (.CI(n50840), .I0(n13698[8]), .I1(n734), .CO(n50841));
    SB_LUT4 add_6100_10_lut (.I0(GND_net), .I1(n13698[7]), .I2(n661), 
            .I3(n50839), .O(n12733[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_10 (.CI(n50839), .I0(n13698[7]), .I1(n661), .CO(n50840));
    SB_LUT4 mux_15_i12_3_lut (.I0(n207[11]), .I1(IntegralLimit[11]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[11] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6100_9_lut (.I0(GND_net), .I1(n13698[6]), .I2(n588), .I3(n50838), 
            .O(n12733[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i71_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6100_9 (.CI(n50838), .I0(n13698[6]), .I1(n588), .CO(n50839));
    SB_LUT4 mult_17_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5171));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51613_4_lut (.I0(n24), .I1(n8_adj_5160), .I2(n45), .I3(n66183), 
            .O(n67299));   // verilog/motorControl.v(55[23:39])
    defparam i51613_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_17_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6100_8_lut (.I0(GND_net), .I1(n13698[5]), .I2(n515), .I3(n50837), 
            .O(n12733[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_add_1221_6_lut (.I0(GND_net), .I1(n12109[3]), .I2(n366_adj_5172), 
            .I3(n49813), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50920_3_lut (.I0(n67657), .I1(n432[12]), .I2(n25), .I3(GND_net), 
            .O(n66606));   // verilog/motorControl.v(55[23:39])
    defparam i50920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n615));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i414_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6100_8 (.CI(n50837), .I0(n13698[5]), .I1(n515), .CO(n50838));
    SB_LUT4 mult_17_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n688));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6100_7_lut (.I0(GND_net), .I1(n13698[4]), .I2(n442_adj_5173), 
            .I3(n50836), .O(n12733[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_6 (.CI(n49813), .I0(n12109[3]), .I1(n366_adj_5172), 
            .CO(n49814));
    SB_LUT4 mult_16_add_1221_5_lut (.I0(GND_net), .I1(n12109[2]), .I2(n293_adj_5174), 
            .I3(n49812), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_7 (.CI(n50836), .I0(n13698[4]), .I1(n442_adj_5173), 
            .CO(n50837));
    SB_LUT4 mult_17_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n761));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6100_6_lut (.I0(GND_net), .I1(n13698[3]), .I2(n369_adj_5175), 
            .I3(n50835), .O(n12733[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_6 (.CI(n50835), .I0(n13698[3]), .I1(n369_adj_5175), 
            .CO(n50836));
    SB_LUT4 add_6100_5_lut (.I0(GND_net), .I1(n13698[2]), .I2(n296_adj_5176), 
            .I3(n50834), .O(n12733[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n834));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n907));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i610_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6100_5 (.CI(n50834), .I0(n13698[2]), .I1(n296_adj_5176), 
            .CO(n50835));
    SB_LUT4 mult_17_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n980));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6100_4_lut (.I0(GND_net), .I1(n13698[1]), .I2(n223), .I3(n50833), 
            .O(n12733[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i11_3_lut (.I0(n130[10]), .I1(n182[10]), .I2(n181), 
            .I3(GND_net), .O(n207[10]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6100_4 (.CI(n50833), .I0(n13698[1]), .I1(n223), .CO(n50834));
    SB_LUT4 i51968_3_lut (.I0(n4), .I1(n432[13]), .I2(n27), .I3(GND_net), 
            .O(n67654));   // verilog/motorControl.v(55[23:39])
    defparam i51968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6100_3_lut (.I0(GND_net), .I1(n13698[0]), .I2(n150), .I3(n50832), 
            .O(n12733[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_3 (.CI(n50832), .I0(n13698[0]), .I1(n150), .CO(n50833));
    SB_LUT4 add_6100_2_lut (.I0(GND_net), .I1(n8_adj_5178), .I2(n77), 
            .I3(GND_net), .O(n12733[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6100_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6100_2 (.CI(GND_net), .I0(n8_adj_5178), .I1(n77), .CO(n50832));
    SB_LUT4 add_6143_22_lut (.I0(GND_net), .I1(n14576[19]), .I2(GND_net), 
            .I3(n50831), .O(n13698[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6143_21_lut (.I0(GND_net), .I1(n14576[18]), .I2(GND_net), 
            .I3(n50830), .O(n13698[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_21 (.CI(n50830), .I0(n14576[18]), .I1(GND_net), 
            .CO(n50831));
    SB_LUT4 add_6143_20_lut (.I0(GND_net), .I1(n14576[17]), .I2(GND_net), 
            .I3(n50829), .O(n13698[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_20 (.CI(n50829), .I0(n14576[17]), .I1(GND_net), 
            .CO(n50830));
    SB_LUT4 mult_16_i743_2_lut (.I0(\Kp[15] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6143_19_lut (.I0(GND_net), .I1(n14576[16]), .I2(GND_net), 
            .I3(n50828), .O(n13698[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i11_3_lut (.I0(n207[10]), .I1(IntegralLimit[10]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[10] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51969_3_lut (.I0(n67654), .I1(n432[14]), .I2(n29), .I3(GND_net), 
            .O(n67655));   // verilog/motorControl.v(55[23:39])
    defparam i51969_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_5179));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i69_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6143_19 (.CI(n50828), .I0(n14576[16]), .I1(GND_net), 
            .CO(n50829));
    SB_LUT4 mult_17_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_5180));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_5181));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n55[13]), .I3(n49226), .O(n130[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6143_18_lut (.I0(GND_net), .I1(n14576[15]), .I2(GND_net), 
            .I3(n50827), .O(n13698[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50519_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n66211), 
            .O(n66205));
    defparam i50519_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_6143_18 (.CI(n50827), .I0(n14576[15]), .I1(GND_net), 
            .CO(n50828));
    SB_LUT4 add_6143_17_lut (.I0(GND_net), .I1(n14576[14]), .I2(GND_net), 
            .I3(n50826), .O(n13698[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_17 (.CI(n50826), .I0(n14576[14]), .I1(GND_net), 
            .CO(n50827));
    SB_LUT4 mult_17_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_5182));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_5183));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i510_2_lut (.I0(\Kp[10] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6143_16_lut (.I0(GND_net), .I1(n14576[13]), .I2(n1102_adj_5184), 
            .I3(n50825), .O(n13698[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_16 (.CI(n50825), .I0(n14576[13]), .I1(n1102_adj_5184), 
            .CO(n50826));
    SB_LUT4 add_6143_15_lut (.I0(GND_net), .I1(n14576[12]), .I2(n1029_adj_5185), 
            .I3(n50824), .O(n13698[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_15 (.CI(n50824), .I0(n14576[12]), .I1(n1029_adj_5185), 
            .CO(n50825));
    SB_LUT4 add_6143_14_lut (.I0(GND_net), .I1(n14576[11]), .I2(n956_adj_5186), 
            .I3(n50823), .O(n13698[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_14 (.CI(n50823), .I0(n14576[11]), .I1(n956_adj_5186), 
            .CO(n50824));
    SB_CARRY mult_16_add_1221_5 (.CI(n49812), .I0(n12109[2]), .I1(n293_adj_5174), 
            .CO(n49813));
    SB_LUT4 add_6143_13_lut (.I0(GND_net), .I1(n14576[10]), .I2(n883_adj_5187), 
            .I3(n50822), .O(n13698[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_13 (.CI(n50822), .I0(n14576[10]), .I1(n883_adj_5187), 
            .CO(n50823));
    SB_LUT4 add_6143_12_lut (.I0(GND_net), .I1(n14576[9]), .I2(n810_adj_5188), 
            .I3(n50821), .O(n13698[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_12 (.CI(n50821), .I0(n14576[9]), .I1(n810_adj_5188), 
            .CO(n50822));
    SB_LUT4 add_6143_11_lut (.I0(GND_net), .I1(n14576[8]), .I2(n737_adj_5189), 
            .I3(n50820), .O(n13698[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_11 (.CI(n50820), .I0(n14576[8]), .I1(n737_adj_5189), 
            .CO(n50821));
    SB_LUT4 add_6143_10_lut (.I0(GND_net), .I1(n14576[7]), .I2(n664_adj_5190), 
            .I3(n50819), .O(n13698[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_10 (.CI(n50819), .I0(n14576[7]), .I1(n664_adj_5190), 
            .CO(n50820));
    SB_LUT4 add_6143_9_lut (.I0(GND_net), .I1(n14576[6]), .I2(n591_adj_5191), 
            .I3(n50818), .O(n13698[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_add_1221_4_lut (.I0(GND_net), .I1(n12109[1]), .I2(n220_adj_5192), 
            .I3(n49811), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_4 (.CI(n49811), .I0(n12109[1]), .I1(n220_adj_5192), 
            .CO(n49812));
    SB_LUT4 mult_16_add_1221_3_lut (.I0(GND_net), .I1(n12109[0]), .I2(n147_adj_5194), 
            .I3(n49810), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_3 (.CI(n49810), .I0(n12109[0]), .I1(n147_adj_5194), 
            .CO(n49811));
    SB_CARRY add_6143_9 (.CI(n50818), .I0(n14576[6]), .I1(n591_adj_5191), 
            .CO(n50819));
    SB_LUT4 i50052_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(n130[3]), .I2(n130[2]), 
            .I3(IntegralLimit[2]), .O(n65738));   // verilog/motorControl.v(46[12:34])
    defparam i50052_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_9_11 (.CI(n49226), .I0(\PID_CONTROLLER.integral [9]), .I1(n55[13]), 
            .CO(n49227));
    SB_LUT4 add_6143_8_lut (.I0(GND_net), .I1(n14576[5]), .I2(n518_adj_5195), 
            .I3(n50817), .O(n13698[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_8 (.CI(n50817), .I0(n14576[5]), .I1(n518_adj_5195), 
            .CO(n50818));
    SB_LUT4 mult_16_add_1221_2_lut (.I0(GND_net), .I1(n5_adj_5196), .I2(n74_adj_5197), 
            .I3(GND_net), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_16_add_1221_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6143_7_lut (.I0(GND_net), .I1(n14576[4]), .I2(n445_adj_5198), 
            .I3(n50816), .O(n13698[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_7 (.CI(n50816), .I0(n14576[4]), .I1(n445_adj_5198), 
            .CO(n50817));
    SB_LUT4 add_6143_6_lut (.I0(GND_net), .I1(n14576[3]), .I2(n372_adj_5199), 
            .I3(n50815), .O(n13698[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_16_add_1221_2 (.CI(GND_net), .I0(n5_adj_5196), .I1(n74_adj_5197), 
            .CO(n49810));
    SB_CARRY add_6143_6 (.CI(n50815), .I0(n14576[3]), .I1(n372_adj_5199), 
            .CO(n50816));
    SB_LUT4 add_6143_5_lut (.I0(GND_net), .I1(n14576[2]), .I2(n299_adj_5200), 
            .I3(n50814), .O(n13698[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_5 (.CI(n50814), .I0(n14576[2]), .I1(n299_adj_5200), 
            .CO(n50815));
    SB_LUT4 add_6143_4_lut (.I0(GND_net), .I1(n14576[1]), .I2(n226_adj_5201), 
            .I3(n50813), .O(n13698[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_4 (.CI(n50813), .I0(n14576[1]), .I1(n226_adj_5201), 
            .CO(n50814));
    SB_LUT4 add_6143_3_lut (.I0(GND_net), .I1(n14576[0]), .I2(n153_adj_5202), 
            .I3(n50812), .O(n13698[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52385_4_lut (.I0(n30_c), .I1(n10), .I2(n35), .I3(n66203), 
            .O(n68071));   // verilog/motorControl.v(55[23:39])
    defparam i52385_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_9_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n55[12]), .I3(n49225), .O(n130[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6143_3 (.CI(n50812), .I0(n14576[0]), .I1(n153_adj_5202), 
            .CO(n50813));
    SB_LUT4 add_6143_2_lut (.I0(GND_net), .I1(n11_adj_5203), .I2(n80_adj_5204), 
            .I3(GND_net), .O(n13698[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6143_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_10 (.CI(n49225), .I0(\PID_CONTROLLER.integral [8]), .I1(n55[12]), 
            .CO(n49226));
    SB_CARRY add_6143_2 (.CI(GND_net), .I0(n11_adj_5203), .I1(n80_adj_5204), 
            .CO(n50812));
    SB_LUT4 add_6440_12_lut (.I0(GND_net), .I1(n19365[9]), .I2(n840_adj_5205), 
            .I3(n50811), .O(n19102[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6440_11_lut (.I0(GND_net), .I1(n19365[8]), .I2(n767_adj_5206), 
            .I3(n50810), .O(n19102[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6336_16_lut (.I0(GND_net), .I1(n18009[13]), .I2(n1120), 
            .I3(n49537), .O(n17530[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6336_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_11 (.CI(n50810), .I0(n19365[8]), .I1(n767_adj_5206), 
            .CO(n50811));
    SB_LUT4 add_6440_10_lut (.I0(GND_net), .I1(n19365[7]), .I2(n694_adj_5207), 
            .I3(n50809), .O(n19102[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_10 (.CI(n50809), .I0(n19365[7]), .I1(n694_adj_5207), 
            .CO(n50810));
    SB_LUT4 add_6336_15_lut (.I0(GND_net), .I1(n18009[12]), .I2(n1047), 
            .I3(n49536), .O(n17530[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6336_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6440_9_lut (.I0(GND_net), .I1(n19365[6]), .I2(n621_adj_5208), 
            .I3(n50808), .O(n19102[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_9 (.CI(n50808), .I0(n19365[6]), .I1(n621_adj_5208), 
            .CO(n50809));
    SB_CARRY add_6336_15 (.CI(n49536), .I0(n18009[12]), .I1(n1047), .CO(n49537));
    SB_LUT4 add_6440_8_lut (.I0(GND_net), .I1(n19365[5]), .I2(n548_adj_5209), 
            .I3(n50807), .O(n19102[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6336_14_lut (.I0(GND_net), .I1(n18009[11]), .I2(n974), 
            .I3(n49535), .O(n17530[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6336_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_8 (.CI(n50807), .I0(n19365[5]), .I1(n548_adj_5209), 
            .CO(n50808));
    SB_LUT4 add_6440_7_lut (.I0(GND_net), .I1(n19365[4]), .I2(n475_adj_5210), 
            .I3(n50806), .O(n19102[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_7 (.CI(n50806), .I0(n19365[4]), .I1(n475_adj_5210), 
            .CO(n50807));
    SB_LUT4 add_6440_6_lut (.I0(GND_net), .I1(n19365[3]), .I2(n402_adj_5211), 
            .I3(n50805), .O(n19102[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_6 (.CI(n50805), .I0(n19365[3]), .I1(n402_adj_5211), 
            .CO(n50806));
    SB_LUT4 add_6440_5_lut (.I0(GND_net), .I1(n19365[2]), .I2(n329_adj_5212), 
            .I3(n50804), .O(n19102[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_5 (.CI(n50804), .I0(n19365[2]), .I1(n329_adj_5212), 
            .CO(n50805));
    SB_LUT4 add_6440_4_lut (.I0(GND_net), .I1(n19365[1]), .I2(n256_adj_5213), 
            .I3(n50803), .O(n19102[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_4 (.CI(n50803), .I0(n19365[1]), .I1(n256_adj_5213), 
            .CO(n50804));
    SB_LUT4 unary_minus_26_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[13]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6440_3_lut (.I0(GND_net), .I1(n19365[0]), .I2(n183_adj_5215), 
            .I3(n50802), .O(n19102[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_3 (.CI(n50802), .I0(n19365[0]), .I1(n183_adj_5215), 
            .CO(n50803));
    SB_LUT4 mult_17_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_5216));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6440_2_lut (.I0(GND_net), .I1(n41_adj_5217), .I2(n110_adj_5218), 
            .I3(GND_net), .O(n19102[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6440_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_5219));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n55[11]), .I3(n49224), .O(n130[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6440_2 (.CI(GND_net), .I0(n41_adj_5217), .I1(n110_adj_5218), 
            .CO(n50802));
    SB_LUT4 add_6183_21_lut (.I0(GND_net), .I1(n15372[18]), .I2(GND_net), 
            .I3(n50801), .O(n14576[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6183_20_lut (.I0(GND_net), .I1(n15372[17]), .I2(GND_net), 
            .I3(n50800), .O(n14576[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i559_2_lut (.I0(\Kp[11] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i559_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6183_20 (.CI(n50800), .I0(n15372[17]), .I1(GND_net), 
            .CO(n50801));
    SB_LUT4 add_6183_19_lut (.I0(GND_net), .I1(n15372[16]), .I2(GND_net), 
            .I3(n50799), .O(n14576[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_19 (.CI(n50799), .I0(n15372[16]), .I1(GND_net), 
            .CO(n50800));
    SB_LUT4 add_6183_18_lut (.I0(GND_net), .I1(n15372[15]), .I2(GND_net), 
            .I3(n50798), .O(n14576[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_18 (.CI(n50798), .I0(n15372[15]), .I1(GND_net), 
            .CO(n50799));
    SB_LUT4 add_6183_17_lut (.I0(GND_net), .I1(n15372[14]), .I2(GND_net), 
            .I3(n50797), .O(n14576[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_17 (.CI(n50797), .I0(n15372[14]), .I1(GND_net), 
            .CO(n50798));
    SB_LUT4 add_6183_16_lut (.I0(GND_net), .I1(n15372[13]), .I2(n1105_adj_5221), 
            .I3(n50796), .O(n14576[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_16 (.CI(n50796), .I0(n15372[13]), .I1(n1105_adj_5221), 
            .CO(n50797));
    SB_LUT4 add_6183_15_lut (.I0(GND_net), .I1(n15372[12]), .I2(n1032_adj_5222), 
            .I3(n50795), .O(n14576[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_15 (.CI(n50795), .I0(n15372[12]), .I1(n1032_adj_5222), 
            .CO(n50796));
    SB_LUT4 add_6183_14_lut (.I0(GND_net), .I1(n15372[11]), .I2(n959_adj_5223), 
            .I3(n50794), .O(n14576[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_14 (.CI(n50794), .I0(n15372[11]), .I1(n959_adj_5223), 
            .CO(n50795));
    SB_LUT4 add_6183_13_lut (.I0(GND_net), .I1(n15372[10]), .I2(n886_adj_5224), 
            .I3(n50793), .O(n14576[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_13 (.CI(n50793), .I0(n15372[10]), .I1(n886_adj_5224), 
            .CO(n50794));
    SB_LUT4 add_6183_12_lut (.I0(GND_net), .I1(n15372[9]), .I2(n813), 
            .I3(n50792), .O(n14576[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_12 (.CI(n50792), .I0(n15372[9]), .I1(n813), .CO(n50793));
    SB_LUT4 add_6183_11_lut (.I0(GND_net), .I1(n15372[8]), .I2(n740), 
            .I3(n50791), .O(n14576[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50922_3_lut (.I0(n67655), .I1(n432[15]), .I2(n31), .I3(GND_net), 
            .O(n66608));   // verilog/motorControl.v(55[23:39])
    defparam i50922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52561_4_lut (.I0(n66608), .I1(n68071), .I2(n35), .I3(n66205), 
            .O(n68247));   // verilog/motorControl.v(55[23:39])
    defparam i52561_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52562_3_lut (.I0(n68247), .I1(n432[18]), .I2(n37), .I3(GND_net), 
            .O(n68248));   // verilog/motorControl.v(55[23:39])
    defparam i52562_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52516_3_lut (.I0(n68248), .I1(n432[19]), .I2(n39_adj_5225), 
            .I3(GND_net), .O(n68202));   // verilog/motorControl.v(55[23:39])
    defparam i52516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50501_4_lut (.I0(n43_c), .I1(n41_adj_5226), .I2(n39_adj_5225), 
            .I3(n68148), .O(n66187));
    defparam i50501_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52242_4_lut (.I0(n66606), .I1(n67299), .I2(n45), .I3(n66185), 
            .O(n67928));   // verilog/motorControl.v(55[23:39])
    defparam i52242_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i50928_3_lut (.I0(n68202), .I1(n432[20]), .I2(n41_adj_5226), 
            .I3(GND_net), .O(n66614));   // verilog/motorControl.v(55[23:39])
    defparam i50928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52439_4_lut (.I0(n66614), .I1(n67928), .I2(n45), .I3(n66187), 
            .O(n68125));   // verilog/motorControl.v(55[23:39])
    defparam i52439_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52440_3_lut (.I0(n68125), .I1(n352[23]), .I2(n432[23]), .I3(GND_net), 
            .O(n68126));   // verilog/motorControl.v(55[23:39])
    defparam i52440_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i5969_3_lut (.I0(control_update), .I1(n405), .I2(n68126), 
            .I3(GND_net), .O(n11610));   // verilog/motorControl.v(20[7:21])
    defparam i5969_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i28859_4_lut (.I0(PWMLimit[0]), .I1(n60219), .I2(n27692), 
            .I3(n11608), .O(n51[0]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i28859_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY add_6183_11 (.CI(n50791), .I0(n15372[8]), .I1(n740), .CO(n50792));
    SB_LUT4 add_6183_10_lut (.I0(GND_net), .I1(n15372[7]), .I2(n667), 
            .I3(n50790), .O(n14576[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_10 (.CI(n50790), .I0(n15372[7]), .I1(n667), .CO(n50791));
    SB_LUT4 add_6183_9_lut (.I0(GND_net), .I1(n15372[6]), .I2(n594), .I3(n50789), 
            .O(n14576[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_5227));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i363_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6183_9 (.CI(n50789), .I0(n15372[6]), .I1(n594), .CO(n50790));
    SB_LUT4 add_6183_8_lut (.I0(GND_net), .I1(n15372[5]), .I2(n521), .I3(n50788), 
            .O(n14576[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_8 (.CI(n50788), .I0(n15372[5]), .I1(n521), .CO(n50789));
    SB_CARRY add_6336_14 (.CI(n49535), .I0(n18009[11]), .I1(n974), .CO(n49536));
    SB_CARRY add_9_9 (.CI(n49224), .I0(\PID_CONTROLLER.integral [7]), .I1(n55[11]), 
            .CO(n49225));
    SB_LUT4 add_6183_7_lut (.I0(GND_net), .I1(n15372[4]), .I2(n448_adj_5228), 
            .I3(n50787), .O(n14576[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_7 (.CI(n50787), .I0(n15372[4]), .I1(n448_adj_5228), 
            .CO(n50788));
    SB_LUT4 add_6183_6_lut (.I0(GND_net), .I1(n15372[3]), .I2(n375_c), 
            .I3(n50786), .O(n14576[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_6 (.CI(n50786), .I0(n15372[3]), .I1(n375_c), .CO(n50787));
    SB_LUT4 add_6183_5_lut (.I0(GND_net), .I1(n15372[2]), .I2(n302), .I3(n50785), 
            .O(n14576[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_5 (.CI(n50785), .I0(n15372[2]), .I1(n302), .CO(n50786));
    SB_LUT4 add_6183_4_lut (.I0(GND_net), .I1(n15372[1]), .I2(n229), .I3(n50784), 
            .O(n14576[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_4 (.CI(n50784), .I0(n15372[1]), .I1(n229), .CO(n50785));
    SB_LUT4 add_6183_3_lut (.I0(GND_net), .I1(n15372[0]), .I2(n156), .I3(n50783), 
            .O(n14576[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6473_11_lut (.I0(GND_net), .I1(n19702[8]), .I2(n770), 
            .I3(n49791), .O(n19506[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n55[10]), .I3(n49223), .O(n130[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_3 (.CI(n50783), .I0(n15372[0]), .I1(n156), .CO(n50784));
    SB_LUT4 add_6183_2_lut (.I0(GND_net), .I1(n14_adj_5229), .I2(n83), 
            .I3(GND_net), .O(n14576[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6183_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6183_2 (.CI(GND_net), .I0(n14_adj_5229), .I1(n83), .CO(n50783));
    SB_LUT4 add_6221_20_lut (.I0(GND_net), .I1(n16090[17]), .I2(GND_net), 
            .I3(n50782), .O(n15372[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6221_19_lut (.I0(GND_net), .I1(n16090[16]), .I2(GND_net), 
            .I3(n50781), .O(n15372[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_19 (.CI(n50781), .I0(n16090[16]), .I1(GND_net), 
            .CO(n50782));
    SB_LUT4 add_6221_18_lut (.I0(GND_net), .I1(n16090[15]), .I2(GND_net), 
            .I3(n50780), .O(n15372[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_18 (.CI(n50780), .I0(n16090[15]), .I1(GND_net), 
            .CO(n50781));
    SB_LUT4 add_6221_17_lut (.I0(GND_net), .I1(n16090[14]), .I2(GND_net), 
            .I3(n50779), .O(n15372[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n612_adj_5230));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i412_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6221_17 (.CI(n50779), .I0(n16090[14]), .I1(GND_net), 
            .CO(n50780));
    SB_LUT4 mult_16_i608_2_lut (.I0(\Kp[12] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6221_16_lut (.I0(GND_net), .I1(n16090[13]), .I2(n1108), 
            .I3(n50778), .O(n15372[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_16 (.CI(n50778), .I0(n16090[13]), .I1(n1108), .CO(n50779));
    SB_LUT4 add_6221_15_lut (.I0(GND_net), .I1(n16090[12]), .I2(n1035), 
            .I3(n50777), .O(n15372[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_15 (.CI(n50777), .I0(n16090[12]), .I1(n1035), .CO(n50778));
    SB_LUT4 add_6221_14_lut (.I0(GND_net), .I1(n16090[11]), .I2(n962), 
            .I3(n50776), .O(n15372[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_14 (.CI(n50776), .I0(n16090[11]), .I1(n962), .CO(n50777));
    SB_LUT4 add_6221_13_lut (.I0(GND_net), .I1(n16090[10]), .I2(n889), 
            .I3(n50775), .O(n15372[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_13 (.CI(n50775), .I0(n16090[10]), .I1(n889), .CO(n50776));
    SB_LUT4 add_6473_10_lut (.I0(GND_net), .I1(n19702[7]), .I2(n697), 
            .I3(n49790), .O(n19506[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6221_12_lut (.I0(GND_net), .I1(n16090[9]), .I2(n816), 
            .I3(n50774), .O(n15372[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6473_10 (.CI(n49790), .I0(n19702[7]), .I1(n697), .CO(n49791));
    SB_CARRY add_6221_12 (.CI(n50774), .I0(n16090[9]), .I1(n816), .CO(n50775));
    SB_LUT4 add_6221_11_lut (.I0(GND_net), .I1(n16090[8]), .I2(n743), 
            .I3(n50773), .O(n15372[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_11 (.CI(n50773), .I0(n16090[8]), .I1(n743), .CO(n50774));
    SB_LUT4 add_6473_9_lut (.I0(GND_net), .I1(n19702[6]), .I2(n624), .I3(n49789), 
            .O(n19506[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6221_10_lut (.I0(GND_net), .I1(n16090[7]), .I2(n670), 
            .I3(n50772), .O(n15372[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_10 (.CI(n50772), .I0(n16090[7]), .I1(n670), .CO(n50773));
    SB_LUT4 add_6221_9_lut (.I0(GND_net), .I1(n16090[6]), .I2(n597), .I3(n50771), 
            .O(n15372[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_9 (.CI(n50771), .I0(n16090[6]), .I1(n597), .CO(n50772));
    SB_LUT4 add_6221_8_lut (.I0(GND_net), .I1(n16090[5]), .I2(n524), .I3(n50770), 
            .O(n15372[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_8 (.CI(n50770), .I0(n16090[5]), .I1(n524), .CO(n50771));
    SB_LUT4 add_6221_7_lut (.I0(GND_net), .I1(n16090[4]), .I2(n451_adj_5231), 
            .I3(n50769), .O(n15372[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_7 (.CI(n50769), .I0(n16090[4]), .I1(n451_adj_5231), 
            .CO(n50770));
    SB_LUT4 add_6221_6_lut (.I0(GND_net), .I1(n16090[3]), .I2(n378), .I3(n50768), 
            .O(n15372[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_6 (.CI(n50768), .I0(n16090[3]), .I1(n378), .CO(n50769));
    SB_LUT4 add_6221_5_lut (.I0(GND_net), .I1(n16090[2]), .I2(n305), .I3(n50767), 
            .O(n15372[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6473_9 (.CI(n49789), .I0(n19702[6]), .I1(n624), .CO(n49790));
    SB_CARRY add_6221_5 (.CI(n50767), .I0(n16090[2]), .I1(n305), .CO(n50768));
    SB_LUT4 add_6221_4_lut (.I0(GND_net), .I1(n16090[1]), .I2(n232), .I3(n50766), 
            .O(n15372[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_4 (.CI(n50766), .I0(n16090[1]), .I1(n232), .CO(n50767));
    SB_LUT4 add_6221_3_lut (.I0(GND_net), .I1(n16090[0]), .I2(n159), .I3(n50765), 
            .O(n15372[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_3 (.CI(n50765), .I0(n16090[0]), .I1(n159), .CO(n50766));
    SB_LUT4 add_6221_2_lut (.I0(GND_net), .I1(n17_adj_5232), .I2(n86), 
            .I3(GND_net), .O(n15372[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6221_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6221_2 (.CI(GND_net), .I0(n17_adj_5232), .I1(n86), .CO(n50765));
    SB_LUT4 add_6461_11_lut (.I0(GND_net), .I1(n19584[8]), .I2(n770_adj_5233), 
            .I3(n50764), .O(n19365[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6461_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6473_8_lut (.I0(GND_net), .I1(n19702[5]), .I2(n551), .I3(n49788), 
            .O(n19506[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6461_10_lut (.I0(GND_net), .I1(n19584[7]), .I2(n697_adj_5234), 
            .I3(n50763), .O(n19365[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6461_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6461_10 (.CI(n50763), .I0(n19584[7]), .I1(n697_adj_5234), 
            .CO(n50764));
    SB_LUT4 add_6336_13_lut (.I0(GND_net), .I1(n18009[10]), .I2(n901), 
            .I3(n49534), .O(n17530[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6336_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6461_9_lut (.I0(GND_net), .I1(n19584[6]), .I2(n624_adj_5235), 
            .I3(n50762), .O(n19365[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6461_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6461_9 (.CI(n50762), .I0(n19584[6]), .I1(n624_adj_5235), 
            .CO(n50763));
    SB_CARRY add_6336_13 (.CI(n49534), .I0(n18009[10]), .I1(n901), .CO(n49535));
    SB_CARRY add_6473_8 (.CI(n49788), .I0(n19702[5]), .I1(n551), .CO(n49789));
    SB_LUT4 add_6473_7_lut (.I0(GND_net), .I1(n19702[4]), .I2(n478), .I3(n49787), 
            .O(n19506[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6461_8_lut (.I0(GND_net), .I1(n19584[5]), .I2(n551_adj_5236), 
            .I3(n50761), .O(n19365[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6461_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6461_8 (.CI(n50761), .I0(n19584[5]), .I1(n551_adj_5236), 
            .CO(n50762));
    SB_LUT4 add_6461_7_lut (.I0(GND_net), .I1(n19584[4]), .I2(n478_adj_5237), 
            .I3(n50760), .O(n19365[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6461_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i6_3_lut_3_lut (.I0(IntegralLimit[3]), .I1(n130[3]), 
            .I2(n130[2]), .I3(GND_net), .O(n6_adj_5238));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_16_i657_2_lut (.I0(\Kp[13] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n685_adj_5239));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i461_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6461_7 (.CI(n50760), .I0(n19584[4]), .I1(n478_adj_5237), 
            .CO(n50761));
    SB_LUT4 add_6461_6_lut (.I0(GND_net), .I1(n19584[3]), .I2(n405_adj_5240), 
            .I3(n50759), .O(n19365[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6461_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6461_6 (.CI(n50759), .I0(n19584[3]), .I1(n405_adj_5240), 
            .CO(n50760));
    SB_LUT4 add_6461_5_lut (.I0(GND_net), .I1(n19584[2]), .I2(n332_adj_5241), 
            .I3(n50758), .O(n19365[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6461_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6461_5 (.CI(n50758), .I0(n19584[2]), .I1(n332_adj_5241), 
            .CO(n50759));
    SB_LUT4 add_6461_4_lut (.I0(GND_net), .I1(n19584[1]), .I2(n259), .I3(n50757), 
            .O(n19365[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6461_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6461_4 (.CI(n50757), .I0(n19584[1]), .I1(n259), .CO(n50758));
    SB_LUT4 add_6461_3_lut (.I0(GND_net), .I1(n19584[0]), .I2(n186_adj_5242), 
            .I3(n50756), .O(n19365[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6461_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6461_3 (.CI(n50756), .I0(n19584[0]), .I1(n186_adj_5242), 
            .CO(n50757));
    SB_LUT4 add_6461_2_lut (.I0(GND_net), .I1(n44), .I2(n113_adj_5243), 
            .I3(GND_net), .O(n19365[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6461_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6461_2 (.CI(GND_net), .I0(n44), .I1(n113_adj_5243), .CO(n50756));
    SB_LUT4 add_6257_19_lut (.I0(GND_net), .I1(n16734[16]), .I2(GND_net), 
            .I3(n50755), .O(n16090[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6257_18_lut (.I0(GND_net), .I1(n16734[15]), .I2(GND_net), 
            .I3(n50754), .O(n16090[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_8 (.CI(n49223), .I0(\PID_CONTROLLER.integral [6]), .I1(n55[10]), 
            .CO(n49224));
    SB_CARRY add_6257_18 (.CI(n50754), .I0(n16734[15]), .I1(GND_net), 
            .CO(n50755));
    SB_LUT4 add_6257_17_lut (.I0(GND_net), .I1(n16734[14]), .I2(GND_net), 
            .I3(n50753), .O(n16090[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6336_12_lut (.I0(GND_net), .I1(n18009[9]), .I2(n828), 
            .I3(n49533), .O(n17530[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6336_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_17 (.CI(n50753), .I0(n16734[14]), .I1(GND_net), 
            .CO(n50754));
    SB_LUT4 add_6257_16_lut (.I0(GND_net), .I1(n16734[13]), .I2(n1111), 
            .I3(n50752), .O(n16090[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_16 (.CI(n50752), .I0(n16734[13]), .I1(n1111), .CO(n50753));
    SB_LUT4 add_6257_15_lut (.I0(GND_net), .I1(n16734[12]), .I2(n1038), 
            .I3(n50751), .O(n16090[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_15 (.CI(n50751), .I0(n16734[12]), .I1(n1038), .CO(n50752));
    SB_CARRY add_6336_12 (.CI(n49533), .I0(n18009[9]), .I1(n828), .CO(n49534));
    SB_LUT4 add_6257_14_lut (.I0(GND_net), .I1(n16734[11]), .I2(n965), 
            .I3(n50750), .O(n16090[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n55[9]), .I3(n49222), .O(n130[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_14 (.CI(n50750), .I0(n16734[11]), .I1(n965), .CO(n50751));
    SB_LUT4 add_6257_13_lut (.I0(GND_net), .I1(n16734[10]), .I2(n892), 
            .I3(n50749), .O(n16090[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_13 (.CI(n50749), .I0(n16734[10]), .I1(n892), .CO(n50750));
    SB_LUT4 add_6257_12_lut (.I0(GND_net), .I1(n16734[9]), .I2(n819), 
            .I3(n50748), .O(n16090[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_12 (.CI(n50748), .I0(n16734[9]), .I1(n819), .CO(n50749));
    SB_LUT4 add_6257_11_lut (.I0(GND_net), .I1(n16734[8]), .I2(n746), 
            .I3(n50747), .O(n16090[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_11 (.CI(n50747), .I0(n16734[8]), .I1(n746), .CO(n50748));
    SB_LUT4 add_6257_10_lut (.I0(GND_net), .I1(n16734[7]), .I2(n673), 
            .I3(n50746), .O(n16090[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_10 (.CI(n50746), .I0(n16734[7]), .I1(n673), .CO(n50747));
    SB_LUT4 add_6257_9_lut (.I0(GND_net), .I1(n16734[6]), .I2(n600), .I3(n50745), 
            .O(n16090[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_9 (.CI(n50745), .I0(n16734[6]), .I1(n600), .CO(n50746));
    SB_LUT4 add_6257_8_lut (.I0(GND_net), .I1(n16734[5]), .I2(n527), .I3(n50744), 
            .O(n16090[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_8 (.CI(n50744), .I0(n16734[5]), .I1(n527), .CO(n50745));
    SB_LUT4 add_6257_7_lut (.I0(GND_net), .I1(n16734[4]), .I2(n454), .I3(n50743), 
            .O(n16090[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_7 (.CI(n50743), .I0(n16734[4]), .I1(n454), .CO(n50744));
    SB_LUT4 add_6257_6_lut (.I0(GND_net), .I1(n16734[3]), .I2(n381), .I3(n50742), 
            .O(n16090[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_6 (.CI(n50742), .I0(n16734[3]), .I1(n381), .CO(n50743));
    SB_LUT4 add_6257_5_lut (.I0(GND_net), .I1(n16734[2]), .I2(n308), .I3(n50741), 
            .O(n16090[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_5 (.CI(n50741), .I0(n16734[2]), .I1(n308), .CO(n50742));
    SB_LUT4 add_6257_4_lut (.I0(GND_net), .I1(n16734[1]), .I2(n235), .I3(n50740), 
            .O(n16090[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_4 (.CI(n50740), .I0(n16734[1]), .I1(n235), .CO(n50741));
    SB_LUT4 add_6257_3_lut (.I0(GND_net), .I1(n16734[0]), .I2(n162), .I3(n50739), 
            .O(n16090[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6473_7 (.CI(n49787), .I0(n19702[4]), .I1(n478), .CO(n49788));
    SB_CARRY add_6257_3 (.CI(n50739), .I0(n16734[0]), .I1(n162), .CO(n50740));
    SB_CARRY add_9_7 (.CI(n49222), .I0(\PID_CONTROLLER.integral [5]), .I1(n55[9]), 
            .CO(n49223));
    SB_LUT4 add_6257_2_lut (.I0(GND_net), .I1(n20_adj_5244), .I2(n89), 
            .I3(GND_net), .O(n16090[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6257_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6257_2 (.CI(GND_net), .I0(n20_adj_5244), .I1(n89), .CO(n50739));
    SB_LUT4 add_6291_18_lut (.I0(GND_net), .I1(n17308[15]), .I2(GND_net), 
            .I3(n50738), .O(n16734[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6291_17_lut (.I0(GND_net), .I1(n17308[14]), .I2(GND_net), 
            .I3(n50737), .O(n16734[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_17 (.CI(n50737), .I0(n17308[14]), .I1(GND_net), 
            .CO(n50738));
    SB_LUT4 add_6291_16_lut (.I0(GND_net), .I1(n17308[13]), .I2(n1114_adj_5245), 
            .I3(n50736), .O(n16734[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_16 (.CI(n50736), .I0(n17308[13]), .I1(n1114_adj_5245), 
            .CO(n50737));
    SB_LUT4 add_6291_15_lut (.I0(GND_net), .I1(n17308[12]), .I2(n1041_adj_5246), 
            .I3(n50735), .O(n16734[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_15 (.CI(n50735), .I0(n17308[12]), .I1(n1041_adj_5246), 
            .CO(n50736));
    SB_LUT4 add_6291_14_lut (.I0(GND_net), .I1(n17308[11]), .I2(n968_adj_5247), 
            .I3(n50734), .O(n16734[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_14 (.CI(n50734), .I0(n17308[11]), .I1(n968_adj_5247), 
            .CO(n50735));
    SB_LUT4 add_6291_13_lut (.I0(GND_net), .I1(n17308[10]), .I2(n895_adj_5248), 
            .I3(n50733), .O(n16734[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_13 (.CI(n50733), .I0(n17308[10]), .I1(n895_adj_5248), 
            .CO(n50734));
    SB_LUT4 add_6291_12_lut (.I0(GND_net), .I1(n17308[9]), .I2(n822_adj_5249), 
            .I3(n50732), .O(n16734[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_12 (.CI(n50732), .I0(n17308[9]), .I1(n822_adj_5249), 
            .CO(n50733));
    SB_LUT4 add_6291_11_lut (.I0(GND_net), .I1(n17308[8]), .I2(n749_adj_5250), 
            .I3(n50731), .O(n16734[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_11 (.CI(n50731), .I0(n17308[8]), .I1(n749_adj_5250), 
            .CO(n50732));
    SB_LUT4 add_6473_6_lut (.I0(GND_net), .I1(n19702[3]), .I2(n405_adj_5251), 
            .I3(n49786), .O(n19506[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6291_10_lut (.I0(GND_net), .I1(n17308[7]), .I2(n676_adj_5252), 
            .I3(n50730), .O(n16734[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_10 (.CI(n50730), .I0(n17308[7]), .I1(n676_adj_5252), 
            .CO(n50731));
    SB_LUT4 add_6291_9_lut (.I0(GND_net), .I1(n17308[6]), .I2(n603_adj_5253), 
            .I3(n50729), .O(n16734[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i53_2_lut (.I0(\Kp[1] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_5254));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6336_11_lut (.I0(GND_net), .I1(n18009[8]), .I2(n755), 
            .I3(n49532), .O(n17530[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6336_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6336_11 (.CI(n49532), .I0(n18009[8]), .I1(n755), .CO(n49533));
    SB_CARRY add_6291_9 (.CI(n50729), .I0(n17308[6]), .I1(n603_adj_5253), 
            .CO(n50730));
    SB_LUT4 add_6291_8_lut (.I0(GND_net), .I1(n17308[5]), .I2(n530_adj_5255), 
            .I3(n50728), .O(n16734[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_8 (.CI(n50728), .I0(n17308[5]), .I1(n530_adj_5255), 
            .CO(n50729));
    SB_LUT4 add_6336_10_lut (.I0(GND_net), .I1(n18009[7]), .I2(n682), 
            .I3(n49531), .O(n17530[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6336_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6291_7_lut (.I0(GND_net), .I1(n17308[4]), .I2(n457_adj_5256), 
            .I3(n50727), .O(n16734[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_7 (.CI(n50727), .I0(n17308[4]), .I1(n457_adj_5256), 
            .CO(n50728));
    SB_LUT4 add_6291_6_lut (.I0(GND_net), .I1(n17308[3]), .I2(n384_adj_5257), 
            .I3(n50726), .O(n16734[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_6 (.CI(n50726), .I0(n17308[3]), .I1(n384_adj_5257), 
            .CO(n50727));
    SB_CARRY add_6336_10 (.CI(n49531), .I0(n18009[7]), .I1(n682), .CO(n49532));
    SB_LUT4 add_6291_5_lut (.I0(GND_net), .I1(n17308[2]), .I2(n311_adj_5258), 
            .I3(n50725), .O(n16734[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_5 (.CI(n50725), .I0(n17308[2]), .I1(n311_adj_5258), 
            .CO(n50726));
    SB_LUT4 add_6291_4_lut (.I0(GND_net), .I1(n17308[1]), .I2(n238_adj_5259), 
            .I3(n50724), .O(n16734[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6473_6 (.CI(n49786), .I0(n19702[3]), .I1(n405_adj_5251), 
            .CO(n49787));
    SB_CARRY add_6291_4 (.CI(n50724), .I0(n17308[1]), .I1(n238_adj_5259), 
            .CO(n50725));
    SB_LUT4 add_6473_5_lut (.I0(GND_net), .I1(n19702[2]), .I2(n332_adj_5260), 
            .I3(n49785), .O(n19506[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6291_3_lut (.I0(GND_net), .I1(n17308[0]), .I2(n165_adj_5261), 
            .I3(n50723), .O(n16734[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6336_9_lut (.I0(GND_net), .I1(n18009[6]), .I2(n609), .I3(n49530), 
            .O(n17530[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6336_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_3 (.CI(n50723), .I0(n17308[0]), .I1(n165_adj_5261), 
            .CO(n50724));
    SB_LUT4 add_9_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n55[8]), .I3(n49221), .O(n130[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6291_2_lut (.I0(GND_net), .I1(n23_adj_5263), .I2(n92_adj_5264), 
            .I3(GND_net), .O(n16734[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6291_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6291_2 (.CI(GND_net), .I0(n23_adj_5263), .I1(n92_adj_5264), 
            .CO(n50723));
    SB_CARRY add_6473_5 (.CI(n49785), .I0(n19702[2]), .I1(n332_adj_5260), 
            .CO(n49786));
    SB_LUT4 mult_16_i6_2_lut (.I0(\Kp[0] ), .I1(n55[6]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_5265));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6480_10_lut (.I0(GND_net), .I1(n19763[7]), .I2(n700), 
            .I3(n50722), .O(n19584[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6480_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6336_9 (.CI(n49530), .I0(n18009[6]), .I1(n609), .CO(n49531));
    SB_LUT4 add_6336_8_lut (.I0(GND_net), .I1(n18009[5]), .I2(n536), .I3(n49529), 
            .O(n17530[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6336_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6480_9_lut (.I0(GND_net), .I1(n19763[6]), .I2(n627), .I3(n50721), 
            .O(n19584[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6480_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_6 (.CI(n49221), .I0(\PID_CONTROLLER.integral [4]), .I1(n55[8]), 
            .CO(n49222));
    SB_LUT4 add_6473_4_lut (.I0(GND_net), .I1(n19702[1]), .I2(n259_adj_5266), 
            .I3(n49784), .O(n19506[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6480_9 (.CI(n50721), .I0(n19763[6]), .I1(n627), .CO(n50722));
    SB_CARRY add_6336_8 (.CI(n49529), .I0(n18009[5]), .I1(n536), .CO(n49530));
    SB_LUT4 add_6336_7_lut (.I0(GND_net), .I1(n18009[4]), .I2(n463), .I3(n49528), 
            .O(n17530[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6336_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6480_8_lut (.I0(GND_net), .I1(n19763[5]), .I2(n554), .I3(n50720), 
            .O(n19584[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6480_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6480_8 (.CI(n50720), .I0(n19763[5]), .I1(n554), .CO(n50721));
    SB_LUT4 mult_17_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n758_adj_5267));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6480_7_lut (.I0(GND_net), .I1(n19763[4]), .I2(n481), .I3(n50719), 
            .O(n19584[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6480_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6480_7 (.CI(n50719), .I0(n19763[4]), .I1(n481), .CO(n50720));
    SB_LUT4 add_6480_6_lut (.I0(GND_net), .I1(n19763[3]), .I2(n408), .I3(n50718), 
            .O(n19584[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6480_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6336_7 (.CI(n49528), .I0(n18009[4]), .I1(n463), .CO(n49529));
    SB_CARRY add_6480_6 (.CI(n50718), .I0(n19763[3]), .I1(n408), .CO(n50719));
    SB_CARRY add_6473_4 (.CI(n49784), .I0(n19702[1]), .I1(n259_adj_5266), 
            .CO(n49785));
    SB_LUT4 add_6480_5_lut (.I0(GND_net), .I1(n19763[2]), .I2(n335_adj_5268), 
            .I3(n50717), .O(n19584[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6480_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6336_6_lut (.I0(GND_net), .I1(n18009[3]), .I2(n390), .I3(n49527), 
            .O(n17530[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6336_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6480_5 (.CI(n50717), .I0(n19763[2]), .I1(n335_adj_5268), 
            .CO(n50718));
    SB_LUT4 add_6480_4_lut (.I0(GND_net), .I1(n19763[1]), .I2(n262), .I3(n50716), 
            .O(n19584[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6480_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6336_6 (.CI(n49527), .I0(n18009[3]), .I1(n390), .CO(n49528));
    SB_CARRY add_6480_4 (.CI(n50716), .I0(n19763[1]), .I1(n262), .CO(n50717));
    SB_LUT4 add_6473_3_lut (.I0(GND_net), .I1(n19702[0]), .I2(n186_adj_5269), 
            .I3(n49783), .O(n19506[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6480_3_lut (.I0(GND_net), .I1(n19763[0]), .I2(n189), .I3(n50715), 
            .O(n19584[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6480_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6480_3 (.CI(n50715), .I0(n19763[0]), .I1(n189), .CO(n50716));
    SB_CARRY add_6473_3 (.CI(n49783), .I0(n19702[0]), .I1(n186_adj_5269), 
            .CO(n49784));
    SB_LUT4 mult_17_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n831_adj_5270));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6480_2_lut (.I0(GND_net), .I1(n47), .I2(n116_adj_5271), 
            .I3(GND_net), .O(n19584[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6480_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6336_5_lut (.I0(GND_net), .I1(n18009[2]), .I2(n317), .I3(n49526), 
            .O(n17530[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6336_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6480_2 (.CI(GND_net), .I0(n47), .I1(n116_adj_5271), .CO(n50715));
    SB_LUT4 add_6323_17_lut (.I0(GND_net), .I1(n17816[14]), .I2(GND_net), 
            .I3(n50714), .O(n17308[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6323_16_lut (.I0(GND_net), .I1(n17816[13]), .I2(n1117_adj_5272), 
            .I3(n50713), .O(n17308[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_16 (.CI(n50713), .I0(n17816[13]), .I1(n1117_adj_5272), 
            .CO(n50714));
    SB_LUT4 add_6323_15_lut (.I0(GND_net), .I1(n17816[12]), .I2(n1044_adj_5273), 
            .I3(n50712), .O(n17308[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_15 (.CI(n50712), .I0(n17816[12]), .I1(n1044_adj_5273), 
            .CO(n50713));
    SB_LUT4 add_6323_14_lut (.I0(GND_net), .I1(n17816[11]), .I2(n971_adj_5274), 
            .I3(n50711), .O(n17308[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_14 (.CI(n50711), .I0(n17816[11]), .I1(n971_adj_5274), 
            .CO(n50712));
    SB_LUT4 mult_16_i102_2_lut (.I0(\Kp[2] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_5275));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6323_13_lut (.I0(GND_net), .I1(n17816[10]), .I2(n898_adj_5276), 
            .I3(n50710), .O(n17308[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_13 (.CI(n50710), .I0(n17816[10]), .I1(n898_adj_5276), 
            .CO(n50711));
    SB_LUT4 add_6323_12_lut (.I0(GND_net), .I1(n17816[9]), .I2(n825_adj_5277), 
            .I3(n50709), .O(n17308[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_12 (.CI(n50709), .I0(n17816[9]), .I1(n825_adj_5277), 
            .CO(n50710));
    SB_LUT4 add_6323_11_lut (.I0(GND_net), .I1(n17816[8]), .I2(n752_adj_5278), 
            .I3(n50708), .O(n17308[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_11 (.CI(n50708), .I0(n17816[8]), .I1(n752_adj_5278), 
            .CO(n50709));
    SB_CARRY add_6336_5 (.CI(n49526), .I0(n18009[2]), .I1(n317), .CO(n49527));
    SB_LUT4 add_6323_10_lut (.I0(GND_net), .I1(n17816[7]), .I2(n679_adj_5279), 
            .I3(n50707), .O(n17308[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6473_2_lut (.I0(GND_net), .I1(n44_adj_5280), .I2(n113_adj_5281), 
            .I3(GND_net), .O(n19506[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6473_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_10 (.CI(n50707), .I0(n17816[7]), .I1(n679_adj_5279), 
            .CO(n50708));
    SB_LUT4 unary_minus_26_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[0]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6323_9_lut (.I0(GND_net), .I1(n17816[6]), .I2(n606_adj_5283), 
            .I3(n50706), .O(n17308[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_9 (.CI(n50706), .I0(n17816[6]), .I1(n606_adj_5283), 
            .CO(n50707));
    SB_LUT4 add_6336_4_lut (.I0(GND_net), .I1(n18009[1]), .I2(n244), .I3(n49525), 
            .O(n17530[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6336_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6336_4 (.CI(n49525), .I0(n18009[1]), .I1(n244), .CO(n49526));
    SB_LUT4 add_6323_8_lut (.I0(GND_net), .I1(n17816[5]), .I2(n533_adj_5284), 
            .I3(n50705), .O(n17308[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_5285));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6336_3_lut (.I0(GND_net), .I1(n18009[0]), .I2(n171), .I3(n49524), 
            .O(n17530[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6336_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_8 (.CI(n50705), .I0(n17816[5]), .I1(n533_adj_5284), 
            .CO(n50706));
    SB_LUT4 add_6323_7_lut (.I0(GND_net), .I1(n17816[4]), .I2(n460_adj_5286), 
            .I3(n50704), .O(n17308[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i706_2_lut (.I0(\Kp[14] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i706_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6323_7 (.CI(n50704), .I0(n17816[4]), .I1(n460_adj_5286), 
            .CO(n50705));
    SB_LUT4 add_6323_6_lut (.I0(GND_net), .I1(n17816[3]), .I2(n387_adj_5287), 
            .I3(n50703), .O(n17308[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_6 (.CI(n50703), .I0(n17816[3]), .I1(n387_adj_5287), 
            .CO(n50704));
    SB_LUT4 add_6323_5_lut (.I0(GND_net), .I1(n17816[2]), .I2(n314_adj_5288), 
            .I3(n50702), .O(n17308[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_5 (.CI(n50702), .I0(n17816[2]), .I1(n314_adj_5288), 
            .CO(n50703));
    SB_LUT4 add_6323_4_lut (.I0(GND_net), .I1(n17816[1]), .I2(n241_adj_5289), 
            .I3(n50701), .O(n17308[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6473_2 (.CI(GND_net), .I0(n44_adj_5280), .I1(n113_adj_5281), 
            .CO(n49783));
    SB_LUT4 add_6050_23_lut (.I0(GND_net), .I1(n13171[20]), .I2(GND_net), 
            .I3(n49782), .O(n12109[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_4 (.CI(n50701), .I0(n17816[1]), .I1(n241_adj_5289), 
            .CO(n50702));
    SB_CARRY add_6336_3 (.CI(n49524), .I0(n18009[0]), .I1(n171), .CO(n49525));
    SB_LUT4 mult_17_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n977_adj_5290));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6336_2_lut (.I0(GND_net), .I1(n29_adj_5291), .I2(n98), 
            .I3(GND_net), .O(n17530[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6336_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n55[7]), .I3(n49220), .O(n130[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6336_2 (.CI(GND_net), .I0(n29_adj_5291), .I1(n98), .CO(n49524));
    SB_LUT4 add_6050_22_lut (.I0(GND_net), .I1(n13171[19]), .I2(GND_net), 
            .I3(n49781), .O(n12109[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6323_3_lut (.I0(GND_net), .I1(n17816[0]), .I2(n168_adj_5292), 
            .I3(n50700), .O(n17308[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6050_22 (.CI(n49781), .I0(n13171[19]), .I1(GND_net), 
            .CO(n49782));
    SB_LUT4 unary_minus_26_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n57[23]), 
            .I3(n49379), .O(n432[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6050_21_lut (.I0(GND_net), .I1(n13171[18]), .I2(GND_net), 
            .I3(n49780), .O(n12109[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6323_3 (.CI(n50700), .I0(n17816[0]), .I1(n168_adj_5292), 
            .CO(n50701));
    SB_LUT4 add_6323_2_lut (.I0(GND_net), .I1(n26_adj_5293), .I2(n95_adj_5294), 
            .I3(GND_net), .O(n17308[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6323_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[14]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n1050_adj_5296));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i706_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6050_21 (.CI(n49780), .I0(n13171[18]), .I1(GND_net), 
            .CO(n49781));
    SB_LUT4 unary_minus_26_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[15]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6323_2 (.CI(GND_net), .I0(n26_adj_5293), .I1(n95_adj_5294), 
            .CO(n50700));
    SB_LUT4 unary_minus_26_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n57[22]), 
            .I3(n49378), .O(n432[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i81_2_lut (.I0(\Kp[1] ), .I1(n55[19]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_5298));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6353_16_lut (.I0(GND_net), .I1(n18262[13]), .I2(n1120_adj_5299), 
            .I3(n50699), .O(n17816[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i34_2_lut (.I0(\Kp[0] ), .I1(n55[20]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6353_15_lut (.I0(GND_net), .I1(n18262[12]), .I2(n1047_adj_5300), 
            .I3(n50698), .O(n17816[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_15 (.CI(n50698), .I0(n18262[12]), .I1(n1047_adj_5300), 
            .CO(n50699));
    SB_LUT4 mult_16_i151_2_lut (.I0(\Kp[3] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_5301));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i151_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_26_add_3_24 (.CI(n49378), .I0(GND_net), .I1(n57[22]), 
            .CO(n49379));
    SB_LUT4 add_6353_14_lut (.I0(GND_net), .I1(n18262[11]), .I2(n974_adj_5302), 
            .I3(n50697), .O(n17816[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_14 (.CI(n50697), .I0(n18262[11]), .I1(n974_adj_5302), 
            .CO(n50698));
    SB_LUT4 add_6050_20_lut (.I0(GND_net), .I1(n13171[17]), .I2(GND_net), 
            .I3(n49779), .O(n12109[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6050_20 (.CI(n49779), .I0(n13171[17]), .I1(GND_net), 
            .CO(n49780));
    SB_LUT4 add_6050_19_lut (.I0(GND_net), .I1(n13171[16]), .I2(GND_net), 
            .I3(n49778), .O(n12109[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6050_19 (.CI(n49778), .I0(n13171[16]), .I1(GND_net), 
            .CO(n49779));
    SB_LUT4 add_6353_13_lut (.I0(GND_net), .I1(n18262[10]), .I2(n901_adj_5303), 
            .I3(n50696), .O(n17816[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_13 (.CI(n50696), .I0(n18262[10]), .I1(n901_adj_5303), 
            .CO(n50697));
    SB_LUT4 add_6050_18_lut (.I0(GND_net), .I1(n13171[15]), .I2(GND_net), 
            .I3(n49777), .O(n12109[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6353_12_lut (.I0(GND_net), .I1(n18262[9]), .I2(n828_adj_5304), 
            .I3(n50695), .O(n17816[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_12 (.CI(n50695), .I0(n18262[9]), .I1(n828_adj_5304), 
            .CO(n50696));
    SB_LUT4 add_6353_11_lut (.I0(GND_net), .I1(n18262[8]), .I2(n755_adj_5305), 
            .I3(n50694), .O(n17816[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n57[21]), 
            .I3(n49377), .O(n432[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6050_18 (.CI(n49777), .I0(n13171[15]), .I1(GND_net), 
            .CO(n49778));
    SB_CARRY unary_minus_26_add_3_23 (.CI(n49377), .I0(GND_net), .I1(n57[21]), 
            .CO(n49378));
    SB_LUT4 add_6050_17_lut (.I0(GND_net), .I1(n13171[14]), .I2(GND_net), 
            .I3(n49776), .O(n12109[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_11 (.CI(n50694), .I0(n18262[8]), .I1(n755_adj_5305), 
            .CO(n50695));
    SB_LUT4 add_6353_10_lut (.I0(GND_net), .I1(n18262[7]), .I2(n682_adj_5307), 
            .I3(n50693), .O(n17816[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n57[20]), 
            .I3(n49376), .O(n432[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_10 (.CI(n50693), .I0(n18262[7]), .I1(n682_adj_5307), 
            .CO(n50694));
    SB_LUT4 mult_16_i200_2_lut (.I0(\Kp[4] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_5309));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i200_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6050_17 (.CI(n49776), .I0(n13171[14]), .I1(GND_net), 
            .CO(n49777));
    SB_LUT4 mult_16_i130_2_lut (.I0(\Kp[2] ), .I1(n55[19]), .I2(GND_net), 
            .I3(GND_net), .O(n192));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6050_16_lut (.I0(GND_net), .I1(n13171[13]), .I2(n1099_adj_5310), 
            .I3(n49775), .O(n12109[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6353_9_lut (.I0(GND_net), .I1(n18262[6]), .I2(n609_adj_5311), 
            .I3(n50692), .O(n17816[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i179_2_lut (.I0(\Kp[3] ), .I1(n55[19]), .I2(GND_net), 
            .I3(GND_net), .O(n265));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i179_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6353_9 (.CI(n50692), .I0(n18262[6]), .I1(n609_adj_5311), 
            .CO(n50693));
    SB_CARRY unary_minus_26_add_3_22 (.CI(n49376), .I0(GND_net), .I1(n57[20]), 
            .CO(n49377));
    SB_CARRY add_6050_16 (.CI(n49775), .I0(n13171[13]), .I1(n1099_adj_5310), 
            .CO(n49776));
    SB_LUT4 unary_minus_26_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n57[19]), 
            .I3(n49375), .O(n432[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_21 (.CI(n49375), .I0(GND_net), .I1(n57[19]), 
            .CO(n49376));
    SB_LUT4 add_6050_15_lut (.I0(GND_net), .I1(n13171[12]), .I2(n1026_adj_5313), 
            .I3(n49774), .O(n12109[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6050_15 (.CI(n49774), .I0(n13171[12]), .I1(n1026_adj_5313), 
            .CO(n49775));
    SB_LUT4 add_6050_14_lut (.I0(GND_net), .I1(n13171[11]), .I2(n953_adj_5314), 
            .I3(n49773), .O(n12109[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6050_14 (.CI(n49773), .I0(n13171[11]), .I1(n953_adj_5314), 
            .CO(n49774));
    SB_LUT4 unary_minus_26_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n57[18]), 
            .I3(n49374), .O(n432[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_20 (.CI(n49374), .I0(GND_net), .I1(n57[18]), 
            .CO(n49375));
    SB_LUT4 add_6353_8_lut (.I0(GND_net), .I1(n18262[5]), .I2(n536_adj_5315), 
            .I3(n50691), .O(n17816[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[16]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6050_13_lut (.I0(GND_net), .I1(n13171[10]), .I2(n880_adj_5317), 
            .I3(n49772), .O(n12109[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6050_13 (.CI(n49772), .I0(n13171[10]), .I1(n880_adj_5317), 
            .CO(n49773));
    SB_LUT4 mult_16_i228_2_lut (.I0(\Kp[4] ), .I1(n55[19]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_5318));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6050_12_lut (.I0(GND_net), .I1(n13171[9]), .I2(n807_adj_5319), 
            .I3(n49771), .O(n12109[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_8 (.CI(n50691), .I0(n18262[5]), .I1(n536_adj_5315), 
            .CO(n50692));
    SB_LUT4 add_6353_7_lut (.I0(GND_net), .I1(n18262[4]), .I2(n463_adj_5320), 
            .I3(n50690), .O(n17816[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i249_2_lut (.I0(\Kp[5] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_5321));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i298_2_lut (.I0(\Kp[6] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_5322));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i298_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6050_12 (.CI(n49771), .I0(n13171[9]), .I1(n807_adj_5319), 
            .CO(n49772));
    SB_LUT4 add_6050_11_lut (.I0(GND_net), .I1(n13171[8]), .I2(n734_adj_5323), 
            .I3(n49770), .O(n12109[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_7 (.CI(n50690), .I0(n18262[4]), .I1(n463_adj_5320), 
            .CO(n50691));
    SB_CARRY add_6050_11 (.CI(n49770), .I0(n13171[8]), .I1(n734_adj_5323), 
            .CO(n49771));
    SB_LUT4 add_6050_10_lut (.I0(GND_net), .I1(n13171[7]), .I2(n661_adj_5324), 
            .I3(n49769), .O(n12109[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6050_10 (.CI(n49769), .I0(n13171[7]), .I1(n661_adj_5324), 
            .CO(n49770));
    SB_LUT4 add_6353_6_lut (.I0(GND_net), .I1(n18262[3]), .I2(n390_adj_5325), 
            .I3(n50689), .O(n17816[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_6 (.CI(n50689), .I0(n18262[3]), .I1(n390_adj_5325), 
            .CO(n50690));
    SB_LUT4 add_6353_5_lut (.I0(GND_net), .I1(n18262[2]), .I2(n317_adj_5326), 
            .I3(n50688), .O(n17816[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_5 (.CI(n50688), .I0(n18262[2]), .I1(n317_adj_5326), 
            .CO(n50689));
    SB_LUT4 add_6353_4_lut (.I0(GND_net), .I1(n18262[1]), .I2(n244_adj_5327), 
            .I3(n50687), .O(n17816[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_4 (.CI(n50687), .I0(n18262[1]), .I1(n244_adj_5327), 
            .CO(n50688));
    SB_LUT4 mult_16_i277_2_lut (.I0(\Kp[5] ), .I1(n55[19]), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i326_2_lut (.I0(\Kp[6] ), .I1(n55[19]), .I2(GND_net), 
            .I3(GND_net), .O(n484));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i347_2_lut (.I0(\Kp[7] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_5328));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i375_2_lut (.I0(\Kp[7] ), .I1(n55[19]), .I2(GND_net), 
            .I3(GND_net), .O(n557));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6050_9_lut (.I0(GND_net), .I1(n13171[6]), .I2(n588_adj_5329), 
            .I3(n49768), .O(n12109[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6353_3_lut (.I0(GND_net), .I1(n18262[0]), .I2(n171_adj_5330), 
            .I3(n50686), .O(n17816[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6353_3 (.CI(n50686), .I0(n18262[0]), .I1(n171_adj_5330), 
            .CO(n50687));
    SB_LUT4 mult_16_i424_2_lut (.I0(\Kp[8] ), .I1(n55[19]), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n57[17]), 
            .I3(n49373), .O(n432[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6353_2_lut (.I0(GND_net), .I1(n29_adj_5332), .I2(n98_adj_5333), 
            .I3(GND_net), .O(n17816[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6353_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i10_3_lut (.I0(n130[9]), .I1(n182[9]), .I2(n181), .I3(GND_net), 
            .O(n207[9]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6353_2 (.CI(GND_net), .I0(n29_adj_5332), .I1(n98_adj_5333), 
            .CO(n50686));
    SB_CARRY add_6050_9 (.CI(n49768), .I0(n13171[6]), .I1(n588_adj_5329), 
            .CO(n49769));
    SB_CARRY add_9_5 (.CI(n49220), .I0(\PID_CONTROLLER.integral [3]), .I1(n55[7]), 
            .CO(n49221));
    SB_CARRY unary_minus_26_add_3_19 (.CI(n49373), .I0(GND_net), .I1(n57[17]), 
            .CO(n49374));
    SB_LUT4 add_6497_9_lut (.I0(GND_net), .I1(n19906[6]), .I2(n630), .I3(n50685), 
            .O(n19763[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6497_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6497_8_lut (.I0(GND_net), .I1(n19906[5]), .I2(n557), .I3(n50684), 
            .O(n19763[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6497_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6050_8_lut (.I0(GND_net), .I1(n13171[5]), .I2(n515_adj_5328), 
            .I3(n49767), .O(n12109[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6497_8 (.CI(n50684), .I0(n19906[5]), .I1(n557), .CO(n50685));
    SB_LUT4 add_6497_7_lut (.I0(GND_net), .I1(n19906[4]), .I2(n484), .I3(n50683), 
            .O(n19763[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6497_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i10_3_lut (.I0(n207[9]), .I1(IntegralLimit[9]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[9] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6050_8 (.CI(n49767), .I0(n13171[5]), .I1(n515_adj_5328), 
            .CO(n49768));
    SB_CARRY add_6497_7 (.CI(n50683), .I0(n19906[4]), .I1(n484), .CO(n50684));
    SB_LUT4 add_6497_6_lut (.I0(GND_net), .I1(n19906[3]), .I2(n411), .I3(n50682), 
            .O(n19763[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6497_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6050_7_lut (.I0(GND_net), .I1(n13171[4]), .I2(n442_adj_5322), 
            .I3(n49766), .O(n12109[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6050_7 (.CI(n49766), .I0(n13171[4]), .I1(n442_adj_5322), 
            .CO(n49767));
    SB_CARRY add_6497_6 (.CI(n50682), .I0(n19906[3]), .I1(n411), .CO(n50683));
    SB_LUT4 mult_17_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_5333));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6050_6_lut (.I0(GND_net), .I1(n13171[3]), .I2(n369_adj_5321), 
            .I3(n49765), .O(n12109[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6050_6 (.CI(n49765), .I0(n13171[3]), .I1(n369_adj_5321), 
            .CO(n49766));
    SB_LUT4 add_6497_5_lut (.I0(GND_net), .I1(n19906[2]), .I2(n338_adj_5318), 
            .I3(n50681), .O(n19763[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6497_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6497_5 (.CI(n50681), .I0(n19906[2]), .I1(n338_adj_5318), 
            .CO(n50682));
    SB_LUT4 unary_minus_26_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n57[16]), 
            .I3(n49372), .O(n432[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5332));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[17]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i63_2_lut (.I0(\Kp[1] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6497_4_lut (.I0(GND_net), .I1(n19906[1]), .I2(n265), .I3(n50680), 
            .O(n19763[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6497_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_5330));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i396_2_lut (.I0(\Kp[8] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_5329));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i16_2_lut (.I0(\Kp[0] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5128));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_9_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n55[6]), .I3(n49219), .O(n130[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6497_4 (.CI(n50680), .I0(n19906[1]), .I1(n265), .CO(n50681));
    SB_LUT4 add_6497_3_lut (.I0(GND_net), .I1(n19906[0]), .I2(n192), .I3(n50679), 
            .O(n19763[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6497_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6050_5_lut (.I0(GND_net), .I1(n13171[2]), .I2(n296_adj_5309), 
            .I3(n49764), .O(n12109[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6050_5 (.CI(n49764), .I0(n13171[2]), .I1(n296_adj_5309), 
            .CO(n49765));
    SB_CARRY add_6497_3 (.CI(n50679), .I0(n19906[0]), .I1(n192), .CO(n50680));
    SB_LUT4 add_6050_4_lut (.I0(GND_net), .I1(n13171[1]), .I2(n223_adj_5301), 
            .I3(n49763), .O(n12109[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6050_4 (.CI(n49763), .I0(n13171[1]), .I1(n223_adj_5301), 
            .CO(n49764));
    SB_LUT4 add_6497_2_lut (.I0(GND_net), .I1(n50), .I2(n119_adj_5298), 
            .I3(GND_net), .O(n19763[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6497_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6497_2 (.CI(GND_net), .I0(n50), .I1(n119_adj_5298), .CO(n50679));
    SB_CARRY unary_minus_26_add_3_18 (.CI(n49372), .I0(GND_net), .I1(n57[16]), 
            .CO(n49373));
    SB_LUT4 unary_minus_26_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n57[15]), 
            .I3(n49371), .O(n432[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_9_4 (.CI(n49219), .I0(\PID_CONTROLLER.integral [2]), .I1(n55[6]), 
            .CO(n49220));
    SB_LUT4 add_6381_15_lut (.I0(GND_net), .I1(n18650[12]), .I2(n1050_adj_5296), 
            .I3(n50678), .O(n18262[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_17 (.CI(n49371), .I0(GND_net), .I1(n57[15]), 
            .CO(n49372));
    SB_LUT4 unary_minus_26_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n57[14]), 
            .I3(n49370), .O(n432[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6381_14_lut (.I0(GND_net), .I1(n18650[11]), .I2(n977_adj_5290), 
            .I3(n50677), .O(n18262[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_14 (.CI(n50677), .I0(n18650[11]), .I1(n977_adj_5290), 
            .CO(n50678));
    SB_LUT4 add_6365_15_lut (.I0(GND_net), .I1(n18428[12]), .I2(n1050), 
            .I3(n49513), .O(n18009[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6365_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n55[5]), .I3(n49218), .O(n130[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6381_13_lut (.I0(GND_net), .I1(n18650[10]), .I2(n904_adj_5285), 
            .I3(n50676), .O(n18262[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6050_3_lut (.I0(GND_net), .I1(n13171[0]), .I2(n150_adj_5275), 
            .I3(n49762), .O(n12109[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6050_3 (.CI(n49762), .I0(n13171[0]), .I1(n150_adj_5275), 
            .CO(n49763));
    SB_CARRY add_6381_13 (.CI(n50676), .I0(n18650[10]), .I1(n904_adj_5285), 
            .CO(n50677));
    SB_CARRY add_9_3 (.CI(n49218), .I0(\PID_CONTROLLER.integral [1]), .I1(n55[5]), 
            .CO(n49219));
    SB_LUT4 add_6381_12_lut (.I0(GND_net), .I1(n18650[9]), .I2(n831_adj_5270), 
            .I3(n50675), .O(n18262[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_5327));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i41_2_lut (.I0(IntegralLimit[20]), .I1(n130[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5335));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6381_12 (.CI(n50675), .I0(n18650[9]), .I1(n831_adj_5270), 
            .CO(n50676));
    SB_LUT4 mult_17_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n317_adj_5326));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6381_11_lut (.I0(GND_net), .I1(n18650[8]), .I2(n758_adj_5267), 
            .I3(n50674), .O(n18262[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_5325));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6050_2_lut (.I0(GND_net), .I1(n8_adj_5265), .I2(n77_adj_5254), 
            .I3(GND_net), .O(n12109[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6050_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_11 (.CI(n50674), .I0(n18650[8]), .I1(n758_adj_5267), 
            .CO(n50675));
    SB_CARRY add_6050_2 (.CI(GND_net), .I0(n8_adj_5265), .I1(n77_adj_5254), 
            .CO(n49762));
    SB_LUT4 add_6381_10_lut (.I0(GND_net), .I1(n18650[7]), .I2(n685_adj_5239), 
            .I3(n50673), .O(n18262[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_9_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n55[4]), .I3(GND_net), .O(n130[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_9_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6365_14_lut (.I0(GND_net), .I1(n18428[11]), .I2(n977), 
            .I3(n49512), .O(n18009[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6365_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6365_14 (.CI(n49512), .I0(n18428[11]), .I1(n977), .CO(n49513));
    SB_CARRY add_9_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), .I1(n55[4]), 
            .CO(n49218));
    SB_LUT4 add_6365_13_lut (.I0(GND_net), .I1(n18428[10]), .I2(n904), 
            .I3(n49511), .O(n18009[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6365_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_10 (.CI(n50673), .I0(n18650[7]), .I1(n685_adj_5239), 
            .CO(n50674));
    SB_LUT4 add_6381_9_lut (.I0(GND_net), .I1(n18650[6]), .I2(n612_adj_5230), 
            .I3(n50672), .O(n18262[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6365_13 (.CI(n49511), .I0(n18428[10]), .I1(n904), .CO(n49512));
    SB_CARRY add_6381_9 (.CI(n50672), .I0(n18650[6]), .I1(n612_adj_5230), 
            .CO(n50673));
    SB_CARRY unary_minus_26_add_3_16 (.CI(n49370), .I0(GND_net), .I1(n57[14]), 
            .CO(n49371));
    SB_LUT4 add_6381_8_lut (.I0(GND_net), .I1(n18650[5]), .I2(n539_adj_5227), 
            .I3(n50671), .O(n18262[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i445_2_lut (.I0(\Kp[9] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_5324));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i494_2_lut (.I0(\Kp[10] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_5323));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_5320));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i543_2_lut (.I0(\Kp[11] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n807_adj_5319));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i592_2_lut (.I0(\Kp[12] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_5317));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i592_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6381_8 (.CI(n50671), .I0(n18650[5]), .I1(n539_adj_5227), 
            .CO(n50672));
    SB_LUT4 add_6365_12_lut (.I0(GND_net), .I1(n18428[9]), .I2(n831), 
            .I3(n49510), .O(n18009[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6365_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6381_7_lut (.I0(GND_net), .I1(n18650[4]), .I2(n466_adj_5219), 
            .I3(n50670), .O(n18262[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_7 (.CI(n50670), .I0(n18650[4]), .I1(n466_adj_5219), 
            .CO(n50671));
    SB_LUT4 mult_17_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n536_adj_5315));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[18]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6365_12 (.CI(n49510), .I0(n18428[9]), .I1(n831), .CO(n49511));
    SB_LUT4 add_6381_6_lut (.I0(GND_net), .I1(n18650[3]), .I2(n393_adj_5216), 
            .I3(n50669), .O(n18262[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n57[13]), 
            .I3(n49369), .O(n432[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_6 (.CI(n50669), .I0(n18650[3]), .I1(n393_adj_5216), 
            .CO(n50670));
    SB_LUT4 sub_8_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(\motor_state[23] ), 
            .I3(n49217), .O(n55[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6365_11_lut (.I0(GND_net), .I1(n18428[8]), .I2(n758), 
            .I3(n49509), .O(n18009[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6365_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6381_5_lut (.I0(GND_net), .I1(n18650[2]), .I2(n320_adj_5183), 
            .I3(n50668), .O(n18262[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_5 (.CI(n50668), .I0(n18650[2]), .I1(n320_adj_5183), 
            .CO(n50669));
    SB_LUT4 add_6381_4_lut (.I0(GND_net), .I1(n18650[1]), .I2(n247_adj_5182), 
            .I3(n50667), .O(n18262[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_4 (.CI(n50667), .I0(n18650[1]), .I1(n247_adj_5182), 
            .CO(n50668));
    SB_LUT4 mult_16_i641_2_lut (.I0(\Kp[13] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_5314));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i39_2_lut (.I0(IntegralLimit[19]), .I1(n130[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5336));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6381_3_lut (.I0(GND_net), .I1(n18650[0]), .I2(n174_adj_5181), 
            .I3(n50666), .O(n18262[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i690_2_lut (.I0(\Kp[14] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_5313));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[19]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6381_3 (.CI(n50666), .I0(n18650[0]), .I1(n174_adj_5181), 
            .CO(n50667));
    SB_LUT4 add_6381_2_lut (.I0(GND_net), .I1(n32_adj_5180), .I2(n101_adj_5179), 
            .I3(GND_net), .O(n18262[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6381_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n609_adj_5311));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_8_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(\motor_state[22] ), 
            .I3(n49216), .O(n55[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6381_2 (.CI(GND_net), .I0(n32_adj_5180), .I1(n101_adj_5179), 
            .CO(n50666));
    SB_LUT4 add_6407_14_lut (.I0(GND_net), .I1(n18984[11]), .I2(n980), 
            .I3(n50665), .O(n18650[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6407_13_lut (.I0(GND_net), .I1(n18984[10]), .I2(n907), 
            .I3(n50664), .O(n18650[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_13 (.CI(n50664), .I0(n18984[10]), .I1(n907), .CO(n50665));
    SB_LUT4 add_6407_12_lut (.I0(GND_net), .I1(n18984[9]), .I2(n834), 
            .I3(n50663), .O(n18650[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_12 (.CI(n50663), .I0(n18984[9]), .I1(n834), .CO(n50664));
    SB_CARRY add_6365_11 (.CI(n49509), .I0(n18428[8]), .I1(n758), .CO(n49510));
    SB_LUT4 add_6407_11_lut (.I0(GND_net), .I1(n18984[8]), .I2(n761), 
            .I3(n50662), .O(n18650[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_11 (.CI(n50662), .I0(n18984[8]), .I1(n761), .CO(n50663));
    SB_LUT4 add_6407_10_lut (.I0(GND_net), .I1(n18984[7]), .I2(n688), 
            .I3(n50661), .O(n18650[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_10 (.CI(n50661), .I0(n18984[7]), .I1(n688), .CO(n50662));
    SB_LUT4 add_6407_9_lut (.I0(GND_net), .I1(n18984[6]), .I2(n615), .I3(n50660), 
            .O(n18650[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_9 (.CI(n50660), .I0(n18984[6]), .I1(n615), .CO(n50661));
    SB_LUT4 mult_16_i739_2_lut (.I0(\Kp[15] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_5310));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[20]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n682_adj_5307));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[21]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n755_adj_5305));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n828_adj_5304));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6407_8_lut (.I0(GND_net), .I1(n18984[5]), .I2(n542), .I3(n50659), 
            .O(n18650[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_8 (.CI(n50659), .I0(n18984[5]), .I1(n542), .CO(n50660));
    SB_LUT4 add_6407_7_lut (.I0(GND_net), .I1(n18984[4]), .I2(n469), .I3(n50658), 
            .O(n18650[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_7 (.CI(n50658), .I0(n18984[4]), .I1(n469), .CO(n50659));
    SB_LUT4 add_6407_6_lut (.I0(GND_net), .I1(n18984[3]), .I2(n396), .I3(n50657), 
            .O(n18650[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n901_adj_5303));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i606_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_8_add_2_24 (.CI(n49216), .I0(setpoint[22]), .I1(\motor_state[22] ), 
            .CO(n49217));
    SB_CARRY add_6407_6 (.CI(n50657), .I0(n18984[3]), .I1(n396), .CO(n50658));
    SB_LUT4 add_6407_5_lut (.I0(GND_net), .I1(n18984[2]), .I2(n323), .I3(n50656), 
            .O(n18650[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_5 (.CI(n50656), .I0(n18984[2]), .I1(n323), .CO(n50657));
    SB_LUT4 add_6407_4_lut (.I0(GND_net), .I1(n18984[1]), .I2(n250), .I3(n50655), 
            .O(n18650[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_4 (.CI(n50655), .I0(n18984[1]), .I1(n250), .CO(n50656));
    SB_LUT4 add_6407_3_lut (.I0(GND_net), .I1(n18984[0]), .I2(n177), .I3(n50654), 
            .O(n18650[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6407_3 (.CI(n50654), .I0(n18984[0]), .I1(n177), .CO(n50655));
    SB_LUT4 add_6407_2_lut (.I0(GND_net), .I1(n35_adj_5171), .I2(n104), 
            .I3(GND_net), .O(n18650[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6407_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i45_2_lut (.I0(IntegralLimit[22]), .I1(n130[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5337));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i45_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6407_2 (.CI(GND_net), .I0(n35_adj_5171), .I1(n104), .CO(n50654));
    SB_LUT4 mult_17_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n974_adj_5302));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6512_8_lut (.I0(GND_net), .I1(n20017[5]), .I2(n560_adj_5168), 
            .I3(n50653), .O(n19906[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6512_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6512_7_lut (.I0(GND_net), .I1(n20017[4]), .I2(n487_adj_5167), 
            .I3(n50652), .O(n19906[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6512_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(\motor_state[21] ), 
            .I3(n49215), .O(n55[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6512_7 (.CI(n50652), .I0(n20017[4]), .I1(n487_adj_5167), 
            .CO(n50653));
    SB_LUT4 add_6365_10_lut (.I0(GND_net), .I1(n18428[7]), .I2(n685), 
            .I3(n49508), .O(n18009[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6365_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6365_10 (.CI(n49508), .I0(n18428[7]), .I1(n685), .CO(n49509));
    SB_LUT4 add_6512_6_lut (.I0(GND_net), .I1(n20017[3]), .I2(n414_adj_5163), 
            .I3(n50651), .O(n19906[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6512_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6512_6 (.CI(n50651), .I0(n20017[3]), .I1(n414_adj_5163), 
            .CO(n50652));
    SB_LUT4 mult_17_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n1047_adj_5300));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i43_2_lut (.I0(IntegralLimit[21]), .I1(n130[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5338));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n1120_adj_5299));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6512_5_lut (.I0(GND_net), .I1(n20017[2]), .I2(n341_adj_5162), 
            .I3(n50650), .O(n19906[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6512_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[22]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_14_i9_3_lut (.I0(n130[8]), .I1(n182[8]), .I2(n181), .I3(GND_net), 
            .O(n207[8]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6512_5 (.CI(n50650), .I0(n20017[2]), .I1(n341_adj_5162), 
            .CO(n50651));
    SB_LUT4 add_6512_4_lut (.I0(GND_net), .I1(n20017[1]), .I2(n268_adj_5161), 
            .I3(n50649), .O(n19906[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6512_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6512_4 (.CI(n50649), .I0(n20017[1]), .I1(n268_adj_5161), 
            .CO(n50650));
    SB_LUT4 mux_15_i9_3_lut (.I0(n207[8]), .I1(IntegralLimit[8]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[8] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6512_3_lut (.I0(GND_net), .I1(n20017[0]), .I2(n195), .I3(n50648), 
            .O(n19906[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6512_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6512_3 (.CI(n50648), .I0(n20017[0]), .I1(n195), .CO(n50649));
    SB_LUT4 mult_17_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_5294));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6512_2_lut (.I0(GND_net), .I1(n53_c), .I2(n122_adj_5154), 
            .I3(GND_net), .O(n19906[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6512_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6512_2 (.CI(GND_net), .I0(n53_c), .I1(n122_adj_5154), 
            .CO(n50648));
    SB_LUT4 add_6431_13_lut (.I0(GND_net), .I1(n19268[10]), .I2(n910), 
            .I3(n50647), .O(n18984[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_15 (.CI(n49369), .I0(GND_net), .I1(n57[13]), 
            .CO(n49370));
    SB_LUT4 add_6431_12_lut (.I0(GND_net), .I1(n19268[9]), .I2(n837), 
            .I3(n50646), .O(n18984[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_12 (.CI(n50646), .I0(n19268[9]), .I1(n837), .CO(n50647));
    SB_LUT4 add_6431_11_lut (.I0(GND_net), .I1(n19268[8]), .I2(n764), 
            .I3(n50645), .O(n18984[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_11 (.CI(n50645), .I0(n19268[8]), .I1(n764), .CO(n50646));
    SB_LUT4 add_6431_10_lut (.I0(GND_net), .I1(n19268[7]), .I2(n691), 
            .I3(n50644), .O(n18984[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_10 (.CI(n50644), .I0(n19268[7]), .I1(n691), .CO(n50645));
    SB_LUT4 add_6431_9_lut (.I0(GND_net), .I1(n19268[6]), .I2(n618), .I3(n50643), 
            .O(n18984[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_5293));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[23]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6431_9 (.CI(n50643), .I0(n19268[6]), .I1(n618), .CO(n50644));
    SB_LUT4 add_6431_8_lut (.I0(GND_net), .I1(n19268[5]), .I2(n545), .I3(n50642), 
            .O(n18984[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_8 (.CI(n50642), .I0(n19268[5]), .I1(n545), .CO(n50643));
    SB_LUT4 add_6431_7_lut (.I0(GND_net), .I1(n19268[4]), .I2(n472), .I3(n50641), 
            .O(n18984[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_7 (.CI(n50641), .I0(n19268[4]), .I1(n472), .CO(n50642));
    SB_LUT4 add_6431_6_lut (.I0(GND_net), .I1(n19268[3]), .I2(n399), .I3(n50640), 
            .O(n18984[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_6 (.CI(n50640), .I0(n19268[3]), .I1(n399), .CO(n50641));
    SB_LUT4 add_6431_5_lut (.I0(GND_net), .I1(n19268[2]), .I2(n326), .I3(n50639), 
            .O(n18984[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_5 (.CI(n50639), .I0(n19268[2]), .I1(n326), .CO(n50640));
    SB_LUT4 add_6365_9_lut (.I0(GND_net), .I1(n18428[6]), .I2(n612), .I3(n49507), 
            .O(n18009[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6365_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6431_4_lut (.I0(GND_net), .I1(n19268[1]), .I2(n253), .I3(n50638), 
            .O(n18984[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_4 (.CI(n50638), .I0(n19268[1]), .I1(n253), .CO(n50639));
    SB_LUT4 add_6431_3_lut (.I0(GND_net), .I1(n19268[0]), .I2(n180), .I3(n50637), 
            .O(n18984[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_3 (.CI(n50637), .I0(n19268[0]), .I1(n180), .CO(n50638));
    SB_LUT4 add_6431_2_lut (.I0(GND_net), .I1(n38), .I2(n107_adj_5139), 
            .I3(GND_net), .O(n18984[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6431_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6119_22_lut (.I0(GND_net), .I1(n14095[19]), .I2(GND_net), 
            .I3(n49744), .O(n13171[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6431_2 (.CI(GND_net), .I0(n38), .I1(n107_adj_5139), .CO(n50637));
    SB_LUT4 add_6453_12_lut (.I0(GND_net), .I1(n19506[9]), .I2(n840), 
            .I3(n50636), .O(n19268[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6453_11_lut (.I0(GND_net), .I1(n19506[8]), .I2(n767), 
            .I3(n50635), .O(n19268[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_5292));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i114_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6453_11 (.CI(n50635), .I0(n19506[8]), .I1(n767), .CO(n50636));
    SB_LUT4 LessThan_10_i37_2_lut (.I0(IntegralLimit[18]), .I1(n130[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5341));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6453_10_lut (.I0(GND_net), .I1(n19506[7]), .I2(n694), 
            .I3(n50634), .O(n19268[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6453_10 (.CI(n50634), .I0(n19506[7]), .I1(n694), .CO(n50635));
    SB_LUT4 add_6453_9_lut (.I0(GND_net), .I1(n19506[6]), .I2(n621), .I3(n50633), 
            .O(n19268[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i67_2_lut (.I0(\Kp[1] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n98));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i67_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6453_9 (.CI(n50633), .I0(n19506[6]), .I1(n621), .CO(n50634));
    SB_LUT4 mult_16_i20_2_lut (.I0(\Kp[0] ), .I1(n55[13]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5291));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6453_8_lut (.I0(GND_net), .I1(n19506[5]), .I2(n548), .I3(n50632), 
            .O(n19268[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6453_8 (.CI(n50632), .I0(n19506[5]), .I1(n548), .CO(n50633));
    SB_LUT4 add_6453_7_lut (.I0(GND_net), .I1(n19506[4]), .I2(n475), .I3(n50631), 
            .O(n19268[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6453_7 (.CI(n50631), .I0(n19506[4]), .I1(n475), .CO(n50632));
    SB_LUT4 unary_minus_26_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n57[12]), 
            .I3(n49368), .O(n432[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_5289));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6453_6_lut (.I0(GND_net), .I1(n19506[3]), .I2(n402), .I3(n50630), 
            .O(n19268[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6119_21_lut (.I0(GND_net), .I1(n14095[18]), .I2(GND_net), 
            .I3(n49743), .O(n13171[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6365_9 (.CI(n49507), .I0(n18428[6]), .I1(n612), .CO(n49508));
    SB_CARRY add_6453_6 (.CI(n50630), .I0(n19506[3]), .I1(n402), .CO(n50631));
    SB_LUT4 add_6453_5_lut (.I0(GND_net), .I1(n19506[2]), .I2(n329), .I3(n50629), 
            .O(n19268[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_14 (.CI(n49368), .I0(GND_net), .I1(n57[12]), 
            .CO(n49369));
    SB_CARRY add_6453_5 (.CI(n50629), .I0(n19506[2]), .I1(n329), .CO(n50630));
    SB_LUT4 add_6453_4_lut (.I0(GND_net), .I1(n19506[1]), .I2(n256), .I3(n50628), 
            .O(n19268[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6119_21 (.CI(n49743), .I0(n14095[18]), .I1(GND_net), 
            .CO(n49744));
    SB_CARRY add_6453_4 (.CI(n50628), .I0(n19506[1]), .I1(n256), .CO(n50629));
    SB_LUT4 add_6453_3_lut (.I0(GND_net), .I1(n19506[0]), .I2(n183_adj_5137), 
            .I3(n50627), .O(n19268[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6453_3 (.CI(n50627), .I0(n19506[0]), .I1(n183_adj_5137), 
            .CO(n50628));
    SB_LUT4 add_6453_2_lut (.I0(GND_net), .I1(n41_adj_5136), .I2(n110), 
            .I3(GND_net), .O(n19268[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6453_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6453_2 (.CI(GND_net), .I0(n41_adj_5136), .I1(n110), .CO(n50627));
    SB_LUT4 add_6525_7_lut (.I0(GND_net), .I1(n59192), .I2(n490_c), .I3(n50626), 
            .O(n20017[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6525_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6119_20_lut (.I0(GND_net), .I1(n14095[17]), .I2(GND_net), 
            .I3(n49742), .O(n13171[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_5288));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_5287));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_5286));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i116_2_lut (.I0(\Kp[2] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n171));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6525_6_lut (.I0(GND_net), .I1(n20100[3]), .I2(n417_c), 
            .I3(n50625), .O(n20017[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6525_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6365_8_lut (.I0(GND_net), .I1(n18428[5]), .I2(n539), .I3(n49506), 
            .O(n18009[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6365_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_23 (.CI(n49215), .I0(setpoint[21]), .I1(\motor_state[21] ), 
            .CO(n49216));
    SB_CARRY add_6365_8 (.CI(n49506), .I0(n18428[5]), .I1(n539), .CO(n49507));
    SB_CARRY add_6525_6 (.CI(n50625), .I0(n20100[3]), .I1(n417_c), .CO(n50626));
    SB_LUT4 add_6365_7_lut (.I0(GND_net), .I1(n18428[4]), .I2(n466), .I3(n49505), 
            .O(n18009[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6365_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6525_5_lut (.I0(GND_net), .I1(n20100[2]), .I2(n344_c), 
            .I3(n50624), .O(n20017[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6525_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n57[11]), 
            .I3(n49367), .O(n432[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_13 (.CI(n49367), .I0(GND_net), .I1(n57[11]), 
            .CO(n49368));
    SB_CARRY add_6525_5 (.CI(n50624), .I0(n20100[2]), .I1(n344_c), .CO(n50625));
    SB_CARRY add_6119_20 (.CI(n49742), .I0(n14095[17]), .I1(GND_net), 
            .CO(n49743));
    SB_LUT4 add_6525_4_lut (.I0(GND_net), .I1(n20100[1]), .I2(n271_c), 
            .I3(n50623), .O(n20017[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6525_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6365_7 (.CI(n49505), .I0(n18428[4]), .I1(n466), .CO(n49506));
    SB_CARRY add_6525_4 (.CI(n50623), .I0(n20100[1]), .I1(n271_c), .CO(n50624));
    SB_LUT4 add_6365_6_lut (.I0(GND_net), .I1(n18428[3]), .I2(n393), .I3(n49504), 
            .O(n18009[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6365_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n57[10]), 
            .I3(n49366), .O(n432[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i23_2_lut (.I0(IntegralLimit[11]), .I1(n130[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5343));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6525_3_lut (.I0(GND_net), .I1(n20100[0]), .I2(n198_c), 
            .I3(n50622), .O(n20017[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6525_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i25_2_lut (.I0(IntegralLimit[12]), .I1(n130[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5344));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_5284));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i165_2_lut (.I0(\Kp[3] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n244));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_5283));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i15_3_lut (.I0(n130[14]), .I1(n182[14]), .I2(n181), 
            .I3(GND_net), .O(n207[14]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i15_3_lut (.I0(n207[14]), .I1(IntegralLimit[14]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[14] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6525_3 (.CI(n50622), .I0(n20100[0]), .I1(n198_c), .CO(n50623));
    SB_LUT4 add_6525_2_lut (.I0(GND_net), .I1(n56_c), .I2(n125_c), .I3(GND_net), 
            .O(n20017[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6525_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6525_2 (.CI(GND_net), .I0(n56_c), .I1(n125_c), .CO(n50622));
    SB_CARRY add_6365_6 (.CI(n49504), .I0(n18428[3]), .I1(n393), .CO(n49505));
    SB_LUT4 sub_8_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(\motor_state[20] ), 
            .I3(n49214), .O(n55[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6119_19_lut (.I0(GND_net), .I1(n14095[16]), .I2(GND_net), 
            .I3(n49741), .O(n13171[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6365_5_lut (.I0(GND_net), .I1(n18428[2]), .I2(n320), .I3(n49503), 
            .O(n18009[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6365_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_12 (.CI(n49366), .I0(GND_net), .I1(n57[10]), 
            .CO(n49367));
    SB_LUT4 mult_17_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_5281));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_5280));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n679_adj_5279));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_5278));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n825_adj_5277));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n57[9]), 
            .I3(n49365), .O(n432[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n898_adj_5276));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i604_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6119_19 (.CI(n49741), .I0(n14095[16]), .I1(GND_net), 
            .CO(n49742));
    SB_CARRY unary_minus_26_add_3_11 (.CI(n49365), .I0(GND_net), .I1(n57[9]), 
            .CO(n49366));
    SB_LUT4 add_6119_18_lut (.I0(GND_net), .I1(n14095[15]), .I2(GND_net), 
            .I3(n49740), .O(n13171[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_5274));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i653_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6119_18 (.CI(n49740), .I0(n14095[15]), .I1(GND_net), 
            .CO(n49741));
    SB_LUT4 add_6119_17_lut (.I0(GND_net), .I1(n14095[14]), .I2(GND_net), 
            .I3(n49739), .O(n13171[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6119_17 (.CI(n49739), .I0(n14095[14]), .I1(GND_net), 
            .CO(n49740));
    SB_LUT4 unary_minus_26_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n57[8]), 
            .I3(n49364), .O(n432[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n1044_adj_5273));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n1117_adj_5272));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i35_2_lut (.I0(IntegralLimit[17]), .I1(n130[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5346));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i214_2_lut (.I0(\Kp[4] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n317));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i79_2_lut (.I0(\Kp[1] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_5271));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i32_2_lut (.I0(\Kp[0] ), .I1(n55[19]), .I2(GND_net), 
            .I3(GND_net), .O(n47));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i128_2_lut (.I0(\Kp[2] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n189));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_5269));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_10_i29_2_lut (.I0(IntegralLimit[14]), .I1(n130[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5347));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i177_2_lut (.I0(\Kp[3] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n262));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6119_16_lut (.I0(GND_net), .I1(n14095[13]), .I2(n1102), 
            .I3(n49738), .O(n13171[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6119_16 (.CI(n49738), .I0(n14095[13]), .I1(n1102), .CO(n49739));
    SB_CARRY add_6365_5 (.CI(n49503), .I0(n18428[2]), .I1(n320), .CO(n49504));
    SB_CARRY unary_minus_26_add_3_10 (.CI(n49364), .I0(GND_net), .I1(n57[8]), 
            .CO(n49365));
    SB_LUT4 add_6365_4_lut (.I0(GND_net), .I1(n18428[1]), .I2(n247), .I3(n49502), 
            .O(n18009[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6365_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_26_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n57[7]), 
            .I3(n49363), .O(n432[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6119_15_lut (.I0(GND_net), .I1(n14095[12]), .I2(n1029), 
            .I3(n49737), .O(n13171[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i31_2_lut (.I0(IntegralLimit[15]), .I1(n130[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5348));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_8_add_2_22 (.CI(n49214), .I0(setpoint[20]), .I1(\motor_state[20] ), 
            .CO(n49215));
    SB_CARRY add_6119_15 (.CI(n49737), .I0(n14095[12]), .I1(n1029), .CO(n49738));
    SB_CARRY unary_minus_26_add_3_9 (.CI(n49363), .I0(GND_net), .I1(n57[7]), 
            .CO(n49364));
    SB_LUT4 mult_16_i263_2_lut (.I0(\Kp[5] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n390));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i226_2_lut (.I0(\Kp[4] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_5268));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i275_2_lut (.I0(\Kp[5] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i324_2_lut (.I0(\Kp[6] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n481));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i373_2_lut (.I0(\Kp[7] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n554));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i312_2_lut (.I0(\Kp[6] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n463));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i312_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6365_4 (.CI(n49502), .I0(n18428[1]), .I1(n247), .CO(n49503));
    SB_LUT4 add_6119_14_lut (.I0(GND_net), .I1(n14095[11]), .I2(n956), 
            .I3(n49736), .O(n13171[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6119_14 (.CI(n49736), .I0(n14095[11]), .I1(n956), .CO(n49737));
    SB_LUT4 add_6119_13_lut (.I0(GND_net), .I1(n14095[10]), .I2(n883), 
            .I3(n49735), .O(n13171[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_5266));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6365_3_lut (.I0(GND_net), .I1(n18428[0]), .I2(n174), .I3(n49501), 
            .O(n18009[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6365_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6119_13 (.CI(n49735), .I0(n14095[10]), .I1(n883), .CO(n49736));
    SB_LUT4 unary_minus_26_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n57[6]), 
            .I3(n49362), .O(n432[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i422_2_lut (.I0(\Kp[8] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n627));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i361_2_lut (.I0(\Kp[7] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n536));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i361_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6365_3 (.CI(n49501), .I0(n18428[0]), .I1(n174), .CO(n49502));
    SB_LUT4 add_6119_12_lut (.I0(GND_net), .I1(n14095[9]), .I2(n810), 
            .I3(n49734), .O(n13171[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6365_2_lut (.I0(GND_net), .I1(n32_c), .I2(n101), .I3(GND_net), 
            .O(n18009[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6365_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6119_12 (.CI(n49734), .I0(n14095[9]), .I1(n810), .CO(n49735));
    SB_LUT4 add_6119_11_lut (.I0(GND_net), .I1(n14095[8]), .I2(n737), 
            .I3(n49733), .O(n13171[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6365_2 (.CI(GND_net), .I0(n32_c), .I1(n101), .CO(n49501));
    SB_CARRY add_6119_11 (.CI(n49733), .I0(n14095[8]), .I1(n737), .CO(n49734));
    SB_LUT4 add_6119_10_lut (.I0(GND_net), .I1(n14095[7]), .I2(n664), 
            .I3(n49732), .O(n13171[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(\motor_state[19] ), 
            .I3(n49213), .O(n55[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6119_10 (.CI(n49732), .I0(n14095[7]), .I1(n664), .CO(n49733));
    SB_LUT4 add_6119_9_lut (.I0(GND_net), .I1(n14095[6]), .I2(n591), .I3(n49731), 
            .O(n13171[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6119_9 (.CI(n49731), .I0(n14095[6]), .I1(n591), .CO(n49732));
    SB_LUT4 add_6119_8_lut (.I0(GND_net), .I1(n14095[5]), .I2(n518), .I3(n49730), 
            .O(n13171[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6119_8 (.CI(n49730), .I0(n14095[5]), .I1(n518), .CO(n49731));
    SB_LUT4 add_6119_7_lut (.I0(GND_net), .I1(n14095[4]), .I2(n445_adj_5126), 
            .I3(n49729), .O(n13171[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i112_2_lut (.I0(\Kp[2] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i112_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6119_7 (.CI(n49729), .I0(n14095[4]), .I1(n445_adj_5126), 
            .CO(n49730));
    SB_LUT4 add_6533_7_lut (.I0(GND_net), .I1(n59684), .I2(n490), .I3(n49500), 
            .O(n20078[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6533_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6119_6_lut (.I0(GND_net), .I1(n14095[3]), .I2(n372_adj_5122), 
            .I3(n49728), .O(n13171[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i161_2_lut (.I0(\Kp[3] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n238));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i161_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6119_6 (.CI(n49728), .I0(n14095[3]), .I1(n372_adj_5122), 
            .CO(n49729));
    SB_LUT4 add_6119_5_lut (.I0(GND_net), .I1(n14095[2]), .I2(n299), .I3(n49727), 
            .O(n13171[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i33_2_lut (.I0(IntegralLimit[16]), .I1(n130[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5350));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6119_5 (.CI(n49727), .I0(n14095[2]), .I1(n299), .CO(n49728));
    SB_LUT4 add_6533_6_lut (.I0(GND_net), .I1(n20146[3]), .I2(n417), .I3(n49499), 
            .O(n20078[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6533_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6119_4_lut (.I0(GND_net), .I1(n14095[1]), .I2(n226), .I3(n49726), 
            .O(n13171[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_21 (.CI(n49213), .I0(setpoint[19]), .I1(\motor_state[19] ), 
            .CO(n49214));
    SB_CARRY add_6119_4 (.CI(n49726), .I0(n14095[1]), .I1(n226), .CO(n49727));
    SB_LUT4 add_6119_3_lut (.I0(GND_net), .I1(n14095[0]), .I2(n153), .I3(n49725), 
            .O(n13171[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6119_3 (.CI(n49725), .I0(n14095[0]), .I1(n153), .CO(n49726));
    SB_CARRY add_6533_6 (.CI(n49499), .I0(n20146[3]), .I1(n417), .CO(n49500));
    SB_LUT4 LessThan_10_i11_2_lut (.I0(IntegralLimit[5]), .I1(n130[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5352));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6119_2_lut (.I0(GND_net), .I1(n11), .I2(n80), .I3(GND_net), 
            .O(n13171[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6119_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6119_2 (.CI(GND_net), .I0(n11), .I1(n80), .CO(n49725));
    SB_CARRY unary_minus_26_add_3_8 (.CI(n49362), .I0(GND_net), .I1(n57[6]), 
            .CO(n49363));
    SB_LUT4 unary_minus_26_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n57[5]), 
            .I3(n49361), .O(n432[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6533_5_lut (.I0(GND_net), .I1(n20149), .I2(n344), .I3(n49498), 
            .O(n20078[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6533_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_7 (.CI(n49361), .I0(GND_net), .I1(n57[5]), 
            .CO(n49362));
    SB_CARRY add_6533_5 (.CI(n49498), .I0(n20149), .I1(n344), .CO(n49499));
    SB_LUT4 unary_minus_26_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n57[4]), 
            .I3(n49360), .O(n432[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i13_2_lut (.I0(IntegralLimit[6]), .I1(n130[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5354));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6533_4_lut (.I0(GND_net), .I1(n20150), .I2(n271), .I3(n49497), 
            .O(n20078[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6533_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i15_2_lut (.I0(IntegralLimit[7]), .I1(n130[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5356));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_26_add_3_6 (.CI(n49360), .I0(GND_net), .I1(n57[4]), 
            .CO(n49361));
    SB_LUT4 mult_16_i210_2_lut (.I0(\Kp[4] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n311));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i259_2_lut (.I0(\Kp[5] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n384));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i308_2_lut (.I0(\Kp[6] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n457));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i357_2_lut (.I0(\Kp[7] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i471_2_lut (.I0(\Kp[9] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i8_3_lut (.I0(n130[7]), .I1(n182[7]), .I2(n181), .I3(GND_net), 
            .O(n207[7]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i8_3_lut (.I0(n207[7]), .I1(IntegralLimit[7]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[7] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_5264));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5263));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i410_2_lut (.I0(\Kp[8] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n609));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_5261));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_5260));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_5259));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_5258));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_5257));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i259_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6533_4 (.CI(n49497), .I0(n20150), .I1(n271), .CO(n49498));
    SB_LUT4 mult_17_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_5256));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i459_2_lut (.I0(\Kp[9] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n682));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_5255));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i406_2_lut (.I0(\Kp[8] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i455_2_lut (.I0(\Kp[9] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i455_2_lut.LUT_INIT = 16'h8888;
    SB_DFFR \PID_CONTROLLER.integral_i0_i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk16MHz), .D(n29641), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_LUT4 unary_minus_26_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n57[3]), 
            .I3(n49359), .O(n432[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i27_2_lut (.I0(IntegralLimit[13]), .I1(n130[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5357));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i9_2_lut (.I0(IntegralLimit[4]), .I1(n130[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5358));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i17_2_lut (.I0(IntegralLimit[8]), .I1(n130[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5359));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i19_2_lut (.I0(IntegralLimit[9]), .I1(n130[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5360));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_10_i21_2_lut (.I0(IntegralLimit[10]), .I1(n130[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5361));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50016_4_lut (.I0(n21_adj_5361), .I1(n19_adj_5360), .I2(n17_adj_5359), 
            .I3(n9_adj_5358), .O(n65702));
    defparam i50016_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_16_i508_2_lut (.I0(\Kp[10] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n755));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n603_adj_5253));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n676_adj_5252));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_5251));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49990_4_lut (.I0(n27_adj_5357), .I1(n15_adj_5356), .I2(n13_adj_5354), 
            .I3(n11_adj_5352), .O(n65676));
    defparam i49990_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_10_i12_3_lut (.I0(n130[7]), .I1(n130[16]), .I2(n33_adj_5350), 
            .I3(GND_net), .O(n12_adj_5362));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_5250));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n822_adj_5249));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i553_2_lut.LUT_INIT = 16'h8888;
    SB_DFFSR counter_1943__i0 (.Q(counter[0]), .C(clk16MHz), .D(n59[0]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_LUT4 mult_17_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n895_adj_5248));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i602_2_lut.LUT_INIT = 16'h8888;
    SB_DFFSR counter_1943__i31 (.Q(counter[31]), .C(clk16MHz), .D(n59[31]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i30 (.Q(counter[30]), .C(clk16MHz), .D(n59[30]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_LUT4 counter_1943_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(counter[31]), 
            .I3(n50495), .O(n59[31])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1943_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(counter[30]), 
            .I3(n50494), .O(n59[30])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR counter_1943__i29 (.Q(counter[29]), .C(clk16MHz), .D(n59[29]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i28 (.Q(counter[28]), .C(clk16MHz), .D(n59[28]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i27 (.Q(counter[27]), .C(clk16MHz), .D(n59[27]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i26 (.Q(counter[26]), .C(clk16MHz), .D(n59[26]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i25 (.Q(counter[25]), .C(clk16MHz), .D(n59[25]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i24 (.Q(counter[24]), .C(clk16MHz), .D(n59[24]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i23 (.Q(counter[23]), .C(clk16MHz), .D(n59[23]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i22 (.Q(counter[22]), .C(clk16MHz), .D(n59[22]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i21 (.Q(counter[21]), .C(clk16MHz), .D(n59[21]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i20 (.Q(counter[20]), .C(clk16MHz), .D(n59[20]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i19 (.Q(counter[19]), .C(clk16MHz), .D(n59[19]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_CARRY counter_1943_add_4_32 (.CI(n50494), .I0(GND_net), .I1(counter[30]), 
            .CO(n50495));
    SB_DFFSR counter_1943__i18 (.Q(counter[18]), .C(clk16MHz), .D(n59[18]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i17 (.Q(counter[17]), .C(clk16MHz), .D(n59[17]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i16 (.Q(counter[16]), .C(clk16MHz), .D(n59[16]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i15 (.Q(counter[15]), .C(clk16MHz), .D(n59[15]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i14 (.Q(counter[14]), .C(clk16MHz), .D(n59[14]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i13 (.Q(counter[13]), .C(clk16MHz), .D(n59[13]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i12 (.Q(counter[12]), .C(clk16MHz), .D(n59[12]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i11 (.Q(counter[11]), .C(clk16MHz), .D(n59[11]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i10 (.Q(counter[10]), .C(clk16MHz), .D(n59[10]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i9 (.Q(counter[9]), .C(clk16MHz), .D(n59[9]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i8 (.Q(counter[8]), .C(clk16MHz), .D(n59[8]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i7 (.Q(counter[7]), .C(clk16MHz), .D(n59[7]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i6 (.Q(counter[6]), .C(clk16MHz), .D(n59[6]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i5 (.Q(counter[5]), .C(clk16MHz), .D(n59[5]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i4 (.Q(counter[4]), .C(clk16MHz), .D(n59[4]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i3 (.Q(counter[3]), .C(clk16MHz), .D(n59[3]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i2 (.Q(counter[2]), .C(clk16MHz), .D(n59[2]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_DFFSR counter_1943__i1 (.Q(counter[1]), .C(clk16MHz), .D(n59[1]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(24[16:25])
    SB_LUT4 counter_1943_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(counter[29]), 
            .I3(n50493), .O(n59[29])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_31 (.CI(n50493), .I0(GND_net), .I1(counter[29]), 
            .CO(n50494));
    SB_LUT4 counter_1943_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(counter[28]), 
            .I3(n50492), .O(n59[28])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_30 (.CI(n50492), .I0(GND_net), .I1(counter[28]), 
            .CO(n50493));
    SB_LUT4 counter_1943_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(counter[27]), 
            .I3(n50491), .O(n59[27])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_29 (.CI(n50491), .I0(GND_net), .I1(counter[27]), 
            .CO(n50492));
    SB_LUT4 counter_1943_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(counter[26]), 
            .I3(n50490), .O(n59[26])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_28 (.CI(n50490), .I0(GND_net), .I1(counter[26]), 
            .CO(n50491));
    SB_LUT4 counter_1943_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(counter[25]), 
            .I3(n50489), .O(n59[25])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_27 (.CI(n50489), .I0(GND_net), .I1(counter[25]), 
            .CO(n50490));
    SB_LUT4 counter_1943_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(counter[24]), 
            .I3(n50488), .O(n59[24])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_26 (.CI(n50488), .I0(GND_net), .I1(counter[24]), 
            .CO(n50489));
    SB_LUT4 counter_1943_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(counter[23]), 
            .I3(n50487), .O(n59[23])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_25 (.CI(n50487), .I0(GND_net), .I1(counter[23]), 
            .CO(n50488));
    SB_LUT4 counter_1943_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(counter[22]), 
            .I3(n50486), .O(n59[22])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_24 (.CI(n50486), .I0(GND_net), .I1(counter[22]), 
            .CO(n50487));
    SB_LUT4 counter_1943_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(counter[21]), 
            .I3(n50485), .O(n59[21])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_23 (.CI(n50485), .I0(GND_net), .I1(counter[21]), 
            .CO(n50486));
    SB_LUT4 counter_1943_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(counter[20]), 
            .I3(n50484), .O(n59[20])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_22 (.CI(n50484), .I0(GND_net), .I1(counter[20]), 
            .CO(n50485));
    SB_LUT4 counter_1943_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(counter[19]), 
            .I3(n50483), .O(n59[19])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_21 (.CI(n50483), .I0(GND_net), .I1(counter[19]), 
            .CO(n50484));
    SB_LUT4 counter_1943_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(counter[18]), 
            .I3(n50482), .O(n59[18])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_20 (.CI(n50482), .I0(GND_net), .I1(counter[18]), 
            .CO(n50483));
    SB_LUT4 counter_1943_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(counter[17]), 
            .I3(n50481), .O(n59[17])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_19 (.CI(n50481), .I0(GND_net), .I1(counter[17]), 
            .CO(n50482));
    SB_LUT4 counter_1943_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(counter[16]), 
            .I3(n50480), .O(n59[16])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_18 (.CI(n50480), .I0(GND_net), .I1(counter[16]), 
            .CO(n50481));
    SB_LUT4 counter_1943_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(counter[15]), 
            .I3(n50479), .O(n59[15])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_17 (.CI(n50479), .I0(GND_net), .I1(counter[15]), 
            .CO(n50480));
    SB_LUT4 counter_1943_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(counter[14]), 
            .I3(n50478), .O(n59[14])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_16 (.CI(n50478), .I0(GND_net), .I1(counter[14]), 
            .CO(n50479));
    SB_LUT4 counter_1943_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(counter[13]), 
            .I3(n50477), .O(n59[13])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_15 (.CI(n50477), .I0(GND_net), .I1(counter[13]), 
            .CO(n50478));
    SB_LUT4 counter_1943_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(counter[12]), 
            .I3(n50476), .O(n59[12])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_14 (.CI(n50476), .I0(GND_net), .I1(counter[12]), 
            .CO(n50477));
    SB_LUT4 counter_1943_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(counter[11]), 
            .I3(n50475), .O(n59[11])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_13 (.CI(n50475), .I0(GND_net), .I1(counter[11]), 
            .CO(n50476));
    SB_LUT4 counter_1943_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(counter[10]), 
            .I3(n50474), .O(n59[10])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_12 (.CI(n50474), .I0(GND_net), .I1(counter[10]), 
            .CO(n50475));
    SB_LUT4 counter_1943_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(counter[9]), 
            .I3(n50473), .O(n59[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_11 (.CI(n50473), .I0(GND_net), .I1(counter[9]), 
            .CO(n50474));
    SB_LUT4 counter_1943_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(counter[8]), 
            .I3(n50472), .O(n59[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_10 (.CI(n50472), .I0(GND_net), .I1(counter[8]), 
            .CO(n50473));
    SB_LUT4 counter_1943_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(counter[7]), 
            .I3(n50471), .O(n59[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_9 (.CI(n50471), .I0(GND_net), .I1(counter[7]), 
            .CO(n50472));
    SB_LUT4 counter_1943_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(counter[6]), 
            .I3(n50470), .O(n59[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result__i23 (.Q(duty[23]), .C(clk16MHz), .E(control_update), 
            .D(n51[23]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_CARRY counter_1943_add_4_8 (.CI(n50470), .I0(GND_net), .I1(counter[6]), 
            .CO(n50471));
    SB_LUT4 add_6533_3_lut (.I0(GND_net), .I1(n20151), .I2(n198), .I3(n49496), 
            .O(n20078[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6533_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_1943_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(counter[5]), 
            .I3(n50469), .O(n59[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i10_3_lut (.I0(n130[5]), .I1(n130[6]), .I2(n13_adj_5354), 
            .I3(GND_net), .O(n10_adj_5391));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY counter_1943_add_4_7 (.CI(n50469), .I0(GND_net), .I1(counter[5]), 
            .CO(n50470));
    SB_LUT4 counter_1943_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n50468), .O(n59[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_6 (.CI(n50468), .I0(GND_net), .I1(counter[4]), 
            .CO(n50469));
    SB_LUT4 counter_1943_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n50467), .O(n59[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_5 (.CI(n50467), .I0(GND_net), .I1(counter[3]), 
            .CO(n50468));
    SB_LUT4 counter_1943_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n50466), .O(n59[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_4 (.CI(n50466), .I0(GND_net), .I1(counter[2]), 
            .CO(n50467));
    SB_LUT4 counter_1943_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n50465), .O(n59[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_10_i30_3_lut (.I0(n12_adj_5362), .I1(n130[17]), .I2(n35_adj_5346), 
            .I3(GND_net), .O(n30_adj_5392));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY counter_1943_add_4_3 (.CI(n50465), .I0(GND_net), .I1(counter[1]), 
            .CO(n50466));
    SB_LUT4 counter_1943_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n59[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1943_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1943_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n50465));
    SB_LUT4 mult_17_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n968_adj_5247));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n1041_adj_5246));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n1114_adj_5245));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i749_2_lut.LUT_INIT = 16'h8888;
    SB_DFFER result__i22 (.Q(duty[22]), .C(clk16MHz), .E(control_update), 
            .D(n51[22]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i21 (.Q(duty[21]), .C(clk16MHz), .E(control_update), 
            .D(n51[21]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i20 (.Q(duty[20]), .C(clk16MHz), .E(control_update), 
            .D(n51[20]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i19 (.Q(duty[19]), .C(clk16MHz), .E(control_update), 
            .D(n51[19]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i18 (.Q(duty[18]), .C(clk16MHz), .E(control_update), 
            .D(n51[18]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i17 (.Q(duty[17]), .C(clk16MHz), .E(control_update), 
            .D(n51[17]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i16 (.Q(duty[16]), .C(clk16MHz), .E(control_update), 
            .D(n51[16]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i15 (.Q(duty[15]), .C(clk16MHz), .E(control_update), 
            .D(n51[15]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i14 (.Q(duty[14]), .C(clk16MHz), .E(control_update), 
            .D(n51[14]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i13 (.Q(duty[13]), .C(clk16MHz), .E(control_update), 
            .D(n51[13]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_CARRY add_6533_3 (.CI(n49496), .I0(n20151), .I1(n198), .CO(n49497));
    SB_DFFER result__i12 (.Q(duty[12]), .C(clk16MHz), .E(control_update), 
            .D(n51[12]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i11 (.Q(duty[11]), .C(clk16MHz), .E(control_update), 
            .D(n51[11]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i10 (.Q(duty[10]), .C(clk16MHz), .E(control_update), 
            .D(n51[10]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_LUT4 add_6533_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n20078[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6533_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result__i9 (.Q(duty[9]), .C(clk16MHz), .E(control_update), 
            .D(n51[9]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i8 (.Q(duty[8]), .C(clk16MHz), .E(control_update), 
            .D(n51[8]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i7 (.Q(duty[7]), .C(clk16MHz), .E(control_update), 
            .D(n51[7]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i6 (.Q(duty[6]), .C(clk16MHz), .E(control_update), 
            .D(n51[6]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i5 (.Q(duty[5]), .C(clk16MHz), .E(control_update), 
            .D(n51[5]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i4 (.Q(duty[4]), .C(clk16MHz), .E(control_update), 
            .D(n51[4]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i3 (.Q(duty[3]), .C(clk16MHz), .E(control_update), 
            .D(n51[3]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i2 (.Q(duty[2]), .C(clk16MHz), .E(control_update), 
            .D(n51[2]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFER result__i1 (.Q(duty[1]), .C(clk16MHz), .E(control_update), 
            .D(n51[1]), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk16MHz), .D(n30463), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk16MHz), .D(n30462), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk16MHz), .D(n30461), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk16MHz), .D(n30460), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk16MHz), .D(n30459), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk16MHz), .D(n30458), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk16MHz), .D(n30457), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk16MHz), .D(n30456), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk16MHz), .D(n30455), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk16MHz), .D(n30454), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk16MHz), .D(n30453), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk16MHz), .D(n30452), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk16MHz), .D(n30451), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk16MHz), .D(n30450), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk16MHz), .D(n30449), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk16MHz), .D(n30448), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk16MHz), .D(n30447), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk16MHz), .D(n30445), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk16MHz), .D(n30443), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk16MHz), .D(n30442), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk16MHz), .D(n30441), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk16MHz), .D(n30440), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk16MHz), .D(n30439), .R(reset));   // verilog/motorControl.v(41[14] 62[8])
    SB_CARRY add_6533_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n49496));
    SB_LUT4 sub_8_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(\motor_state[18] ), 
            .I3(n49212), .O(n55[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_5 (.CI(n49359), .I0(GND_net), .I1(n57[3]), 
            .CO(n49360));
    SB_LUT4 i50725_2_lut_4_lut (.I0(n130[21]), .I1(n182[21]), .I2(n130[9]), 
            .I3(n182[9]), .O(n66411));
    defparam i50725_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 unary_minus_26_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n57[2]), 
            .I3(n49358), .O(n432[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_14_i7_3_lut (.I0(n130[6]), .I1(n182[6]), .I2(n181), .I3(GND_net), 
            .O(n207[6]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_26_add_3_4 (.CI(n49358), .I0(GND_net), .I1(n57[2]), 
            .CO(n49359));
    SB_LUT4 mux_15_i7_3_lut (.I0(n207[6]), .I1(IntegralLimit[6]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[6] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5244));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50955_4_lut (.I0(n13_adj_5354), .I1(n11_adj_5352), .I2(n9_adj_5358), 
            .I3(n65738), .O(n66641));
    defparam i50955_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50945_4_lut (.I0(n19_adj_5360), .I1(n17_adj_5359), .I2(n15_adj_5356), 
            .I3(n66641), .O(n66631));
    defparam i50945_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52226_4_lut (.I0(n25_adj_5344), .I1(n23_adj_5343), .I2(n21_adj_5361), 
            .I3(n66631), .O(n67912));
    defparam i52226_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51595_4_lut (.I0(n31_adj_5348), .I1(n29_adj_5347), .I2(n27_adj_5357), 
            .I3(n67912), .O(n67281));
    defparam i51595_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52429_4_lut (.I0(n37_adj_5341), .I1(n35_adj_5346), .I2(n33_adj_5350), 
            .I3(n67281), .O(n68115));
    defparam i52429_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_10_i16_3_lut (.I0(n130[9]), .I1(n130[21]), .I2(n43_adj_5338), 
            .I3(GND_net), .O(n16_adj_5404));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52224_3_lut (.I0(n6_adj_5238), .I1(n130[10]), .I2(n21_adj_5361), 
            .I3(GND_net), .O(n67910));   // verilog/motorControl.v(46[12:34])
    defparam i52224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52225_3_lut (.I0(n67910), .I1(n130[11]), .I2(n23_adj_5343), 
            .I3(GND_net), .O(n67911));   // verilog/motorControl.v(46[12:34])
    defparam i52225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i8_3_lut (.I0(n130[4]), .I1(n130[8]), .I2(n17_adj_5359), 
            .I3(GND_net), .O(n8_adj_5405));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i24_3_lut (.I0(n16_adj_5404), .I1(n130[22]), .I2(n45_adj_5337), 
            .I3(GND_net), .O(n24_adj_5406));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49913_4_lut (.I0(n43_adj_5338), .I1(n25_adj_5344), .I2(n23_adj_5343), 
            .I3(n65702), .O(n65599));
    defparam i49913_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51603_4_lut (.I0(n24_adj_5406), .I1(n8_adj_5405), .I2(n45_adj_5337), 
            .I3(n65581), .O(n67289));   // verilog/motorControl.v(46[12:34])
    defparam i51603_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51921_3_lut (.I0(n67911), .I1(n130[12]), .I2(n25_adj_5344), 
            .I3(GND_net), .O(n67607));   // verilog/motorControl.v(46[12:34])
    defparam i51921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_10_i4_4_lut (.I0(n130[0]), .I1(n130[1]), .I2(IntegralLimit[1]), 
            .I3(IntegralLimit[0]), .O(n4_adj_5407));   // verilog/motorControl.v(46[12:34])
    defparam LessThan_10_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i52173_3_lut (.I0(n4_adj_5407), .I1(n130[13]), .I2(n27_adj_5357), 
            .I3(GND_net), .O(n67859));   // verilog/motorControl.v(46[12:34])
    defparam i52173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52174_3_lut (.I0(n67859), .I1(n130[14]), .I2(n29_adj_5347), 
            .I3(GND_net), .O(n67860));   // verilog/motorControl.v(46[12:34])
    defparam i52174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49978_4_lut (.I0(n33_adj_5350), .I1(n31_adj_5348), .I2(n29_adj_5347), 
            .I3(n65676), .O(n65664));
    defparam i49978_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52466_4_lut (.I0(n30_adj_5392), .I1(n10_adj_5391), .I2(n35_adj_5346), 
            .I3(n65657), .O(n68152));   // verilog/motorControl.v(46[12:34])
    defparam i52466_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51923_3_lut (.I0(n67860), .I1(n130[15]), .I2(n31_adj_5348), 
            .I3(GND_net), .O(n67609));   // verilog/motorControl.v(46[12:34])
    defparam i51923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52601_4_lut (.I0(n67609), .I1(n68152), .I2(n35_adj_5346), 
            .I3(n65664), .O(n68287));   // verilog/motorControl.v(46[12:34])
    defparam i52601_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52602_3_lut (.I0(n68287), .I1(n130[18]), .I2(n37_adj_5341), 
            .I3(GND_net), .O(n68288));   // verilog/motorControl.v(46[12:34])
    defparam i52602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52564_3_lut (.I0(n68288), .I1(n130[19]), .I2(n39_adj_5336), 
            .I3(GND_net), .O(n68250));   // verilog/motorControl.v(46[12:34])
    defparam i52564_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49928_4_lut (.I0(n43_adj_5338), .I1(n41_adj_5335), .I2(n39_adj_5336), 
            .I3(n68115), .O(n65614));
    defparam i49928_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51926_4_lut (.I0(n67607), .I1(n67289), .I2(n45_adj_5337), 
            .I3(n65599), .O(n67612));   // verilog/motorControl.v(46[12:34])
    defparam i51926_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52510_3_lut (.I0(n68250), .I1(n130[20]), .I2(n41_adj_5335), 
            .I3(GND_net), .O(n40_adj_5408));   // verilog/motorControl.v(46[12:34])
    defparam i52510_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52232_4_lut (.I0(n40_adj_5408), .I1(n67612), .I2(n45_adj_5337), 
            .I3(n65614), .O(n67918));   // verilog/motorControl.v(46[12:34])
    defparam i52232_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52233_3_lut (.I0(n67918), .I1(IntegralLimit[23]), .I2(n130[23]), 
            .I3(GND_net), .O(n155));   // verilog/motorControl.v(46[12:34])
    defparam i52233_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_12_i41_2_lut (.I0(n130[20]), .I1(n182[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35081_2_lut_3_lut (.I0(\Kp[1] ), .I1(n55[22]), .I2(n62_adj_5133), 
            .I3(GND_net), .O(n20100[0]));   // verilog/motorControl.v(51[18:24])
    defparam i35081_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i1_3_lut_4_lut (.I0(\Kp[1] ), .I1(n55[22]), .I2(n62_adj_5133), 
            .I3(n61894), .O(n20100[1]));   // verilog/motorControl.v(51[18:24])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 add_6161_21_lut (.I0(GND_net), .I1(n14934[18]), .I2(GND_net), 
            .I3(n49708), .O(n14095[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i39_2_lut (.I0(n130[19]), .I1(n182[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i45_2_lut (.I0(n130[22]), .I1(n182[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_5120));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i43_2_lut (.I0(n130[21]), .I1(n182[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5119));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6161_20_lut (.I0(GND_net), .I1(n14934[17]), .I2(GND_net), 
            .I3(n49707), .O(n14095[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6161_20 (.CI(n49707), .I0(n14934[17]), .I1(GND_net), 
            .CO(n49708));
    SB_LUT4 LessThan_12_i37_2_lut (.I0(n130[18]), .I1(n182[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5409));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6161_19_lut (.I0(GND_net), .I1(n14934[16]), .I2(GND_net), 
            .I3(n49706), .O(n14095[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6161_19 (.CI(n49706), .I0(n14934[16]), .I1(GND_net), 
            .CO(n49707));
    SB_LUT4 unary_minus_26_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n57[1]), 
            .I3(n49357), .O(n455)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6161_18_lut (.I0(GND_net), .I1(n14934[15]), .I2(GND_net), 
            .I3(n49705), .O(n14095[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_26_add_3_3 (.CI(n49357), .I0(GND_net), .I1(n57[1]), 
            .CO(n49358));
    SB_CARRY add_6161_18 (.CI(n49705), .I0(n14934[15]), .I1(GND_net), 
            .CO(n49706));
    SB_LUT4 unary_minus_26_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[1]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6161_17_lut (.I0(GND_net), .I1(n14934[14]), .I2(GND_net), 
            .I3(n49704), .O(n14095[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i29_2_lut (.I0(n130[14]), .I1(n182[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5411));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_26_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n57[0]), 
            .I3(VCC_net), .O(n456)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_26_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6161_17 (.CI(n49704), .I0(n14934[14]), .I1(GND_net), 
            .CO(n49705));
    SB_LUT4 add_6161_16_lut (.I0(GND_net), .I1(n14934[13]), .I2(n1105), 
            .I3(n49703), .O(n14095[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6161_16 (.CI(n49703), .I0(n14934[13]), .I1(n1105), .CO(n49704));
    SB_LUT4 add_6161_15_lut (.I0(GND_net), .I1(n14934[12]), .I2(n1032), 
            .I3(n49702), .O(n14095[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i31_2_lut (.I0(n130[15]), .I1(n182[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5412));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6161_15 (.CI(n49702), .I0(n14934[12]), .I1(n1032), .CO(n49703));
    SB_LUT4 add_6161_14_lut (.I0(GND_net), .I1(n14934[11]), .I2(n959), 
            .I3(n49701), .O(n14095[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6161_14 (.CI(n49701), .I0(n14934[11]), .I1(n959), .CO(n49702));
    SB_CARRY sub_8_add_2_20 (.CI(n49212), .I0(setpoint[18]), .I1(\motor_state[18] ), 
            .CO(n49213));
    SB_LUT4 add_6161_13_lut (.I0(GND_net), .I1(n14934[10]), .I2(n886), 
            .I3(n49700), .O(n14095[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i23_2_lut (.I0(n130[11]), .I1(n182[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5413));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_26_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n57[0]), 
            .CO(n49357));
    SB_CARRY add_6161_13 (.CI(n49700), .I0(n14934[10]), .I1(n886), .CO(n49701));
    SB_LUT4 add_6392_14_lut (.I0(GND_net), .I1(n18791[11]), .I2(n980_adj_5414), 
            .I3(n49486), .O(n18428[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6392_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6161_12_lut (.I0(GND_net), .I1(n14934[9]), .I2(n813_adj_5415), 
            .I3(n49699), .O(n14095[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6392_13_lut (.I0(GND_net), .I1(n18791[10]), .I2(n907_adj_5416), 
            .I3(n49485), .O(n18428[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6392_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_25_lut (.I0(n352[23]), .I1(GND_net), .I2(n61[23]), 
            .I3(n49356), .O(n47_adj_5417)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6161_12 (.CI(n49699), .I0(n14934[9]), .I1(n813_adj_5415), 
            .CO(n49700));
    SB_LUT4 add_6161_11_lut (.I0(GND_net), .I1(n14934[8]), .I2(n740_adj_5419), 
            .I3(n49698), .O(n14095[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6392_13 (.CI(n49485), .I0(n18791[10]), .I1(n907_adj_5416), 
            .CO(n49486));
    SB_CARRY add_6161_11 (.CI(n49698), .I0(n14934[8]), .I1(n740_adj_5419), 
            .CO(n49699));
    SB_LUT4 add_6161_10_lut (.I0(GND_net), .I1(n14934[7]), .I2(n667_adj_5420), 
            .I3(n49697), .O(n14095[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6161_10 (.CI(n49697), .I0(n14934[7]), .I1(n667_adj_5420), 
            .CO(n49698));
    SB_LUT4 add_6161_9_lut (.I0(GND_net), .I1(n14934[6]), .I2(n594_adj_5421), 
            .I3(n49696), .O(n14095[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6161_9 (.CI(n49696), .I0(n14934[6]), .I1(n594_adj_5421), 
            .CO(n49697));
    SB_LUT4 add_6161_8_lut (.I0(GND_net), .I1(n14934[5]), .I2(n521_adj_5422), 
            .I3(n49695), .O(n14095[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n61[22]), 
            .I3(n49355), .O(n63[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_24 (.CI(n49355), .I0(GND_net), .I1(n61[22]), 
            .CO(n49356));
    SB_CARRY add_6161_8 (.CI(n49695), .I0(n14934[5]), .I1(n521_adj_5422), 
            .CO(n49696));
    SB_LUT4 add_6392_12_lut (.I0(GND_net), .I1(n18791[9]), .I2(n834_adj_5424), 
            .I3(n49484), .O(n18428[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6392_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6161_7_lut (.I0(GND_net), .I1(n14934[4]), .I2(n448_adj_5425), 
            .I3(n49694), .O(n14095[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6392_12 (.CI(n49484), .I0(n18791[9]), .I1(n834_adj_5424), 
            .CO(n49485));
    SB_CARRY add_6161_7 (.CI(n49694), .I0(n14934[4]), .I1(n448_adj_5425), 
            .CO(n49695));
    SB_LUT4 add_6161_6_lut (.I0(GND_net), .I1(n14934[3]), .I2(n375_adj_5426), 
            .I3(n49693), .O(n14095[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(\motor_state[17] ), 
            .I3(n49211), .O(n55[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6392_11_lut (.I0(GND_net), .I1(n18791[8]), .I2(n761_adj_5427), 
            .I3(n49483), .O(n18428[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6392_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n61[21]), 
            .I3(n49354), .O(n63[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6161_6 (.CI(n49693), .I0(n14934[3]), .I1(n375_adj_5426), 
            .CO(n49694));
    SB_CARRY unary_minus_20_add_3_23 (.CI(n49354), .I0(GND_net), .I1(n61[21]), 
            .CO(n49355));
    SB_CARRY add_6392_11 (.CI(n49483), .I0(n18791[8]), .I1(n761_adj_5427), 
            .CO(n49484));
    SB_LUT4 add_6161_5_lut (.I0(GND_net), .I1(n14934[2]), .I2(n302_adj_5430), 
            .I3(n49692), .O(n14095[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6392_10_lut (.I0(GND_net), .I1(n18791[7]), .I2(n688_adj_5431), 
            .I3(n49482), .O(n18428[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6392_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6161_5 (.CI(n49692), .I0(n14934[2]), .I1(n302_adj_5430), 
            .CO(n49693));
    SB_LUT4 add_6161_4_lut (.I0(GND_net), .I1(n14934[1]), .I2(n229_adj_5432), 
            .I3(n49691), .O(n14095[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6161_4 (.CI(n49691), .I0(n14934[1]), .I1(n229_adj_5432), 
            .CO(n49692));
    SB_LUT4 add_6161_3_lut (.I0(GND_net), .I1(n14934[0]), .I2(n156_adj_5433), 
            .I3(n49690), .O(n14095[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6161_3 (.CI(n49690), .I0(n14934[0]), .I1(n156_adj_5433), 
            .CO(n49691));
    SB_CARRY sub_8_add_2_19 (.CI(n49211), .I0(setpoint[17]), .I1(\motor_state[17] ), 
            .CO(n49212));
    SB_CARRY add_6392_10 (.CI(n49482), .I0(n18791[7]), .I1(n688_adj_5431), 
            .CO(n49483));
    SB_LUT4 unary_minus_20_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n61[20]), 
            .I3(n49353), .O(n63[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_22 (.CI(n49353), .I0(GND_net), .I1(n61[20]), 
            .CO(n49354));
    SB_LUT4 add_6161_2_lut (.I0(GND_net), .I1(n14_adj_5435), .I2(n83_adj_5436), 
            .I3(GND_net), .O(n14095[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6161_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6392_9_lut (.I0(GND_net), .I1(n18791[6]), .I2(n615_adj_5437), 
            .I3(n49481), .O(n18428[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6392_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6392_9 (.CI(n49481), .I0(n18791[6]), .I1(n615_adj_5437), 
            .CO(n49482));
    SB_LUT4 unary_minus_20_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n61[19]), 
            .I3(n49352), .O(n63[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6161_2 (.CI(GND_net), .I0(n14_adj_5435), .I1(n83_adj_5436), 
            .CO(n49690));
    SB_LUT4 add_6392_8_lut (.I0(GND_net), .I1(n18791[5]), .I2(n542_adj_5439), 
            .I3(n49480), .O(n18428[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6392_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_21 (.CI(n49352), .I0(GND_net), .I1(n61[19]), 
            .CO(n49353));
    SB_CARRY add_6392_8 (.CI(n49480), .I0(n18791[5]), .I1(n542_adj_5439), 
            .CO(n49481));
    SB_LUT4 add_6392_7_lut (.I0(GND_net), .I1(n18791[4]), .I2(n469_adj_5440), 
            .I3(n49479), .O(n18428[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6392_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6392_7 (.CI(n49479), .I0(n18791[4]), .I1(n469_adj_5440), 
            .CO(n49480));
    SB_LUT4 add_6392_6_lut (.I0(GND_net), .I1(n18791[3]), .I2(n396_adj_5441), 
            .I3(n49478), .O(n18428[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6392_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n61[18]), 
            .I3(n49351), .O(n63[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6491_10_lut (.I0(GND_net), .I1(n19860[7]), .I2(n700_adj_5444), 
            .I3(n49689), .O(n19702[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6491_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(n20), 
            .I3(n49210), .O(n55[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6491_9_lut (.I0(GND_net), .I1(n19860[6]), .I2(n627_adj_5446), 
            .I3(n49688), .O(n19702[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6491_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_20 (.CI(n49351), .I0(GND_net), .I1(n61[18]), 
            .CO(n49352));
    SB_LUT4 unary_minus_20_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n61[17]), 
            .I3(n49350), .O(n63[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6491_9 (.CI(n49688), .I0(n19860[6]), .I1(n627_adj_5446), 
            .CO(n49689));
    SB_LUT4 LessThan_12_i25_2_lut (.I0(n130[12]), .I1(n182[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5448));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_8_add_2_18 (.CI(n49210), .I0(setpoint[16]), .I1(n20), 
            .CO(n49211));
    SB_CARRY add_6392_6 (.CI(n49478), .I0(n18791[3]), .I1(n396_adj_5441), 
            .CO(n49479));
    SB_LUT4 add_6491_8_lut (.I0(GND_net), .I1(n19860[5]), .I2(n554_adj_5449), 
            .I3(n49687), .O(n19702[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6491_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(\motor_state[15] ), 
            .I3(n49209), .O(n55[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6491_8 (.CI(n49687), .I0(n19860[5]), .I1(n554_adj_5449), 
            .CO(n49688));
    SB_CARRY unary_minus_20_add_3_19 (.CI(n49350), .I0(GND_net), .I1(n61[17]), 
            .CO(n49351));
    SB_CARRY sub_8_add_2_17 (.CI(n49209), .I0(setpoint[15]), .I1(\motor_state[15] ), 
            .CO(n49210));
    SB_LUT4 sub_8_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(\motor_state[14] ), 
            .I3(n49208), .O(n55[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6491_7_lut (.I0(GND_net), .I1(n19860[4]), .I2(n481_adj_5450), 
            .I3(n49686), .O(n19702[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6491_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_16 (.CI(n49208), .I0(setpoint[14]), .I1(\motor_state[14] ), 
            .CO(n49209));
    SB_CARRY add_6491_7 (.CI(n49686), .I0(n19860[4]), .I1(n481_adj_5450), 
            .CO(n49687));
    SB_LUT4 add_6491_6_lut (.I0(GND_net), .I1(n19860[3]), .I2(n408_adj_5451), 
            .I3(n49685), .O(n19702[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6491_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6491_6 (.CI(n49685), .I0(n19860[3]), .I1(n408_adj_5451), 
            .CO(n49686));
    SB_LUT4 unary_minus_20_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n61[16]), 
            .I3(n49349), .O(n63[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6491_5_lut (.I0(GND_net), .I1(n19860[2]), .I2(n335_adj_5453), 
            .I3(n49684), .O(n19702[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6491_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6491_5 (.CI(n49684), .I0(n19860[2]), .I1(n335_adj_5453), 
            .CO(n49685));
    SB_CARRY unary_minus_20_add_3_18 (.CI(n49349), .I0(GND_net), .I1(n61[16]), 
            .CO(n49350));
    SB_LUT4 add_6491_4_lut (.I0(GND_net), .I1(n19860[1]), .I2(n262_adj_5454), 
            .I3(n49683), .O(n19702[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6491_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6491_4 (.CI(n49683), .I0(n19860[1]), .I1(n262_adj_5454), 
            .CO(n49684));
    SB_LUT4 add_6392_5_lut (.I0(GND_net), .I1(n18791[2]), .I2(n323_adj_5455), 
            .I3(n49477), .O(n18428[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6392_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6392_5 (.CI(n49477), .I0(n18791[2]), .I1(n323_adj_5455), 
            .CO(n49478));
    SB_LUT4 add_6491_3_lut (.I0(GND_net), .I1(n19860[0]), .I2(n189_adj_5456), 
            .I3(n49682), .O(n19702[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6491_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(\motor_state[13] ), 
            .I3(n49207), .O(n55[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6392_4_lut (.I0(GND_net), .I1(n18791[1]), .I2(n250_adj_5457), 
            .I3(n49476), .O(n18428[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6392_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6491_3 (.CI(n49682), .I0(n19860[0]), .I1(n189_adj_5456), 
            .CO(n49683));
    SB_LUT4 add_6491_2_lut (.I0(GND_net), .I1(n47_adj_5458), .I2(n116_adj_5459), 
            .I3(GND_net), .O(n19702[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6491_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_15 (.CI(n49207), .I0(setpoint[13]), .I1(\motor_state[13] ), 
            .CO(n49208));
    SB_LUT4 unary_minus_20_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n61[15]), 
            .I3(n49348), .O(n63[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6491_2 (.CI(GND_net), .I0(n47_adj_5458), .I1(n116_adj_5459), 
            .CO(n49682));
    SB_CARRY add_6392_4 (.CI(n49476), .I0(n18791[1]), .I1(n250_adj_5457), 
            .CO(n49477));
    SB_CARRY unary_minus_20_add_3_17 (.CI(n49348), .I0(GND_net), .I1(n61[15]), 
            .CO(n49349));
    SB_LUT4 sub_8_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(\motor_state[12] ), 
            .I3(n49206), .O(n55[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6392_3_lut (.I0(GND_net), .I1(n18791[0]), .I2(n177_adj_5462), 
            .I3(n49475), .O(n18428[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6392_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6392_3 (.CI(n49475), .I0(n18791[0]), .I1(n177_adj_5462), 
            .CO(n49476));
    SB_CARRY sub_8_add_2_14 (.CI(n49206), .I0(setpoint[12]), .I1(\motor_state[12] ), 
            .CO(n49207));
    SB_LUT4 sub_8_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(n1), 
            .I3(n49205), .O(n55[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n61[14]), 
            .I3(n49347), .O(n63[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_16 (.CI(n49347), .I0(GND_net), .I1(n61[14]), 
            .CO(n49348));
    SB_CARRY sub_8_add_2_13 (.CI(n49205), .I0(setpoint[11]), .I1(n1), 
            .CO(n49206));
    SB_LUT4 unary_minus_20_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n61[13]), 
            .I3(n49346), .O(n63[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6392_2_lut (.I0(GND_net), .I1(n35_adj_5465), .I2(n104_adj_5466), 
            .I3(GND_net), .O(n18428[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6392_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(\motor_state[10] ), 
            .I3(n49204), .O(n55[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6392_2 (.CI(GND_net), .I0(n35_adj_5465), .I1(n104_adj_5466), 
            .CO(n49475));
    SB_CARRY unary_minus_20_add_3_15 (.CI(n49346), .I0(GND_net), .I1(n61[13]), 
            .CO(n49347));
    SB_LUT4 unary_minus_20_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n61[12]), 
            .I3(n49345), .O(n63[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_14 (.CI(n49345), .I0(GND_net), .I1(n61[12]), 
            .CO(n49346));
    SB_LUT4 unary_minus_20_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n61[11]), 
            .I3(n49344), .O(n63[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_13 (.CI(n49344), .I0(GND_net), .I1(n61[11]), 
            .CO(n49345));
    SB_LUT4 unary_minus_20_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n61[10]), 
            .I3(n49343), .O(n63[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_12 (.CI(n49343), .I0(GND_net), .I1(n61[10]), 
            .CO(n49344));
    SB_LUT4 unary_minus_20_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n61[9]), 
            .I3(n49342), .O(n63[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_12 (.CI(n49204), .I0(setpoint[10]), .I1(\motor_state[10] ), 
            .CO(n49205));
    SB_CARRY unary_minus_20_add_3_11 (.CI(n49342), .I0(GND_net), .I1(n61[9]), 
            .CO(n49343));
    SB_LUT4 unary_minus_20_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n61[8]), 
            .I3(n49341), .O(n63[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_10 (.CI(n49341), .I0(GND_net), .I1(n61[8]), 
            .CO(n49342));
    SB_LUT4 sub_8_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(\motor_state[9] ), 
            .I3(n49203), .O(n55[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_25_lut (.I0(GND_net), .I1(n11650[0]), .I2(n12226[0]), 
            .I3(n49263), .O(n352[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6200_20_lut (.I0(GND_net), .I1(n15693[17]), .I2(GND_net), 
            .I3(n49666), .O(n14934[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n61[7]), 
            .I3(n49340), .O(n63[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6200_19_lut (.I0(GND_net), .I1(n15693[16]), .I2(GND_net), 
            .I3(n49665), .O(n14934[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6200_19 (.CI(n49665), .I0(n15693[16]), .I1(GND_net), 
            .CO(n49666));
    SB_CARRY unary_minus_20_add_3_9 (.CI(n49340), .I0(GND_net), .I1(n61[7]), 
            .CO(n49341));
    SB_LUT4 add_6200_18_lut (.I0(GND_net), .I1(n15693[15]), .I2(GND_net), 
            .I3(n49664), .O(n14934[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n61[6]), 
            .I3(n49339), .O(n63[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_11 (.CI(n49203), .I0(setpoint[9]), .I1(\motor_state[9] ), 
            .CO(n49204));
    SB_CARRY add_6200_18 (.CI(n49664), .I0(n15693[15]), .I1(GND_net), 
            .CO(n49665));
    SB_LUT4 add_6200_17_lut (.I0(GND_net), .I1(n15693[14]), .I2(GND_net), 
            .I3(n49663), .O(n14934[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6200_17 (.CI(n49663), .I0(n15693[14]), .I1(GND_net), 
            .CO(n49664));
    SB_LUT4 add_18_24_lut (.I0(GND_net), .I1(n257[22]), .I2(n49[22]), 
            .I3(n49262), .O(n352[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6200_16_lut (.I0(GND_net), .I1(n15693[13]), .I2(n1108_adj_5477), 
            .I3(n49662), .O(n14934[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_8 (.CI(n49339), .I0(GND_net), .I1(n61[6]), 
            .CO(n49340));
    SB_CARRY add_6200_16 (.CI(n49662), .I0(n15693[13]), .I1(n1108_adj_5477), 
            .CO(n49663));
    SB_LUT4 add_6200_15_lut (.I0(GND_net), .I1(n15693[12]), .I2(n1035_adj_5478), 
            .I3(n49661), .O(n14934[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_24 (.CI(n49262), .I0(n257[22]), .I1(n49[22]), .CO(n49263));
    SB_CARRY add_6200_15 (.CI(n49661), .I0(n15693[12]), .I1(n1035_adj_5478), 
            .CO(n49662));
    SB_LUT4 unary_minus_20_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n61[5]), 
            .I3(n49338), .O(n63[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6200_14_lut (.I0(GND_net), .I1(n15693[11]), .I2(n962_adj_5480), 
            .I3(n49660), .O(n14934[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6200_14 (.CI(n49660), .I0(n15693[11]), .I1(n962_adj_5480), 
            .CO(n49661));
    SB_LUT4 add_6200_13_lut (.I0(GND_net), .I1(n15693[10]), .I2(n889_adj_5481), 
            .I3(n49659), .O(n14934[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_7 (.CI(n49338), .I0(GND_net), .I1(n61[5]), 
            .CO(n49339));
    SB_LUT4 add_18_23_lut (.I0(GND_net), .I1(n257[21]), .I2(n49[21]), 
            .I3(n49261), .O(n352[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6200_13 (.CI(n49659), .I0(n15693[10]), .I1(n889_adj_5481), 
            .CO(n49660));
    SB_LUT4 add_6200_12_lut (.I0(GND_net), .I1(n15693[9]), .I2(n816_adj_5482), 
            .I3(n49658), .O(n14934[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n61[4]), 
            .I3(n49337), .O(n63[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_6 (.CI(n49337), .I0(GND_net), .I1(n61[4]), 
            .CO(n49338));
    SB_LUT4 unary_minus_20_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n61[3]), 
            .I3(n49336), .O(n63[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6200_12 (.CI(n49658), .I0(n15693[9]), .I1(n816_adj_5482), 
            .CO(n49659));
    SB_LUT4 add_6200_11_lut (.I0(GND_net), .I1(n15693[8]), .I2(n743_adj_5486), 
            .I3(n49657), .O(n14934[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6200_11 (.CI(n49657), .I0(n15693[8]), .I1(n743_adj_5486), 
            .CO(n49658));
    SB_LUT4 sub_8_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(\motor_state[8] ), 
            .I3(n49202), .O(n55[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_5 (.CI(n49336), .I0(GND_net), .I1(n61[3]), 
            .CO(n49337));
    SB_CARRY add_18_23 (.CI(n49261), .I0(n257[21]), .I1(n49[21]), .CO(n49262));
    SB_LUT4 add_6200_10_lut (.I0(GND_net), .I1(n15693[7]), .I2(n670_adj_5487), 
            .I3(n49656), .O(n14934[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_22_lut (.I0(GND_net), .I1(n257[20]), .I2(n49[20]), 
            .I3(n49260), .O(n352[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n61[2]), 
            .I3(n49335), .O(n63[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_4 (.CI(n49335), .I0(GND_net), .I1(n61[2]), 
            .CO(n49336));
    SB_CARRY add_6200_10 (.CI(n49656), .I0(n15693[7]), .I1(n670_adj_5487), 
            .CO(n49657));
    SB_LUT4 add_6200_9_lut (.I0(GND_net), .I1(n15693[6]), .I2(n597_adj_5489), 
            .I3(n49655), .O(n14934[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n61[1]), 
            .I3(n49334), .O(n401)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6200_9 (.CI(n49655), .I0(n15693[6]), .I1(n597_adj_5489), 
            .CO(n49656));
    SB_CARRY add_18_22 (.CI(n49260), .I0(n257[20]), .I1(n49[20]), .CO(n49261));
    SB_LUT4 add_6200_8_lut (.I0(GND_net), .I1(n15693[5]), .I2(n524_adj_5491), 
            .I3(n49654), .O(n14934[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6200_8 (.CI(n49654), .I0(n15693[5]), .I1(n524_adj_5491), 
            .CO(n49655));
    SB_LUT4 add_6200_7_lut (.I0(GND_net), .I1(n15693[4]), .I2(n451_adj_5492), 
            .I3(n49653), .O(n14934[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6200_7 (.CI(n49653), .I0(n15693[4]), .I1(n451_adj_5492), 
            .CO(n49654));
    SB_LUT4 add_6200_6_lut (.I0(GND_net), .I1(n15693[3]), .I2(n378_adj_5493), 
            .I3(n49652), .O(n14934[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_21_lut (.I0(GND_net), .I1(n257[19]), .I2(n49[19]), 
            .I3(n49259), .O(n352[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6200_6 (.CI(n49652), .I0(n15693[3]), .I1(n378_adj_5493), 
            .CO(n49653));
    SB_LUT4 add_6200_5_lut (.I0(GND_net), .I1(n15693[2]), .I2(n305_adj_5494), 
            .I3(n49651), .O(n14934[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6200_5 (.CI(n49651), .I0(n15693[2]), .I1(n305_adj_5494), 
            .CO(n49652));
    SB_LUT4 add_6200_4_lut (.I0(GND_net), .I1(n15693[1]), .I2(n232_adj_5495), 
            .I3(n49650), .O(n14934[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6200_4 (.CI(n49650), .I0(n15693[1]), .I1(n232_adj_5495), 
            .CO(n49651));
    SB_CARRY unary_minus_20_add_3_3 (.CI(n49334), .I0(GND_net), .I1(n61[1]), 
            .CO(n49335));
    SB_LUT4 add_6200_3_lut (.I0(GND_net), .I1(n15693[0]), .I2(n159_adj_5496), 
            .I3(n49649), .O(n14934[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_2_lut (.I0(n37174), .I1(GND_net), .I2(n61[0]), 
            .I3(VCC_net), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_6200_3 (.CI(n49649), .I0(n15693[0]), .I1(n159_adj_5496), 
            .CO(n49650));
    SB_LUT4 add_6200_2_lut (.I0(GND_net), .I1(n17_adj_5499), .I2(n86_adj_5500), 
            .I3(GND_net), .O(n14934[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6200_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_21 (.CI(n49259), .I0(n257[19]), .I1(n49[19]), .CO(n49260));
    SB_CARRY add_6200_2 (.CI(GND_net), .I0(n17_adj_5499), .I1(n86_adj_5500), 
            .CO(n49649));
    SB_CARRY unary_minus_20_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n61[0]), 
            .CO(n49334));
    SB_LUT4 add_18_20_lut (.I0(GND_net), .I1(n257[18]), .I2(n49[18]), 
            .I3(n49258), .O(n352[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n65[23]), 
            .I3(n49333), .O(n182[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_20 (.CI(n49258), .I0(n257[18]), .I1(n49[18]), .CO(n49259));
    SB_LUT4 unary_minus_13_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n65[22]), 
            .I3(n49332), .O(n182[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_10 (.CI(n49202), .I0(setpoint[8]), .I1(\motor_state[8] ), 
            .CO(n49203));
    SB_LUT4 add_18_19_lut (.I0(GND_net), .I1(n257[17]), .I2(n49[17]), 
            .I3(n49257), .O(n352[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_19 (.CI(n49257), .I0(n257[17]), .I1(n49[17]), .CO(n49258));
    SB_LUT4 add_18_18_lut (.I0(GND_net), .I1(n257[16]), .I2(n49[16]), 
            .I3(n49256), .O(n352[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_8_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(\motor_state[7] ), 
            .I3(n49201), .O(n55[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_9 (.CI(n49201), .I0(setpoint[7]), .I1(\motor_state[7] ), 
            .CO(n49202));
    SB_LUT4 sub_8_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(n41622), 
            .I3(n49200), .O(n55[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_8 (.CI(n49200), .I0(setpoint[6]), .I1(n41622), 
            .CO(n49201));
    SB_LUT4 sub_8_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(\motor_state[5] ), 
            .I3(n49199), .O(n55[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_18 (.CI(n49256), .I0(n257[16]), .I1(n49[16]), .CO(n49257));
    SB_CARRY unary_minus_13_add_3_24 (.CI(n49332), .I0(GND_net), .I1(n65[22]), 
            .CO(n49333));
    SB_LUT4 unary_minus_13_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n65[21]), 
            .I3(n49331), .O(n182[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_23 (.CI(n49331), .I0(GND_net), .I1(n65[21]), 
            .CO(n49332));
    SB_LUT4 unary_minus_13_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n65[20]), 
            .I3(n49330), .O(n182[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_22 (.CI(n49330), .I0(GND_net), .I1(n65[20]), 
            .CO(n49331));
    SB_LUT4 unary_minus_13_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n65[19]), 
            .I3(n49329), .O(n182[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_17_lut (.I0(GND_net), .I1(n257[15]), .I2(n49[15]), 
            .I3(n49255), .O(n361)) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6237_19_lut (.I0(GND_net), .I1(n16376[16]), .I2(GND_net), 
            .I3(n49634), .O(n15693[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6237_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_7 (.CI(n49199), .I0(setpoint[5]), .I1(\motor_state[5] ), 
            .CO(n49200));
    SB_CARRY add_18_17 (.CI(n49255), .I0(n257[15]), .I1(n49[15]), .CO(n49256));
    SB_LUT4 add_6237_18_lut (.I0(GND_net), .I1(n16376[15]), .I2(GND_net), 
            .I3(n49633), .O(n15693[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6237_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_16_lut (.I0(GND_net), .I1(n257[14]), .I2(n49[14]), 
            .I3(n49254), .O(n352[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6237_18 (.CI(n49633), .I0(n16376[15]), .I1(GND_net), 
            .CO(n49634));
    SB_LUT4 sub_8_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(\motor_state[4] ), 
            .I3(n49198), .O(n55[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_8_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6237_17_lut (.I0(GND_net), .I1(n16376[14]), .I2(GND_net), 
            .I3(n49632), .O(n15693[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6237_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_21 (.CI(n49329), .I0(GND_net), .I1(n65[19]), 
            .CO(n49330));
    SB_LUT4 unary_minus_13_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n65[18]), 
            .I3(n49328), .O(n182[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_20 (.CI(n49328), .I0(GND_net), .I1(n65[18]), 
            .CO(n49329));
    SB_CARRY add_6237_17 (.CI(n49632), .I0(n16376[14]), .I1(GND_net), 
            .CO(n49633));
    SB_LUT4 unary_minus_13_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n65[17]), 
            .I3(n49327), .O(n182[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6237_16_lut (.I0(GND_net), .I1(n16376[13]), .I2(n1111_adj_5509), 
            .I3(n49631), .O(n15693[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6237_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6237_16 (.CI(n49631), .I0(n16376[13]), .I1(n1111_adj_5509), 
            .CO(n49632));
    SB_CARRY sub_8_add_2_6 (.CI(n49198), .I0(setpoint[4]), .I1(\motor_state[4] ), 
            .CO(n49199));
    SB_LUT4 add_6237_15_lut (.I0(GND_net), .I1(n16376[12]), .I2(n1038_adj_5510), 
            .I3(n49630), .O(n15693[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6237_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6237_15 (.CI(n49630), .I0(n16376[12]), .I1(n1038_adj_5510), 
            .CO(n49631));
    SB_CARRY add_18_16 (.CI(n49254), .I0(n257[14]), .I1(n49[14]), .CO(n49255));
    SB_CARRY unary_minus_13_add_3_19 (.CI(n49327), .I0(GND_net), .I1(n65[17]), 
            .CO(n49328));
    SB_LUT4 add_6237_14_lut (.I0(GND_net), .I1(n16376[11]), .I2(n965_adj_5511), 
            .I3(n49629), .O(n15693[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6237_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_5 (.CI(n49197), .I0(setpoint[3]), .I1(n42235), 
            .CO(n49198));
    SB_CARRY add_6237_14 (.CI(n49629), .I0(n16376[11]), .I1(n965_adj_5511), 
            .CO(n49630));
    SB_LUT4 add_18_15_lut (.I0(GND_net), .I1(n257[13]), .I2(n49[13]), 
            .I3(n49253), .O(n352[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_4 (.CI(n49196), .I0(setpoint[2]), .I1(\motor_state[2] ), 
            .CO(n49197));
    SB_LUT4 unary_minus_13_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n65[16]), 
            .I3(n49326), .O(n182[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6237_13_lut (.I0(GND_net), .I1(n16376[10]), .I2(n892_adj_5513), 
            .I3(n49628), .O(n15693[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6237_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_18 (.CI(n49326), .I0(GND_net), .I1(n65[16]), 
            .CO(n49327));
    SB_LUT4 add_6417_13_lut (.I0(GND_net), .I1(n19102[10]), .I2(n910_adj_5514), 
            .I3(n49448), .O(n18791[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6417_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6417_12_lut (.I0(GND_net), .I1(n19102[9]), .I2(n837_adj_5515), 
            .I3(n49447), .O(n18791[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6417_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6237_13 (.CI(n49628), .I0(n16376[10]), .I1(n892_adj_5513), 
            .CO(n49629));
    SB_CARRY sub_8_add_2_3 (.CI(n49195), .I0(setpoint[1]), .I1(\motor_state[1] ), 
            .CO(n49196));
    SB_CARRY add_18_15 (.CI(n49253), .I0(n257[13]), .I1(n49[13]), .CO(n49254));
    SB_CARRY add_6417_12 (.CI(n49447), .I0(n19102[9]), .I1(n837_adj_5515), 
            .CO(n49448));
    SB_LUT4 unary_minus_13_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n65[15]), 
            .I3(n49325), .O(n182[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_17 (.CI(n49325), .I0(GND_net), .I1(n65[15]), 
            .CO(n49326));
    SB_LUT4 add_18_14_lut (.I0(GND_net), .I1(n257[12]), .I2(n49[12]), 
            .I3(n49252), .O(n352[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_8_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(\motor_state[0] ), 
            .CO(n49195));
    SB_LUT4 add_6417_11_lut (.I0(GND_net), .I1(n19102[8]), .I2(n764_adj_5517), 
            .I3(n49446), .O(n18791[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6417_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6237_12_lut (.I0(GND_net), .I1(n16376[9]), .I2(n819_adj_5518), 
            .I3(n49627), .O(n15693[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6237_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6237_12 (.CI(n49627), .I0(n16376[9]), .I1(n819_adj_5518), 
            .CO(n49628));
    SB_CARRY add_6417_11 (.CI(n49446), .I0(n19102[8]), .I1(n764_adj_5517), 
            .CO(n49447));
    SB_CARRY add_18_14 (.CI(n49252), .I0(n257[12]), .I1(n49[12]), .CO(n49253));
    SB_LUT4 add_18_13_lut (.I0(GND_net), .I1(n257[11]), .I2(n49[11]), 
            .I3(n49251), .O(n352[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n65[14]), 
            .I3(n49324), .O(n182[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_13 (.CI(n49251), .I0(n257[11]), .I1(n49[11]), .CO(n49252));
    SB_LUT4 add_6417_10_lut (.I0(GND_net), .I1(n19102[7]), .I2(n691_adj_5520), 
            .I3(n49445), .O(n18791[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6417_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6417_10 (.CI(n49445), .I0(n19102[7]), .I1(n691_adj_5520), 
            .CO(n49446));
    SB_LUT4 add_6417_9_lut (.I0(GND_net), .I1(n19102[6]), .I2(n618_adj_5521), 
            .I3(n49444), .O(n18791[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6417_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6237_11_lut (.I0(GND_net), .I1(n16376[8]), .I2(n746_adj_5522), 
            .I3(n49626), .O(n15693[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6237_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6237_11 (.CI(n49626), .I0(n16376[8]), .I1(n746_adj_5522), 
            .CO(n49627));
    SB_LUT4 add_18_12_lut (.I0(GND_net), .I1(n257[10]), .I2(n49[10]), 
            .I3(n49250), .O(n352[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6237_10_lut (.I0(GND_net), .I1(n16376[7]), .I2(n673_adj_5523), 
            .I3(n49625), .O(n15693[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6237_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6417_9 (.CI(n49444), .I0(n19102[6]), .I1(n618_adj_5521), 
            .CO(n49445));
    SB_CARRY add_6237_10 (.CI(n49625), .I0(n16376[7]), .I1(n673_adj_5523), 
            .CO(n49626));
    SB_LUT4 mult_17_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i257_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_18_12 (.CI(n49250), .I0(n257[10]), .I1(n49[10]), .CO(n49251));
    SB_CARRY unary_minus_13_add_3_16 (.CI(n49324), .I0(GND_net), .I1(n65[14]), 
            .CO(n49325));
    SB_LUT4 add_6237_9_lut (.I0(GND_net), .I1(n16376[6]), .I2(n600_adj_5524), 
            .I3(n49624), .O(n15693[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6237_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6237_9 (.CI(n49624), .I0(n16376[6]), .I1(n600_adj_5524), 
            .CO(n49625));
    SB_LUT4 add_6417_8_lut (.I0(GND_net), .I1(n19102[5]), .I2(n545_adj_5525), 
            .I3(n49443), .O(n18791[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6417_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6417_8 (.CI(n49443), .I0(n19102[5]), .I1(n545_adj_5525), 
            .CO(n49444));
    SB_LUT4 add_18_11_lut (.I0(GND_net), .I1(n257[9]), .I2(n49[9]), .I3(n49249), 
            .O(n352[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n65[13]), 
            .I3(n49323), .O(n182[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6417_7_lut (.I0(GND_net), .I1(n19102[4]), .I2(n472_adj_5527), 
            .I3(n49442), .O(n18791[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6417_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_11 (.CI(n49249), .I0(n257[9]), .I1(n49[9]), .CO(n49250));
    SB_CARRY add_6417_7 (.CI(n49442), .I0(n19102[4]), .I1(n472_adj_5527), 
            .CO(n49443));
    SB_CARRY unary_minus_13_add_3_15 (.CI(n49323), .I0(GND_net), .I1(n65[13]), 
            .CO(n49324));
    SB_LUT4 add_6417_6_lut (.I0(GND_net), .I1(n19102[3]), .I2(n399_adj_5528), 
            .I3(n49441), .O(n18791[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6417_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6417_6 (.CI(n49441), .I0(n19102[3]), .I1(n399_adj_5528), 
            .CO(n49442));
    SB_LUT4 unary_minus_13_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n65[12]), 
            .I3(n49322), .O(n182[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_14 (.CI(n49322), .I0(GND_net), .I1(n65[12]), 
            .CO(n49323));
    SB_LUT4 add_18_10_lut (.I0(GND_net), .I1(n257[8]), .I2(n49[8]), .I3(n49248), 
            .O(n352[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6417_5_lut (.I0(GND_net), .I1(n19102[2]), .I2(n326_adj_5530), 
            .I3(n49440), .O(n18791[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6417_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6237_8_lut (.I0(GND_net), .I1(n16376[5]), .I2(n527_adj_5531), 
            .I3(n49623), .O(n15693[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6237_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6237_8 (.CI(n49623), .I0(n16376[5]), .I1(n527_adj_5531), 
            .CO(n49624));
    SB_CARRY add_18_10 (.CI(n49248), .I0(n257[8]), .I1(n49[8]), .CO(n49249));
    SB_LUT4 unary_minus_13_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n65[11]), 
            .I3(n49321), .O(n182[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6237_7_lut (.I0(GND_net), .I1(n16376[4]), .I2(n454_adj_5533), 
            .I3(n49622), .O(n15693[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6237_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6417_5 (.CI(n49440), .I0(n19102[2]), .I1(n326_adj_5530), 
            .CO(n49441));
    SB_CARRY add_6237_7 (.CI(n49622), .I0(n16376[4]), .I1(n454_adj_5533), 
            .CO(n49623));
    SB_CARRY unary_minus_13_add_3_13 (.CI(n49321), .I0(GND_net), .I1(n65[11]), 
            .CO(n49322));
    SB_LUT4 add_6237_6_lut (.I0(GND_net), .I1(n16376[3]), .I2(n381_adj_5534), 
            .I3(n49621), .O(n15693[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6237_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_9_lut (.I0(GND_net), .I1(n257[7]), .I2(n49[7]), .I3(n49247), 
            .O(n352[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6417_4_lut (.I0(GND_net), .I1(n19102[1]), .I2(n253_adj_5535), 
            .I3(n49439), .O(n18791[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6417_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6237_6 (.CI(n49621), .I0(n16376[3]), .I1(n381_adj_5534), 
            .CO(n49622));
    SB_CARRY add_6417_4 (.CI(n49439), .I0(n19102[1]), .I1(n253_adj_5535), 
            .CO(n49440));
    SB_LUT4 add_6237_5_lut (.I0(GND_net), .I1(n16376[2]), .I2(n308_adj_5536), 
            .I3(n49620), .O(n15693[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6237_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6237_5 (.CI(n49620), .I0(n16376[2]), .I1(n308_adj_5536), 
            .CO(n49621));
    SB_CARRY add_18_9 (.CI(n49247), .I0(n257[7]), .I1(n49[7]), .CO(n49248));
    SB_LUT4 unary_minus_13_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n65[10]), 
            .I3(n49320), .O(n182[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6417_3_lut (.I0(GND_net), .I1(n19102[0]), .I2(n180_adj_5538), 
            .I3(n49438), .O(n18791[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6417_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_8_lut (.I0(GND_net), .I1(n257[6]), .I2(n49[6]), .I3(n49246), 
            .O(n352[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6237_4_lut (.I0(GND_net), .I1(n16376[1]), .I2(n235_adj_5539), 
            .I3(n49619), .O(n15693[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6237_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6417_3 (.CI(n49438), .I0(n19102[0]), .I1(n180_adj_5538), 
            .CO(n49439));
    SB_CARRY add_18_8 (.CI(n49246), .I0(n257[6]), .I1(n49[6]), .CO(n49247));
    SB_CARRY add_6237_4 (.CI(n49619), .I0(n16376[1]), .I1(n235_adj_5539), 
            .CO(n49620));
    SB_CARRY unary_minus_13_add_3_12 (.CI(n49320), .I0(GND_net), .I1(n65[10]), 
            .CO(n49321));
    SB_LUT4 add_6237_3_lut (.I0(GND_net), .I1(n16376[0]), .I2(n162_adj_5540), 
            .I3(n49618), .O(n15693[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6237_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6417_2_lut (.I0(GND_net), .I1(n38_adj_5541), .I2(n107_adj_5542), 
            .I3(GND_net), .O(n18791[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6417_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6237_3 (.CI(n49618), .I0(n16376[0]), .I1(n162_adj_5540), 
            .CO(n49619));
    SB_CARRY add_6417_2 (.CI(GND_net), .I0(n38_adj_5541), .I1(n107_adj_5542), 
            .CO(n49438));
    SB_LUT4 add_6237_2_lut (.I0(GND_net), .I1(n20_adj_5543), .I2(n89_adj_5544), 
            .I3(GND_net), .O(n15693[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6237_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6237_2 (.CI(GND_net), .I0(n20_adj_5543), .I1(n89_adj_5544), 
            .CO(n49618));
    SB_LUT4 add_18_7_lut (.I0(GND_net), .I1(n257[5]), .I2(n49[5]), .I3(n49245), 
            .O(n352[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6507_9_lut (.I0(GND_net), .I1(n19984[6]), .I2(n630_adj_5545), 
            .I3(n49617), .O(n19860[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6507_8_lut (.I0(GND_net), .I1(n19984[5]), .I2(n557_adj_5546), 
            .I3(n49616), .O(n19860[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n65[9]), 
            .I3(n49319), .O(n182[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_11 (.CI(n49319), .I0(GND_net), .I1(n65[9]), 
            .CO(n49320));
    SB_CARRY add_6507_8 (.CI(n49616), .I0(n19984[5]), .I1(n557_adj_5546), 
            .CO(n49617));
    SB_LUT4 mult_17_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i306_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_18_7 (.CI(n49245), .I0(n257[5]), .I1(n49[5]), .CO(n49246));
    SB_LUT4 unary_minus_13_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n65[8]), 
            .I3(n49318), .O(n182[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_10 (.CI(n49318), .I0(GND_net), .I1(n65[8]), 
            .CO(n49319));
    SB_LUT4 unary_minus_13_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n65[7]), 
            .I3(n49317), .O(n182[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6507_7_lut (.I0(GND_net), .I1(n19984[4]), .I2(n484_adj_5550), 
            .I3(n49615), .O(n19860[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6507_7 (.CI(n49615), .I0(n19984[4]), .I1(n484_adj_5550), 
            .CO(n49616));
    SB_LUT4 add_6507_6_lut (.I0(GND_net), .I1(n19984[3]), .I2(n411_adj_5551), 
            .I3(n49614), .O(n19860[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_6_lut (.I0(GND_net), .I1(n257[4]), .I2(n49[4]), .I3(n49244), 
            .O(n352[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_17_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n600));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n673));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i35_2_lut (.I0(n130[17]), .I1(n182[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5552));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i33_2_lut (.I0(n130[16]), .I1(n182[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5553));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i11_2_lut (.I0(n130[5]), .I1(n182[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5554));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n819));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i551_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_13_add_3_9 (.CI(n49317), .I0(GND_net), .I1(n65[7]), 
            .CO(n49318));
    SB_CARRY add_6507_6 (.CI(n49614), .I0(n19984[3]), .I1(n411_adj_5551), 
            .CO(n49615));
    SB_LUT4 unary_minus_13_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n65[6]), 
            .I3(n49316), .O(n182[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_8 (.CI(n49316), .I0(GND_net), .I1(n65[6]), 
            .CO(n49317));
    SB_LUT4 add_6507_5_lut (.I0(GND_net), .I1(n19984[2]), .I2(n338_adj_5556), 
            .I3(n49613), .O(n19860[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n65[5]), 
            .I3(n49315), .O(n182[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_18_6 (.CI(n49244), .I0(n257[4]), .I1(n49[4]), .CO(n49245));
    SB_CARRY add_6507_5 (.CI(n49613), .I0(n19984[2]), .I1(n338_adj_5556), 
            .CO(n49614));
    SB_LUT4 add_6507_4_lut (.I0(GND_net), .I1(n19984[1]), .I2(n265_adj_5558), 
            .I3(n49612), .O(n19860[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_18_5_lut (.I0(GND_net), .I1(n257[3]), .I2(n49[3]), .I3(n49243), 
            .O(n352[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6507_4 (.CI(n49612), .I0(n19984[1]), .I1(n265_adj_5558), 
            .CO(n49613));
    SB_CARRY unary_minus_13_add_3_7 (.CI(n49315), .I0(GND_net), .I1(n65[5]), 
            .CO(n49316));
    SB_LUT4 add_6507_3_lut (.I0(GND_net), .I1(n19984[0]), .I2(n192_adj_5559), 
            .I3(n49611), .O(n19860[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6507_3 (.CI(n49611), .I0(n19984[0]), .I1(n192_adj_5559), 
            .CO(n49612));
    SB_LUT4 LessThan_12_i13_2_lut (.I0(n130[6]), .I1(n182[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5560));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n892));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i15_2_lut (.I0(n130[7]), .I1(n182[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5561));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_17_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n965));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n1038));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n1111));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i557_2_lut (.I0(\Kp[11] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i27_2_lut (.I0(n130[13]), .I1(n182[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5562));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_12_i9_2_lut (.I0(n130[4]), .I1(n182[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5563));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6507_2_lut (.I0(GND_net), .I1(n50_adj_5564), .I2(n119_adj_5565), 
            .I3(GND_net), .O(n19860[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6507_2 (.CI(GND_net), .I0(n50_adj_5564), .I1(n119_adj_5565), 
            .CO(n49611));
    SB_LUT4 LessThan_12_i17_2_lut (.I0(n130[8]), .I1(n182[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5566));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_13_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n65[4]), 
            .I3(n49314), .O(n182[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_6 (.CI(n49314), .I0(GND_net), .I1(n65[4]), 
            .CO(n49315));
    SB_CARRY add_18_5 (.CI(n49243), .I0(n257[3]), .I1(n49[3]), .CO(n49244));
    SB_LUT4 unary_minus_13_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n65[3]), 
            .I3(n49313), .O(n182[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i77_2_lut (.I0(\Kp[1] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_5243));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i30_2_lut (.I0(\Kp[0] ), .I1(n55[18]), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i126_2_lut (.I0(\Kp[2] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_5242));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i175_2_lut (.I0(\Kp[3] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n259));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i224_2_lut (.I0(\Kp[4] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_5241));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i273_2_lut (.I0(\Kp[5] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n405_adj_5240));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_18_4_lut (.I0(GND_net), .I1(n257[2]), .I2(n49[2]), .I3(n49242), 
            .O(n352[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_16_i322_2_lut (.I0(\Kp[6] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_5237));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i371_2_lut (.I0(\Kp[7] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_5236));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i420_2_lut (.I0(\Kp[8] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_5235));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i606_2_lut (.I0(\Kp[12] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i469_2_lut (.I0(\Kp[9] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_5234));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i19_2_lut (.I0(n130[9]), .I1(n182[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5569));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i19_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_18_4 (.CI(n49242), .I0(n257[2]), .I1(n49[2]), .CO(n49243));
    SB_CARRY unary_minus_13_add_3_5 (.CI(n49313), .I0(GND_net), .I1(n65[3]), 
            .CO(n49314));
    SB_LUT4 unary_minus_13_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n65[2]), 
            .I3(n49312), .O(n182[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_4 (.CI(n49312), .I0(GND_net), .I1(n65[2]), 
            .CO(n49313));
    SB_LUT4 add_18_3_lut (.I0(GND_net), .I1(n257[1]), .I2(n49[1]), .I3(n49241), 
            .O(n375)) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_13_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n65[1]), 
            .I3(n49311), .O(n182[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_13_add_3_3 (.CI(n49311), .I0(GND_net), .I1(n65[1]), 
            .CO(n49312));
    SB_LUT4 unary_minus_13_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n65[0]), 
            .I3(VCC_net), .O(n182[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_13_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_12_i21_2_lut (.I0(n130[10]), .I1(n182[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5574));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i11_2_lut (.I0(PWMLimit[5]), .I1(n352[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5575));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i13_2_lut (.I0(PWMLimit[6]), .I1(n352[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5576));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_13_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n65[0]), 
            .CO(n49311));
    SB_LUT4 LessThan_23_i9_2_lut (.I0(PWMLimit[4]), .I1(n352[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5577));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i17_2_lut (.I0(PWMLimit[8]), .I1(n352[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5578));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_18_3 (.CI(n49241), .I0(n257[1]), .I1(n49[1]), .CO(n49242));
    SB_LUT4 LessThan_23_i7_2_lut (.I0(PWMLimit[3]), .I1(n352[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5579));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_18_2_lut (.I0(GND_net), .I1(n257[0]), .I2(n49[0]), .I3(GND_net), 
            .O(n376)) /* synthesis syn_instantiated=1 */ ;
    defparam add_18_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_23_i19_2_lut (.I0(PWMLimit[9]), .I1(n352[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5580));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i21_2_lut (.I0(PWMLimit[10]), .I1(n352[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5581));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49844_4_lut (.I0(n21_adj_5574), .I1(n19_adj_5569), .I2(n17_adj_5566), 
            .I3(n9_adj_5563), .O(n65530));
    defparam i49844_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_23_i23_2_lut (.I0(PWMLimit[11]), .I1(n352[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5582));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i15_2_lut (.I0(PWMLimit[7]), .I1(n352[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5583));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i25_2_lut (.I0(PWMLimit[12]), .I1(n352[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5584));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_16_i518_2_lut (.I0(\Kp[10] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_5233));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i6_3_lut (.I0(n130[5]), .I1(n182[5]), .I2(n181), .I3(GND_net), 
            .O(n207[5]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i6_3_lut (.I0(n207[5]), .I1(IntegralLimit[5]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[5] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49836_4_lut (.I0(n27_adj_5562), .I1(n15_adj_5561), .I2(n13_adj_5560), 
            .I3(n11_adj_5554), .O(n65522));
    defparam i49836_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_17_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5232));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_5231));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n597));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n670));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n624));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_26_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[2]));   // verilog/motorControl.v(56[22:31])
    defparam unary_minus_26_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n816));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n697));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n889));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n962));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n1035));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n1108));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i12_3_lut (.I0(n182[7]), .I1(n182[16]), .I2(n33_adj_5553), 
            .I3(GND_net), .O(n12_adj_5586));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i5_3_lut (.I0(n130[4]), .I1(n182[4]), .I2(n181), .I3(GND_net), 
            .O(n207[4]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i5_3_lut (.I0(n207[4]), .I1(IntegralLimit[4]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[4] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5229));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i14_3_lut (.I0(n130[13]), .I1(n182[13]), .I2(n181), 
            .I3(GND_net), .O(n207[13]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i14_3_lut (.I0(n207[13]), .I1(IntegralLimit[13]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[13] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n770));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n375_c));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_5228));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n594));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n667));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i10_3_lut (.I0(n182[5]), .I1(n182[6]), .I2(n13_adj_5560), 
            .I3(GND_net), .O(n10_adj_5587));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n813));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_5224));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_5223));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_5222));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_5221));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i75_2_lut (.I0(\Kp[1] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_5218));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i28_2_lut (.I0(\Kp[0] ), .I1(n55[17]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5217));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i124_2_lut (.I0(\Kp[2] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_5215));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[0]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[1]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[2]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i173_2_lut (.I0(\Kp[3] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_5213));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i222_2_lut (.I0(\Kp[4] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_5212));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i271_2_lut (.I0(\Kp[5] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_5211));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i320_2_lut (.I0(\Kp[6] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_5210));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i655_2_lut (.I0(\Kp[13] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i369_2_lut (.I0(\Kp[7] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_5209));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i418_2_lut (.I0(\Kp[8] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_5208));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i704_2_lut (.I0(\Kp[14] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i467_2_lut (.I0(\Kp[9] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_5207));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i753_2_lut (.I0(\Kp[15] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i516_2_lut (.I0(\Kp[10] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_5206));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[3]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i565_2_lut (.I0(\Kp[11] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_5205));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[4]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_5565));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_5564));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_5559));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_5558));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[5]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_5556));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[6]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_5551));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_5550));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[7]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_12_i30_3_lut (.I0(n12_adj_5586), .I1(n182[17]), .I2(n35_adj_5552), 
            .I3(GND_net), .O(n30_adj_5588));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_13_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[8]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[9]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_5546));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i4_3_lut (.I0(n130[3]), .I1(n182[3]), .I2(n181), .I3(GND_net), 
            .O(n207[3]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n630_adj_5545));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i4_3_lut (.I0(n207[3]), .I1(IntegralLimit[3]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[3] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_5204));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5203));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i61_2_lut (.I0(\Kp[1] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n89_adj_5544));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i14_2_lut (.I0(\Kp[0] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_5543));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i73_2_lut (.I0(\Kp[1] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_5542));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i26_2_lut (.I0(\Kp[0] ), .I1(n55[16]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_5541));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i110_2_lut (.I0(\Kp[2] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n162_adj_5540));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i159_2_lut (.I0(\Kp[3] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_5539));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i122_2_lut (.I0(\Kp[2] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_5538));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[10]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i208_2_lut (.I0(\Kp[4] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_5536));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_5202));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_5201));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i171_2_lut (.I0(\Kp[3] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_5535));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i257_2_lut (.I0(\Kp[5] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n381_adj_5534));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i306_2_lut (.I0(\Kp[6] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_5533));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_5200));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[11]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i355_2_lut (.I0(\Kp[7] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n527_adj_5531));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i220_2_lut (.I0(\Kp[4] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_5530));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[12]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i269_2_lut (.I0(\Kp[5] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_5528));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i318_2_lut (.I0(\Kp[6] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_5527));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_5199));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_5198));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[13]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i51_2_lut (.I0(\Kp[1] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_5197));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i4_2_lut (.I0(\Kp[0] ), .I1(n55[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_5196));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_5195));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i367_2_lut (.I0(\Kp[7] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_5525));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i404_2_lut (.I0(\Kp[8] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n600_adj_5524));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i453_2_lut (.I0(\Kp[9] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n673_adj_5523));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i502_2_lut (.I0(\Kp[10] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_5522));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i416_2_lut (.I0(\Kp[8] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_5521));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i465_2_lut (.I0(\Kp[9] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_5520));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50768_4_lut (.I0(n13_adj_5560), .I1(n11_adj_5554), .I2(n9_adj_5563), 
            .I3(n65576), .O(n66454));
    defparam i50768_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 unary_minus_13_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[14]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i551_2_lut (.I0(\Kp[11] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_5518));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i514_2_lut (.I0(\Kp[10] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_5517));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[15]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i563_2_lut (.I0(\Kp[11] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_5515));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50762_4_lut (.I0(n19_adj_5569), .I1(n17_adj_5566), .I2(n15_adj_5561), 
            .I3(n66454), .O(n66448));
    defparam i50762_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_16_i612_2_lut (.I0(\Kp[12] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_5514));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i600_2_lut (.I0(\Kp[12] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_5513));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[16]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i100_2_lut (.I0(\Kp[2] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_5194));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i149_2_lut (.I0(\Kp[3] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_5192));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n591_adj_5191));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n664_adj_5190));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_5189));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n810_adj_5188));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n883_adj_5187));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n956_adj_5186));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_5185));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n1102_adj_5184));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i3_3_lut (.I0(n130[2]), .I1(n182[2]), .I2(n181), .I3(GND_net), 
            .O(n207[2]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i3_3_lut (.I0(n207[2]), .I1(IntegralLimit[2]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[2] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i649_2_lut (.I0(\Kp[13] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_5511));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i698_2_lut (.I0(\Kp[14] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1038_adj_5510));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5178));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_5176));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_5175));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i747_2_lut (.I0(\Kp[15] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1111_adj_5509));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[17]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i198_2_lut (.I0(\Kp[4] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_5174));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_5173));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i247_2_lut (.I0(\Kp[5] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_5172));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n588));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[18]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n661));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n807));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n880));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i296_2_lut (.I0(\Kp[6] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_5166));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n953));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52181_4_lut (.I0(n25_adj_5448), .I1(n23_adj_5413), .I2(n21_adj_5574), 
            .I3(n66448), .O(n67867));
    defparam i52181_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_13_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[19]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[20]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[21]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i49827_2_lut_4_lut (.I0(n130[16]), .I1(n182[16]), .I2(n130[7]), 
            .I3(n182[7]), .O(n65513));
    defparam i49827_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i504_2_lut (.I0(\Kp[10] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_13_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[22]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_13_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n65[23]));   // verilog/motorControl.v(49[22:36])
    defparam unary_minus_13_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i59_2_lut (.I0(\Kp[1] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_5500));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n1026));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n1099));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i12_2_lut (.I0(\Kp[0] ), .I1(n55[9]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5499));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i18_3_lut (.I0(n130[17]), .I1(n182[17]), .I2(n181), 
            .I3(GND_net), .O(n214));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_5165));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23214_1_lut (.I0(n376), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37174));   // verilog/motorControl.v(51[18:38])
    defparam i23214_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i1_1_lut (.I0(deadband[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[0]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i108_2_lut (.I0(\Kp[2] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n159_adj_5496));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i157_2_lut (.I0(\Kp[3] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n232_adj_5495));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i206_2_lut (.I0(\Kp[4] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_5494));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i255_2_lut (.I0(\Kp[5] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_5493));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i304_2_lut (.I0(\Kp[6] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_5492));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i353_2_lut (.I0(\Kp[7] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n524_adj_5491));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i2_1_lut (.I0(deadband[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[1]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i402_2_lut (.I0(\Kp[8] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n597_adj_5489));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i3_1_lut (.I0(deadband[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[2]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i451_2_lut (.I0(\Kp[9] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_5487));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i500_2_lut (.I0(\Kp[10] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_5486));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i4_1_lut (.I0(deadband[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[3]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i5_1_lut (.I0(deadband[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[4]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i549_2_lut (.I0(\Kp[11] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_5482));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i598_2_lut (.I0(\Kp[12] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_5481));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i647_2_lut (.I0(\Kp[13] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n962_adj_5480));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i6_1_lut (.I0(deadband[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[5]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i345_2_lut (.I0(\Kp[7] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n512_adj_5159));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i2_3_lut (.I0(n130[1]), .I1(n182[1]), .I2(n181), .I3(GND_net), 
            .O(n207[1]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i2_3_lut (.I0(n207[1]), .I1(IntegralLimit[1]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[1] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_5158));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35120_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[22] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3715[21] ), .I3(\Ki[1] ), 
            .O(n20229[0]));   // verilog/motorControl.v(51[27:38])
    defparam i35120_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_16_i696_2_lut (.I0(\Kp[14] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_5478));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i394_2_lut (.I0(\Kp[8] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_5157));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i745_2_lut (.I0(\Kp[15] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_5477));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i51533_4_lut (.I0(n31_adj_5412), .I1(n29_adj_5411), .I2(n27_adj_5562), 
            .I3(n67867), .O(n67219));
    defparam i51533_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 unary_minus_20_inv_0_i7_1_lut (.I0(deadband[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[6]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i443_2_lut (.I0(\Kp[9] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_5155));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i8_1_lut (.I0(deadband[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[7]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_17_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35122_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[22] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3715[21] ), .I3(\Ki[1] ), 
            .O(n49008));   // verilog/motorControl.v(51[27:38])
    defparam i35122_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 unary_minus_20_inv_0_i9_1_lut (.I0(deadband[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[8]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i10_1_lut (.I0(deadband[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[9]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i11_1_lut (.I0(deadband[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[10]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i12_1_lut (.I0(deadband[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[11]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i13_1_lut (.I0(deadband[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[12]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i71_2_lut (.I0(\Kp[1] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_5466));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i24_2_lut (.I0(\Kp[0] ), .I1(n55[15]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5465));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i553_2_lut (.I0(\Kp[11] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n822));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35170_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[21] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3715[20] ), .I3(\Ki[1] ), 
            .O(n20220[0]));   // verilog/motorControl.v(51[27:38])
    defparam i35170_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_16_i602_2_lut (.I0(\Kp[12] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35172_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[21] ), 
            .I2(\PID_CONTROLLER.integral_23__N_3715[20] ), .I3(\Ki[1] ), 
            .O(n49059));   // verilog/motorControl.v(51[27:38])
    defparam i35172_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 unary_minus_20_inv_0_i14_1_lut (.I0(deadband[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[13]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i15_1_lut (.I0(deadband[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[14]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_3_lut (.I0(counter[19]), .I1(counter[24]), .I2(counter[29]), 
            .I3(GND_net), .O(n14_adj_5590));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut (.I0(counter[28]), .I1(counter[27]), .I2(counter[16]), 
            .I3(counter[30]), .O(n15_adj_5591));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1801 (.I0(counter[2]), .I1(counter[0]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_5592));
    defparam i1_2_lut_adj_1801.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(counter[4]), .I1(counter[6]), .I2(counter[1]), 
            .I3(counter[3]), .O(n12_adj_5593));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4912_4_lut (.I0(counter[5]), .I1(counter[7]), .I2(n12_adj_5593), 
            .I3(n8_adj_5592), .O(n16_adj_5594));
    defparam i4912_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i4_4_lut (.I0(counter[13]), .I1(counter[9]), .I2(counter[10]), 
            .I3(counter[11]), .O(n10_adj_5595));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut_adj_1802 (.I0(counter[12]), .I1(n10_adj_5595), .I2(n16_adj_5594), 
            .I3(counter[8]), .O(n59568));
    defparam i5_4_lut_adj_1802.LUT_INIT = 16'h8880;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5591), .I1(counter[20]), .I2(n14_adj_5590), 
            .I3(counter[14]), .O(n59846));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1803 (.I0(counter[23]), .I1(n59846), .I2(n59568), 
            .I3(counter[17]), .O(n16_adj_5596));
    defparam i6_4_lut_adj_1803.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut (.I0(counter[15]), .I1(counter[25]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5597));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut (.I0(counter[21]), .I1(counter[22]), .I2(counter[26]), 
            .I3(counter[18]), .O(n17_adj_5598));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i28949_4_lut (.I0(n17_adj_5598), .I1(counter[31]), .I2(n15_adj_5597), 
            .I3(n16_adj_5596), .O(counter_31__N_3714));   // verilog/motorControl.v(26[8:41])
    defparam i28949_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 mult_16_i492_2_lut (.I0(\Kp[10] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_5153));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i541_2_lut (.I0(\Kp[11] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_5151));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i651_2_lut (.I0(\Kp[13] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_5150));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_5149));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i700_2_lut (.I0(\Kp[14] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52425_4_lut (.I0(n37_adj_5409), .I1(n35_adj_5552), .I2(n33_adj_5553), 
            .I3(n67219), .O(n68111));
    defparam i52425_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_16_i749_2_lut (.I0(\Kp[15] ), .I1(n55[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i120_2_lut (.I0(\Kp[2] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_5462));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i16_3_lut (.I0(n182[9]), .I1(n182[21]), .I2(n43_adj_5119), 
            .I3(GND_net), .O(n16_adj_5599));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_20_inv_0_i16_1_lut (.I0(deadband[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[15]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52169_3_lut (.I0(n6_c), .I1(n182[10]), .I2(n21_adj_5574), 
            .I3(GND_net), .O(n67855));   // verilog/motorControl.v(48[21:44])
    defparam i52169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52170_3_lut (.I0(n67855), .I1(n182[11]), .I2(n23_adj_5413), 
            .I3(GND_net), .O(n67856));   // verilog/motorControl.v(48[21:44])
    defparam i52170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_5459));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i590_2_lut (.I0(\Kp[12] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_5148));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_5147));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i639_2_lut (.I0(\Kp[13] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_5145));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_5458));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i688_2_lut (.I0(\Kp[14] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_5144));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i737_2_lut (.I0(\Kp[15] ), .I1(n55[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_5143));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i169_2_lut (.I0(\Kp[3] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_5457));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_5456));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49895_2_lut_4_lut (.I0(IntegralLimit[21]), .I1(n130[21]), .I2(IntegralLimit[9]), 
            .I3(n130[9]), .O(n65581));
    defparam i49895_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_17_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_14_i17_3_lut (.I0(n130[16]), .I1(n182[16]), .I2(n181), 
            .I3(GND_net), .O(n207[16]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i218_2_lut (.I0(\Kp[4] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_5455));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i17_3_lut (.I0(n207[16]), .I1(IntegralLimit[16]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[16] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n585));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_5454));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_5453));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i65_2_lut (.I0(\Kp[1] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n95));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i17_1_lut (.I0(deadband[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[16]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i18_2_lut (.I0(\Kp[0] ), .I1(n55[12]), .I2(GND_net), 
            .I3(GND_net), .O(n26));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_5451));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i114_2_lut (.I0(\Kp[2] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i163_2_lut (.I0(\Kp[3] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n241));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n950));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_5450));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3715[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49971_2_lut_4_lut (.I0(IntegralLimit[16]), .I1(n130[16]), .I2(IntegralLimit[7]), 
            .I3(n130[7]), .O(n65657));
    defparam i49971_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_16_i212_2_lut (.I0(\Kp[4] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n314));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i261_2_lut (.I0(\Kp[5] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n387));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_12_i8_3_lut (.I0(n182[4]), .I1(n182[8]), .I2(n17_adj_5566), 
            .I3(GND_net), .O(n8_adj_5600));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35206_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n20220[0]), 
            .O(n4_adj_32));   // verilog/motorControl.v(51[27:38])
    defparam i35206_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 LessThan_12_i24_3_lut (.I0(n16_adj_5599), .I1(n182[22]), .I2(n45_adj_5120), 
            .I3(GND_net), .O(n24_adj_5604));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_17_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_5449));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i50729_4_lut (.I0(n43_adj_5119), .I1(n25_adj_5448), .I2(n23_adj_5413), 
            .I3(n65530), .O(n66415));
    defparam i50729_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_3_lut_4_lut_adj_1804 (.I0(n62), .I1(n131), .I2(n204), .I3(n20220[0]), 
            .O(n20195));   // verilog/motorControl.v(51[27:38])
    defparam i1_3_lut_4_lut_adj_1804.LUT_INIT = 16'h8778;
    SB_LUT4 unary_minus_20_inv_0_i18_1_lut (.I0(deadband[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[17]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_14_i16_3_lut (.I0(n130[15]), .I1(n182[15]), .I2(n181), 
            .I3(GND_net), .O(n207[15]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i310_2_lut (.I0(\Kp[6] ), .I1(n55[11]), .I2(GND_net), 
            .I3(GND_net), .O(n460));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_17_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n627_adj_5446));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_15_i16_3_lut (.I0(n207[15]), .I1(IntegralLimit[15]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[15] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_14_i24_3_lut (.I0(n130[23]), .I1(n182[23]), .I2(n181), 
            .I3(GND_net), .O(n207[23]));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_14_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_15_i24_3_lut (.I0(n207[23]), .I1(IntegralLimit[23]), .I2(n155), 
            .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715[23] ));   // verilog/motorControl.v(48[18] 50[12])
    defparam mux_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29444_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43349));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29444_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51605_4_lut (.I0(n24_adj_5604), .I1(n8_adj_5600), .I2(n45_adj_5120), 
            .I3(n66411), .O(n67291));   // verilog/motorControl.v(48[21:44])
    defparam i51605_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51929_3_lut (.I0(n67856), .I1(n182[12]), .I2(n25_adj_5448), 
            .I3(GND_net), .O(n67615));   // verilog/motorControl.v(48[21:44])
    defparam i51929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_12_i4_4_lut (.I0(n130[0]), .I1(n182[1]), .I2(n130[1]), 
            .I3(n182[0]), .O(n4_adj_5605));   // verilog/motorControl.v(48[21:44])
    defparam LessThan_12_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i52167_3_lut (.I0(n4_adj_5605), .I1(n182[13]), .I2(n27_adj_5562), 
            .I3(GND_net), .O(n67853));   // verilog/motorControl.v(48[21:44])
    defparam i52167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52168_3_lut (.I0(n67853), .I1(n182[14]), .I2(n29_adj_5411), 
            .I3(GND_net), .O(n67854));   // verilog/motorControl.v(48[21:44])
    defparam i52168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29324_4_lut (.I0(PWMLimit[1]), .I1(n60219), .I2(n37189), 
            .I3(n11608), .O(n51[1]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29324_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_17_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3715[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n700_adj_5444));   // verilog/motorControl.v(51[27:38])
    defparam mult_17_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i19_1_lut (.I0(deadband[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[18]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i267_2_lut (.I0(\Kp[5] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_5441));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i316_2_lut (.I0(\Kp[6] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_5440));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i365_2_lut (.I0(\Kp[7] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_5439));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i20_1_lut (.I0(deadband[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[19]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i414_2_lut (.I0(\Kp[8] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_5437));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i57_2_lut (.I0(\Kp[1] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_5436));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i10_2_lut (.I0(\Kp[0] ), .I1(n55[8]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_5435));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i21_1_lut (.I0(deadband[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[20]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i106_2_lut (.I0(\Kp[2] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_5433));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13894_3_lut (.I0(n352[2]), .I1(n432[2]), .I2(n11610), .I3(GND_net), 
            .O(n27892));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49829_4_lut (.I0(n33_adj_5553), .I1(n31_adj_5412), .I2(n29_adj_5411), 
            .I3(n65522), .O(n65515));
    defparam i49829_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52375_4_lut (.I0(n30_adj_5588), .I1(n10_adj_5587), .I2(n35_adj_5552), 
            .I3(n65513), .O(n68061));   // verilog/motorControl.v(48[21:44])
    defparam i52375_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29323_4_lut (.I0(PWMLimit[2]), .I1(n60219), .I2(n27892), 
            .I3(n11608), .O(n51[2]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29323_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_16_i155_2_lut (.I0(\Kp[3] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_5432));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13889_3_lut (.I0(n352[3]), .I1(n432[3]), .I2(n11610), .I3(GND_net), 
            .O(n27887));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29322_4_lut (.I0(PWMLimit[3]), .I1(n60219), .I2(n27887), 
            .I3(n11608), .O(n51[3]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29322_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_16_i463_2_lut (.I0(\Kp[9] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_5431));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i204_2_lut (.I0(\Kp[4] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_5430));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13884_3_lut (.I0(n352[4]), .I1(n432[4]), .I2(n11610), .I3(GND_net), 
            .O(n27882));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29321_4_lut (.I0(PWMLimit[4]), .I1(n60219), .I2(n27882), 
            .I3(n11608), .O(n51[4]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29321_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 unary_minus_20_inv_0_i22_1_lut (.I0(deadband[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[21]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_16_i512_2_lut (.I0(\Kp[10] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n761_adj_5427));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i253_2_lut (.I0(\Kp[5] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_5426));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i302_2_lut (.I0(\Kp[6] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_5425));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i561_2_lut (.I0(\Kp[11] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_5424));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i23_1_lut (.I0(deadband[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[22]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i51931_3_lut (.I0(n67854), .I1(n182[15]), .I2(n31_adj_5412), 
            .I3(GND_net), .O(n28_adj_5606));   // verilog/motorControl.v(48[21:44])
    defparam i51931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_16_i351_2_lut (.I0(\Kp[7] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_5422));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13879_3_lut (.I0(n352[5]), .I1(n432[5]), .I2(n11610), .I3(GND_net), 
            .O(n27877));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29320_4_lut (.I0(PWMLimit[5]), .I1(n60219), .I2(n27877), 
            .I3(n11608), .O(n51[5]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29320_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_16_i400_2_lut (.I0(\Kp[8] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_5421));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52525_4_lut (.I0(n28_adj_5606), .I1(n68061), .I2(n35_adj_5552), 
            .I3(n65515), .O(n68211));   // verilog/motorControl.v(48[21:44])
    defparam i52525_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_16_i449_2_lut (.I0(\Kp[9] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n667_adj_5420));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13874_3_lut (.I0(n352[6]), .I1(n432[6]), .I2(n11610), .I3(GND_net), 
            .O(n27872));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29319_4_lut (.I0(PWMLimit[6]), .I1(n60219), .I2(n27872), 
            .I3(n11608), .O(n51[6]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29319_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_16_i498_2_lut (.I0(\Kp[10] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_5419));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13869_3_lut (.I0(n352[7]), .I1(n432[7]), .I2(n11610), .I3(GND_net), 
            .O(n27867));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29318_4_lut (.I0(PWMLimit[7]), .I1(n60219), .I2(n27867), 
            .I3(n11608), .O(n51[7]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29318_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 unary_minus_20_inv_0_i24_1_lut (.I0(deadband[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n61[23]));   // verilog/motorControl.v(52[43:52])
    defparam unary_minus_20_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13864_3_lut (.I0(n352[8]), .I1(n432[8]), .I2(n11610), .I3(GND_net), 
            .O(n27862));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29317_4_lut (.I0(PWMLimit[8]), .I1(n60219), .I2(n27862), 
            .I3(n11608), .O(n51[8]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29317_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_16_i610_2_lut (.I0(\Kp[12] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_5416));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13859_3_lut (.I0(n352[9]), .I1(n432[9]), .I2(n11610), .I3(GND_net), 
            .O(n27857));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29316_4_lut (.I0(PWMLimit[9]), .I1(n60219), .I2(n27857), 
            .I3(n11608), .O(n51[9]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29316_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mult_16_i547_2_lut (.I0(\Kp[11] ), .I1(n55[7]), .I2(GND_net), 
            .I3(GND_net), .O(n813_adj_5415));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_16_i659_2_lut (.I0(\Kp[13] ), .I1(n55[14]), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_5414));   // verilog/motorControl.v(51[18:24])
    defparam mult_16_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i33_2_lut (.I0(deadband[16]), .I1(n352[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5607));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i31_2_lut (.I0(deadband[15]), .I1(n361), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5608));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i37_2_lut (.I0(deadband[18]), .I1(n352[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5609));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i35_2_lut (.I0(deadband[17]), .I1(n352[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5610));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i25_2_lut (.I0(deadband[12]), .I1(n352[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5611));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i27_2_lut (.I0(deadband[13]), .I1(n352[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5612));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i29_2_lut (.I0(deadband[14]), .I1(n352[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5613));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50497_2_lut_4_lut (.I0(n352[21]), .I1(n432[21]), .I2(n352[9]), 
            .I3(n432[9]), .O(n66183));
    defparam i50497_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_19_i21_2_lut (.I0(deadband[10]), .I1(n352[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5614));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i23_2_lut (.I0(deadband[11]), .I1(n352[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5615));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i13_2_lut (.I0(deadband[6]), .I1(n352[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5616));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i15_2_lut (.I0(deadband[7]), .I1(n352[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5617));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i17_2_lut (.I0(deadband[8]), .I1(n352[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5618));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i9_2_lut (.I0(deadband[4]), .I1(n352[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5619));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i11_2_lut (.I0(deadband[5]), .I1(n352[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5620));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i19_2_lut (.I0(deadband[9]), .I1(n352[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5621));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i43_2_lut (.I0(PWMLimit[21]), .I1(n352[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5622));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13854_3_lut (.I0(n352[10]), .I1(n432[10]), .I2(n11610), .I3(GND_net), 
            .O(n27852));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29315_4_lut (.I0(PWMLimit[10]), .I1(n60219), .I2(n27852), 
            .I3(n11608), .O(n51[10]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29315_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 LessThan_23_i41_2_lut (.I0(PWMLimit[20]), .I1(n352[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5623));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i37_2_lut (.I0(PWMLimit[18]), .I1(n352[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5624));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i39_2_lut (.I0(PWMLimit[19]), .I1(n352[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5625));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_23_i5_2_lut (.I0(PWMLimit[2]), .I1(n352[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_5626));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50582_4_lut (.I0(n11_adj_5575), .I1(n9_adj_5577), .I2(n7_adj_5579), 
            .I3(n5_adj_5626), .O(n66268));
    defparam i50582_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50578_4_lut (.I0(n17_adj_5578), .I1(n15_adj_5583), .I2(n13_adj_5576), 
            .I3(n66268), .O(n66264));
    defparam i50578_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_23_i10_3_lut (.I0(n352[5]), .I1(n352[6]), .I2(n13_adj_5576), 
            .I3(GND_net), .O(n10_adj_5627));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13849_3_lut (.I0(n352[11]), .I1(n432[11]), .I2(n11610), .I3(GND_net), 
            .O(n27847));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29314_4_lut (.I0(PWMLimit[11]), .I1(n60219), .I2(n27847), 
            .I3(n11608), .O(n51[11]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29314_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13844_3_lut (.I0(n352[12]), .I1(n432[12]), .I2(n11610), .I3(GND_net), 
            .O(n27842));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29313_4_lut (.I0(PWMLimit[12]), .I1(n60219), .I2(n27842), 
            .I3(n11608), .O(n51[12]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29313_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 LessThan_23_i12_3_lut (.I0(n10_adj_5627), .I1(n352[7]), .I2(n15_adj_5583), 
            .I3(GND_net), .O(n12_adj_5628));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i8_3_lut (.I0(n352[4]), .I1(n352[8]), .I2(n17_adj_5578), 
            .I3(GND_net), .O(n8_adj_5629));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13839_3_lut (.I0(n352[13]), .I1(n432[13]), .I2(n11610), .I3(GND_net), 
            .O(n27837));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29312_4_lut (.I0(PWMLimit[13]), .I1(n60219), .I2(n27837), 
            .I3(n11608), .O(n51[13]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29312_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13834_3_lut (.I0(n352[14]), .I1(n432[14]), .I2(n11610), .I3(GND_net), 
            .O(n27832));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29311_4_lut (.I0(PWMLimit[14]), .I1(n60219), .I2(n27832), 
            .I3(n11608), .O(n51[14]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29311_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 LessThan_23_i6_3_lut (.I0(n352[2]), .I1(n352[3]), .I2(n7_adj_5579), 
            .I3(GND_net), .O(n6_adj_5630));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13829_3_lut (.I0(n361), .I1(n432[15]), .I2(n11610), .I3(GND_net), 
            .O(n27827));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_23_i16_3_lut (.I0(n8_adj_5629), .I1(n352[9]), .I2(n19_adj_5580), 
            .I3(GND_net), .O(n16_adj_5631));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29310_4_lut (.I0(PWMLimit[15]), .I1(n60219), .I2(n27827), 
            .I3(n11608), .O(n51[15]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29310_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i52383_4_lut (.I0(n16_adj_5631), .I1(n6_adj_5630), .I2(n19_adj_5580), 
            .I3(n66260), .O(n68069));   // verilog/motorControl.v(53[14:29])
    defparam i52383_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52384_3_lut (.I0(n68069), .I1(n352[10]), .I2(n21_adj_5581), 
            .I3(GND_net), .O(n68070));   // verilog/motorControl.v(53[14:29])
    defparam i52384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52263_3_lut (.I0(n68070), .I1(n352[11]), .I2(n23_adj_5582), 
            .I3(GND_net), .O(n67949));   // verilog/motorControl.v(53[14:29])
    defparam i52263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52113_4_lut (.I0(n23_adj_5582), .I1(n21_adj_5581), .I2(n19_adj_5580), 
            .I3(n66264), .O(n67799));
    defparam i52113_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13824_3_lut (.I0(n352[16]), .I1(n432[16]), .I2(n11610), .I3(GND_net), 
            .O(n27822));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29309_4_lut (.I0(PWMLimit[16]), .I1(n60219), .I2(n27822), 
            .I3(n11608), .O(n51[16]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29309_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i52161_4_lut (.I0(n12_adj_5628), .I1(n4_adj_33), .I2(n15_adj_5583), 
            .I3(n66266), .O(n67847));   // verilog/motorControl.v(53[14:29])
    defparam i52161_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50915_3_lut (.I0(n67949), .I1(n352[12]), .I2(n25_adj_5584), 
            .I3(GND_net), .O(n66601));   // verilog/motorControl.v(53[14:29])
    defparam i50915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52389_4_lut (.I0(n66601), .I1(n67847), .I2(n25_adj_5584), 
            .I3(n67799), .O(n68075));   // verilog/motorControl.v(53[14:29])
    defparam i52389_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52390_3_lut (.I0(n68075), .I1(n352[13]), .I2(PWMLimit[13]), 
            .I3(GND_net), .O(n68076));   // verilog/motorControl.v(53[14:29])
    defparam i52390_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52241_3_lut (.I0(n68076), .I1(n352[14]), .I2(PWMLimit[14]), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(53[14:29])
    defparam i52241_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i13819_3_lut (.I0(n352[17]), .I1(n432[17]), .I2(n11610), .I3(GND_net), 
            .O(n27817));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29308_4_lut (.I0(PWMLimit[17]), .I1(n60219), .I2(n27817), 
            .I3(n11608), .O(n51[17]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29308_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13814_3_lut (.I0(n352[18]), .I1(n432[18]), .I2(n11610), .I3(GND_net), 
            .O(n27812));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29307_4_lut (.I0(PWMLimit[18]), .I1(n60219), .I2(n27812), 
            .I3(n11608), .O(n51[18]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29307_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13809_3_lut (.I0(n352[19]), .I1(n432[19]), .I2(n11610), .I3(GND_net), 
            .O(n27807));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29306_4_lut (.I0(PWMLimit[19]), .I1(n60219), .I2(n27807), 
            .I3(n11608), .O(n51[19]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29306_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13804_3_lut (.I0(n352[20]), .I1(n432[20]), .I2(n11610), .I3(GND_net), 
            .O(n27802));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29305_4_lut (.I0(PWMLimit[20]), .I1(n60219), .I2(n27802), 
            .I3(n11608), .O(n51[20]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29305_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i51976_3_lut (.I0(n32), .I1(n352[19]), .I2(n39_adj_5625), 
            .I3(GND_net), .O(n67662));   // verilog/motorControl.v(53[14:29])
    defparam i51976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51977_3_lut (.I0(n67662), .I1(n352[20]), .I2(n41_adj_5623), 
            .I3(GND_net), .O(n67663));   // verilog/motorControl.v(53[14:29])
    defparam i51977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35043_2_lut_3_lut (.I0(\Kp[0] ), .I1(n55[23]), .I2(\Kp[1] ), 
            .I3(GND_net), .O(n48918));   // verilog/motorControl.v(51[18:24])
    defparam i35043_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i13799_3_lut (.I0(n352[21]), .I1(n432[21]), .I2(n11610), .I3(GND_net), 
            .O(n27797));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29304_4_lut (.I0(PWMLimit[21]), .I1(n60219), .I2(n27797), 
            .I3(n11608), .O(n51[21]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29304_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i13794_3_lut (.I0(n352[22]), .I1(n432[22]), .I2(n11610), .I3(GND_net), 
            .O(n27792));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29303_4_lut (.I0(PWMLimit[22]), .I1(n60219), .I2(n27792), 
            .I3(n11608), .O(n51[22]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29303_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i2_2_lut_3_lut (.I0(\Kp[2] ), .I1(\Kp[0] ), .I2(\Kp[1] ), 
            .I3(GND_net), .O(n60074));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i51425_4_lut (.I0(n41_adj_5623), .I1(n39_adj_5625), .I2(n37_adj_5624), 
            .I3(n66246), .O(n67111));
    defparam i51425_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51936_3_lut (.I0(n34_adj_5635), .I1(n352[18]), .I2(n37_adj_5624), 
            .I3(GND_net), .O(n67622));   // verilog/motorControl.v(53[14:29])
    defparam i51936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50917_3_lut (.I0(n67663), .I1(n352[21]), .I2(n43_adj_5622), 
            .I3(GND_net), .O(n66603));   // verilog/motorControl.v(53[14:29])
    defparam i50917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51974_4_lut (.I0(n66603), .I1(n67622), .I2(n43_adj_5622), 
            .I3(n67111), .O(n67660));   // verilog/motorControl.v(53[14:29])
    defparam i51974_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51975_3_lut (.I0(n67660), .I1(n352[22]), .I2(PWMLimit[22]), 
            .I3(GND_net), .O(n67661));   // verilog/motorControl.v(53[14:29])
    defparam i51975_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_23_i48_3_lut (.I0(n67661), .I1(PWMLimit[23]), .I2(n352[23]), 
            .I3(GND_net), .O(n405));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50670_4_lut (.I0(n352[6]), .I1(n352[5]), .I2(n63[6]), .I3(n63[5]), 
            .O(n66356));
    defparam i50670_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i51485_3_lut (.I0(n352[7]), .I1(n66356), .I2(n63[7]), .I3(GND_net), 
            .O(n67171));
    defparam i51485_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 LessThan_21_i27_rep_81_2_lut (.I0(n352[13]), .I1(n63[13]), .I2(GND_net), 
            .I3(GND_net), .O(n69591));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i27_rep_81_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51473_4_lut (.I0(n352[14]), .I1(n69591), .I2(n63[14]), .I3(n67171), 
            .O(n67159));
    defparam i51473_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_21_i31_rep_75_2_lut (.I0(n361), .I1(n63[15]), .I2(GND_net), 
            .I3(GND_net), .O(n69585));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i31_rep_75_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_21_i12_3_lut (.I0(n63[7]), .I1(n63[16]), .I2(n352[16]), 
            .I3(GND_net), .O(n12_adj_5636));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50634_4_lut (.I0(n352[16]), .I1(n352[7]), .I2(n63[16]), .I3(n63[7]), 
            .O(n66320));
    defparam i50634_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_21_i35_rep_100_2_lut (.I0(n352[17]), .I1(n63[17]), 
            .I2(GND_net), .I3(GND_net), .O(n69610));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i35_rep_100_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_21_i10_3_lut (.I0(n63[5]), .I1(n63[6]), .I2(n352[6]), 
            .I3(GND_net), .O(n10_adj_5637));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_21_i30_3_lut (.I0(n12_adj_5636), .I1(n63[17]), .I2(n352[17]), 
            .I3(GND_net), .O(n30_adj_5638));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50666_4_lut (.I0(n352[8]), .I1(n352[4]), .I2(n63[8]), .I3(n63[4]), 
            .O(n66352));
    defparam i50666_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i51481_3_lut (.I0(n352[9]), .I1(n66352), .I2(n63[9]), .I3(GND_net), 
            .O(n67167));
    defparam i51481_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 LessThan_21_i21_rep_94_2_lut (.I0(n352[10]), .I1(n63[10]), .I2(GND_net), 
            .I3(GND_net), .O(n69604));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i21_rep_94_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51479_4_lut (.I0(n352[11]), .I1(n69604), .I2(n63[11]), .I3(n67167), 
            .O(n67165));
    defparam i51479_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_21_i25_rep_89_2_lut (.I0(n352[12]), .I1(n63[12]), .I2(GND_net), 
            .I3(GND_net), .O(n69599));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i25_rep_89_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_21_i16_3_lut (.I0(n63[9]), .I1(n63[21]), .I2(n352[21]), 
            .I3(GND_net), .O(n16_adj_5639));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50592_4_lut (.I0(n352[21]), .I1(n352[9]), .I2(n63[21]), .I3(n63[9]), 
            .O(n66278));
    defparam i50592_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_21_i8_3_lut (.I0(n63[4]), .I1(n63[8]), .I2(n352[8]), 
            .I3(GND_net), .O(n8_adj_5640));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_21_i24_3_lut (.I0(n16_adj_5639), .I1(n63[22]), .I2(n352[22]), 
            .I3(GND_net), .O(n24_adj_5641));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50675_4_lut (.I0(n352[3]), .I1(n352[2]), .I2(n63[3]), .I3(n63[2]), 
            .O(n66361));
    defparam i50675_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_21_i9_rep_120_2_lut (.I0(n352[4]), .I1(n63[4]), .I2(GND_net), 
            .I3(GND_net), .O(n69630));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i9_rep_120_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50672_4_lut (.I0(n352[5]), .I1(n69630), .I2(n63[5]), .I3(n66361), 
            .O(n66358));
    defparam i50672_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_21_i13_rep_113_2_lut (.I0(n352[6]), .I1(n63[6]), .I2(GND_net), 
            .I3(GND_net), .O(n69623));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i13_rep_113_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50543_3_lut_4_lut (.I0(n352[3]), .I1(n432[3]), .I2(n432[2]), 
            .I3(n352[2]), .O(n66229));   // verilog/motorControl.v(55[23:39])
    defparam i50543_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51845_4_lut (.I0(n352[7]), .I1(n69623), .I2(n63[7]), .I3(n66358), 
            .O(n67531));
    defparam i51845_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_21_i17_rep_116_2_lut (.I0(n352[8]), .I1(n63[8]), .I2(GND_net), 
            .I3(GND_net), .O(n69626));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i17_rep_116_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51483_4_lut (.I0(n352[9]), .I1(n69626), .I2(n63[9]), .I3(n67531), 
            .O(n67169));
    defparam i51483_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_25_i6_3_lut_3_lut (.I0(n352[3]), .I1(n432[3]), .I2(n432[2]), 
            .I3(GND_net), .O(n6_adj_5141));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i52119_4_lut (.I0(n352[11]), .I1(n69604), .I2(n63[11]), .I3(n67169), 
            .O(n67805));
    defparam i52119_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i50651_4_lut (.I0(n352[13]), .I1(n69599), .I2(n63[13]), .I3(n67805), 
            .O(n66337));
    defparam i50651_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_21_i29_rep_79_2_lut (.I0(n352[14]), .I1(n63[14]), .I2(GND_net), 
            .I3(GND_net), .O(n69589));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i29_rep_79_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51839_4_lut (.I0(n361), .I1(n69589), .I2(n63[15]), .I3(n66337), 
            .O(n67525));
    defparam i51839_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_21_i33_rep_105_2_lut (.I0(n352[16]), .I1(n63[16]), 
            .I2(GND_net), .I3(GND_net), .O(n69615));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i33_rep_105_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52381_4_lut (.I0(n352[17]), .I1(n69615), .I2(n63[17]), .I3(n67525), 
            .O(n68067));
    defparam i52381_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_21_i37_rep_70_2_lut (.I0(n352[18]), .I1(n63[18]), .I2(GND_net), 
            .I3(GND_net), .O(n69580));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i37_rep_70_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52574_4_lut (.I0(n352[19]), .I1(n69580), .I2(n63[19]), .I3(n68067), 
            .O(n68260));
    defparam i52574_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_21_i41_rep_67_2_lut (.I0(n352[20]), .I1(n63[20]), .I2(GND_net), 
            .I3(GND_net), .O(n69577));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i41_rep_67_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i10_3_lut (.I0(n352[5]), .I1(n352[9]), .I2(n19_adj_5621), 
            .I3(GND_net), .O(n10_adj_5642));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51519_4_lut (.I0(n11_adj_5620), .I1(n9_adj_5619), .I2(deadband[3]), 
            .I3(n352[3]), .O(n67205));
    defparam i51519_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i51859_4_lut (.I0(n17_adj_5618), .I1(n15_adj_5617), .I2(n13_adj_5616), 
            .I3(n67205), .O(n67545));
    defparam i51859_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50517_2_lut_4_lut (.I0(n352[16]), .I1(n432[16]), .I2(n352[7]), 
            .I3(n432[7]), .O(n66203));
    defparam i50517_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51857_4_lut (.I0(n23_adj_5615), .I1(n21_adj_5614), .I2(n19_adj_5621), 
            .I3(n67545), .O(n67543));
    defparam i51857_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50705_4_lut (.I0(n29_adj_5613), .I1(n27_adj_5612), .I2(n25_adj_5611), 
            .I3(n67543), .O(n66391));
    defparam i50705_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50002_4_lut (.I0(deadband[1]), .I1(n376), .I2(n375), .I3(deadband[0]), 
            .O(n65316));   // verilog/motorControl.v(52[12:29])
    defparam i50002_4_lut.LUT_INIT = 16'h50d4;
    SB_LUT4 LessThan_19_i6_3_lut (.I0(n65316), .I1(n352[2]), .I2(deadband[2]), 
            .I3(GND_net), .O(n6_adj_5643));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51994_3_lut (.I0(n6_adj_5643), .I1(n352[14]), .I2(n29_adj_5613), 
            .I3(GND_net), .O(n67680));   // verilog/motorControl.v(52[12:29])
    defparam i51994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i14_3_lut (.I0(n352[8]), .I1(n352[17]), .I2(n35_adj_5610), 
            .I3(GND_net), .O(n14_adj_5644));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i12_3_lut (.I0(n352[6]), .I1(n352[7]), .I2(n15_adj_5617), 
            .I3(GND_net), .O(n12_adj_5645));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i32_3_lut (.I0(n14_adj_5644), .I1(n352[18]), .I2(n37_adj_5609), 
            .I3(GND_net), .O(n32_adj_5646));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50702_4_lut (.I0(n29_adj_5613), .I1(n17_adj_5618), .I2(n15_adj_5617), 
            .I3(n13_adj_5616), .O(n66388));
    defparam i50702_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51995_3_lut (.I0(n67680), .I1(n361), .I2(n31_adj_5608), .I3(GND_net), 
            .O(n67681));   // verilog/motorControl.v(52[12:29])
    defparam i51995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50698_4_lut (.I0(n35_adj_5610), .I1(n33_adj_5607), .I2(n31_adj_5608), 
            .I3(n66388), .O(n66384));
    defparam i50698_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52377_4_lut (.I0(n32_adj_5646), .I1(n12_adj_5645), .I2(n37_adj_5609), 
            .I3(n66382), .O(n68063));   // verilog/motorControl.v(52[12:29])
    defparam i52377_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50895_3_lut (.I0(n67681), .I1(n352[16]), .I2(n33_adj_5607), 
            .I3(GND_net), .O(n66581));   // verilog/motorControl.v(52[12:29])
    defparam i50895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_21_i6_3_lut (.I0(n63[2]), .I1(n63[3]), .I2(n352[3]), 
            .I3(GND_net), .O(n6_adj_5647));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51990_3_lut (.I0(n6_adj_5647), .I1(n63[10]), .I2(n352[10]), 
            .I3(GND_net), .O(n67676));   // verilog/motorControl.v(52[33:53])
    defparam i51990_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51991_3_lut (.I0(n67676), .I1(n63[11]), .I2(n352[11]), .I3(GND_net), 
            .O(n67677));   // verilog/motorControl.v(52[33:53])
    defparam i51991_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51984_3_lut (.I0(n4_adj_34), .I1(n63[13]), .I2(n352[13]), 
            .I3(GND_net), .O(n67670));   // verilog/motorControl.v(52[33:53])
    defparam i51984_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51985_3_lut (.I0(n67670), .I1(n63[14]), .I2(n352[14]), .I3(GND_net), 
            .O(n67671));   // verilog/motorControl.v(52[33:53])
    defparam i51985_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50636_4_lut (.I0(n352[16]), .I1(n69585), .I2(n63[16]), .I3(n67159), 
            .O(n66322));
    defparam i50636_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i52379_4_lut (.I0(n30_adj_5638), .I1(n10_adj_5637), .I2(n69610), 
            .I3(n66320), .O(n68065));   // verilog/motorControl.v(52[33:53])
    defparam i52379_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50905_3_lut (.I0(n67671), .I1(n63[15]), .I2(n361), .I3(GND_net), 
            .O(n66591));   // verilog/motorControl.v(52[33:53])
    defparam i50905_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52559_4_lut (.I0(n66591), .I1(n68065), .I2(n69610), .I3(n66322), 
            .O(n68245));   // verilog/motorControl.v(52[33:53])
    defparam i52559_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52560_3_lut (.I0(n68245), .I1(n63[18]), .I2(n352[18]), .I3(GND_net), 
            .O(n68246));   // verilog/motorControl.v(52[33:53])
    defparam i52560_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52522_3_lut (.I0(n68246), .I1(n63[19]), .I2(n352[19]), .I3(GND_net), 
            .O(n68208));   // verilog/motorControl.v(52[33:53])
    defparam i52522_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50596_4_lut (.I0(n352[21]), .I1(n69599), .I2(n63[21]), .I3(n67165), 
            .O(n66282));
    defparam i50596_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_21_i45_rep_64_2_lut (.I0(n352[22]), .I1(n63[22]), .I2(GND_net), 
            .I3(GND_net), .O(n69574));   // verilog/motorControl.v(52[33:53])
    defparam LessThan_21_i45_rep_64_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51609_4_lut (.I0(n24_adj_5641), .I1(n8_adj_5640), .I2(n69574), 
            .I3(n66278), .O(n67295));   // verilog/motorControl.v(52[33:53])
    defparam i51609_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50903_3_lut (.I0(n67677), .I1(n63[12]), .I2(n352[12]), .I3(GND_net), 
            .O(n66589));   // verilog/motorControl.v(52[33:53])
    defparam i50903_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50603_4_lut (.I0(n352[21]), .I1(n69577), .I2(n63[21]), .I3(n68260), 
            .O(n66289));
    defparam i50603_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i52238_4_lut (.I0(n66589), .I1(n67295), .I2(n69574), .I3(n66282), 
            .O(n67924));   // verilog/motorControl.v(52[33:53])
    defparam i52238_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i50911_3_lut (.I0(n68208), .I1(n63[20]), .I2(n352[20]), .I3(GND_net), 
            .O(n66597));   // verilog/motorControl.v(52[33:53])
    defparam i50911_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_19_i8_3_lut (.I0(n352[3]), .I1(n352[4]), .I2(n9_adj_5619), 
            .I3(GND_net), .O(n8_adj_5649));   // verilog/motorControl.v(52[12:29])
    defparam LessThan_19_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51996_3_lut (.I0(n8_adj_5649), .I1(n352[11]), .I2(n23_adj_5615), 
            .I3(GND_net), .O(n67682));   // verilog/motorControl.v(52[12:29])
    defparam i51996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51997_3_lut (.I0(n67682), .I1(n352[12]), .I2(n25_adj_5611), 
            .I3(GND_net), .O(n67683));   // verilog/motorControl.v(52[12:29])
    defparam i51997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51509_4_lut (.I0(n25_adj_5611), .I1(n23_adj_5615), .I2(n21_adj_5614), 
            .I3(n66398), .O(n67195));
    defparam i51509_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51607_3_lut (.I0(n10_adj_5642), .I1(n352[10]), .I2(n21_adj_5614), 
            .I3(GND_net), .O(n67293));   // verilog/motorControl.v(52[12:29])
    defparam i51607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50893_3_lut (.I0(n67683), .I1(n352[13]), .I2(n27_adj_5612), 
            .I3(GND_net), .O(n66579));   // verilog/motorControl.v(52[12:29])
    defparam i50893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52125_4_lut (.I0(n35_adj_5610), .I1(n33_adj_5607), .I2(n31_adj_5608), 
            .I3(n66391), .O(n67811));
    defparam i52125_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52557_4_lut (.I0(n66581), .I1(n68063), .I2(n37_adj_5609), 
            .I3(n66384), .O(n68243));   // verilog/motorControl.v(52[12:29])
    defparam i52557_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52165_4_lut (.I0(n66579), .I1(n67293), .I2(n27_adj_5612), 
            .I3(n67195), .O(n67851));   // verilog/motorControl.v(52[12:29])
    defparam i52165_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52621_4_lut (.I0(n67851), .I1(n68243), .I2(n37_adj_5609), 
            .I3(n67811), .O(n68307));   // verilog/motorControl.v(52[12:29])
    defparam i52621_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52622_3_lut (.I0(n68307), .I1(n352[19]), .I2(deadband[19]), 
            .I3(GND_net), .O(n68308));   // verilog/motorControl.v(52[12:29])
    defparam i52622_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52468_3_lut (.I0(n68308), .I1(n352[20]), .I2(deadband[20]), 
            .I3(GND_net), .O(n68154));   // verilog/motorControl.v(52[12:29])
    defparam i52468_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52391_3_lut (.I0(n68154), .I1(n352[21]), .I2(deadband[21]), 
            .I3(GND_net), .O(n68077));   // verilog/motorControl.v(52[12:29])
    defparam i52391_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52392_3_lut (.I0(n68077), .I1(n352[22]), .I2(deadband[22]), 
            .I3(GND_net), .O(n68078));   // verilog/motorControl.v(52[12:29])
    defparam i52392_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52437_4_lut (.I0(n66597), .I1(n67924), .I2(n69574), .I3(n66289), 
            .O(n68123));   // verilog/motorControl.v(52[33:53])
    defparam i52437_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1805 (.I0(n68078), .I1(control_update), .I2(deadband[23]), 
            .I3(n352[23]), .O(n61858));
    defparam i1_4_lut_adj_1805.LUT_INIT = 16'h4c04;
    SB_LUT4 i1_4_lut_adj_1806 (.I0(n61858), .I1(n68123), .I2(n352[23]), 
            .I3(n47_adj_5417), .O(n60219));
    defparam i1_4_lut_adj_1806.LUT_INIT = 16'h0a22;
    SB_LUT4 i13789_3_lut (.I0(n352[23]), .I1(n432[23]), .I2(n11610), .I3(GND_net), 
            .O(n27787));   // verilog/motorControl.v(41[14] 62[8])
    defparam i13789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29302_4_lut (.I0(PWMLimit[23]), .I1(n60219), .I2(n27787), 
            .I3(n11608), .O(n51[23]));   // verilog/motorControl.v(41[14] 62[8])
    defparam i29302_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i35193_2_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3715[20] ), 
            .I2(n36694), .I3(\Ki[1] ), .O(n20196));   // verilog/motorControl.v(51[27:38])
    defparam i35193_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 LessThan_25_i41_2_lut (.I0(n352[20]), .I1(n432[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5226));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_25_i39_2_lut (.I0(n352[19]), .I1(n432[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5225));   // verilog/motorControl.v(55[23:39])
    defparam LessThan_25_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i52526_3_lut (.I0(n68211), .I1(n182[18]), .I2(n37_adj_5409), 
            .I3(GND_net), .O(n68212));   // verilog/motorControl.v(48[21:44])
    defparam i52526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50560_3_lut_4_lut (.I0(PWMLimit[17]), .I1(n352[17]), .I2(n352[16]), 
            .I3(PWMLimit[16]), .O(n66246));   // verilog/motorControl.v(53[14:29])
    defparam i50560_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_23_i34_3_lut_3_lut (.I0(PWMLimit[17]), .I1(n352[17]), 
            .I2(n352[16]), .I3(GND_net), .O(n34_adj_5635));   // verilog/motorControl.v(53[14:29])
    defparam LessThan_23_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1) 
//

module \quadrature_decoder(1)  (b_prev, GND_net, a_new, position_31__N_3827, 
            ENCODER1_B_N_keep, n1779, ENCODER1_A_N_keep, n29704, n1784, 
            n1824, n1786, n1788, n1790, n1792, n1794, n1796, \encoder1_position[25] , 
            \encoder1_position[24] , \encoder1_position[23] , \encoder1_position[22] , 
            \encoder1_position[21] , \encoder1_position[20] , \encoder1_position[19] , 
            \encoder1_position[18] , \encoder1_position[17] , \encoder1_position[16] , 
            \encoder1_position[15] , \encoder1_position[14] , \encoder1_position[13] , 
            \encoder1_position[12] , \encoder1_position[11] , \encoder1_position[10] , 
            \encoder1_position[9] , \encoder1_position[8] , \encoder1_position[7] , 
            \encoder1_position[6] , \encoder1_position[5] , \encoder1_position[4] , 
            \encoder1_position[3] , \encoder1_position[2] , n1822, VCC_net) /* synthesis lattice_noprune=1 */ ;
    output b_prev;
    input GND_net;
    output [1:0]a_new;
    output position_31__N_3827;
    input ENCODER1_B_N_keep;
    input n1779;
    input ENCODER1_A_N_keep;
    input n29704;
    output n1784;
    output n1824;
    output n1786;
    output n1788;
    output n1790;
    output n1792;
    output n1794;
    output n1796;
    output \encoder1_position[25] ;
    output \encoder1_position[24] ;
    output \encoder1_position[23] ;
    output \encoder1_position[22] ;
    output \encoder1_position[21] ;
    output \encoder1_position[20] ;
    output \encoder1_position[19] ;
    output \encoder1_position[18] ;
    output \encoder1_position[17] ;
    output \encoder1_position[16] ;
    output \encoder1_position[15] ;
    output \encoder1_position[14] ;
    output \encoder1_position[13] ;
    output \encoder1_position[12] ;
    output \encoder1_position[11] ;
    output \encoder1_position[10] ;
    output \encoder1_position[9] ;
    output \encoder1_position[8] ;
    output \encoder1_position[7] ;
    output \encoder1_position[6] ;
    output \encoder1_position[5] ;
    output \encoder1_position[4] ;
    output \encoder1_position[3] ;
    output \encoder1_position[2] ;
    output n1822;
    input VCC_net;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire position_31__N_3830, debounce_cnt, a_prev, direction_N_3832;
    wire [1:0]a_new_c;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire a_prev_N_3835, n29752;
    wire [31:0]n133;
    
    wire n50526, n50525, n50524, n50523, n50522, n50521, n50520, 
        n50519, n50518, n50517, n50516, n50515, n50514, n50513, 
        n50512, n50511, n50510, n50509, n50508, n50507, n50506, 
        n50505, n50504, n50503, n50502, n50501, n50500, n50499, 
        n50498, n50497, n50496, n29477;
    
    SB_LUT4 b_prev_I_0_43_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(position_31__N_3830));   // vhdl/quadrature_decoder.vhd(63[37:56])
    defparam b_prev_I_0_43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(position_31__N_3830), 
            .I3(a_new[1]), .O(position_31__N_3827));   // vhdl/quadrature_decoder.vhd(62[7] 63[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 b_prev_I_0_45_2_lut (.I0(b_prev), .I1(a_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3832));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_45_2_lut.LUT_INIT = 16'h9999;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1779), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new_c[0]), .C(n1779), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 i52693_4_lut (.I0(a_new_c[0]), .I1(b_new[0]), .I2(a_new[1]), 
            .I3(b_new[1]), .O(a_prev_N_3835));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i52693_4_lut.LUT_INIT = 16'h8421;
    SB_DFF debounce_cnt_37 (.Q(debounce_cnt), .C(n1779), .D(a_prev_N_3835));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_prev_38 (.Q(a_prev), .C(n1779), .D(n29752));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_40 (.Q(n1784), .C(n1779), .D(n29704));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_1944__i0 (.Q(n1824), .C(n1779), .E(position_31__N_3827), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 position_1944_add_4_33_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1786), .I3(n50526), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_1944_add_4_32_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1788), .I3(n50525), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_32 (.CI(n50525), .I0(direction_N_3832), 
            .I1(n1788), .CO(n50526));
    SB_LUT4 position_1944_add_4_31_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1790), .I3(n50524), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_31 (.CI(n50524), .I0(direction_N_3832), 
            .I1(n1790), .CO(n50525));
    SB_LUT4 position_1944_add_4_30_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1792), .I3(n50523), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_30 (.CI(n50523), .I0(direction_N_3832), 
            .I1(n1792), .CO(n50524));
    SB_LUT4 position_1944_add_4_29_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1794), .I3(n50522), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_29 (.CI(n50522), .I0(direction_N_3832), 
            .I1(n1794), .CO(n50523));
    SB_LUT4 position_1944_add_4_28_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1796), .I3(n50521), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_28 (.CI(n50521), .I0(direction_N_3832), 
            .I1(n1796), .CO(n50522));
    SB_LUT4 position_1944_add_4_27_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[25] ), .I3(n50520), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_27 (.CI(n50520), .I0(direction_N_3832), 
            .I1(\encoder1_position[25] ), .CO(n50521));
    SB_LUT4 position_1944_add_4_26_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[24] ), .I3(n50519), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_26 (.CI(n50519), .I0(direction_N_3832), 
            .I1(\encoder1_position[24] ), .CO(n50520));
    SB_LUT4 position_1944_add_4_25_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[23] ), .I3(n50518), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_25 (.CI(n50518), .I0(direction_N_3832), 
            .I1(\encoder1_position[23] ), .CO(n50519));
    SB_LUT4 position_1944_add_4_24_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[22] ), .I3(n50517), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_24 (.CI(n50517), .I0(direction_N_3832), 
            .I1(\encoder1_position[22] ), .CO(n50518));
    SB_LUT4 position_1944_add_4_23_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[21] ), .I3(n50516), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_23 (.CI(n50516), .I0(direction_N_3832), 
            .I1(\encoder1_position[21] ), .CO(n50517));
    SB_LUT4 position_1944_add_4_22_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[20] ), .I3(n50515), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_22 (.CI(n50515), .I0(direction_N_3832), 
            .I1(\encoder1_position[20] ), .CO(n50516));
    SB_LUT4 position_1944_add_4_21_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[19] ), .I3(n50514), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_21 (.CI(n50514), .I0(direction_N_3832), 
            .I1(\encoder1_position[19] ), .CO(n50515));
    SB_LUT4 position_1944_add_4_20_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[18] ), .I3(n50513), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_20 (.CI(n50513), .I0(direction_N_3832), 
            .I1(\encoder1_position[18] ), .CO(n50514));
    SB_LUT4 position_1944_add_4_19_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[17] ), .I3(n50512), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_19 (.CI(n50512), .I0(direction_N_3832), 
            .I1(\encoder1_position[17] ), .CO(n50513));
    SB_LUT4 position_1944_add_4_18_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[16] ), .I3(n50511), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_DFFE position_1944__i31 (.Q(n1786), .C(n1779), .E(position_31__N_3827), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_CARRY position_1944_add_4_18 (.CI(n50511), .I0(direction_N_3832), 
            .I1(\encoder1_position[16] ), .CO(n50512));
    SB_LUT4 position_1944_add_4_17_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[15] ), .I3(n50510), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_17 (.CI(n50510), .I0(direction_N_3832), 
            .I1(\encoder1_position[15] ), .CO(n50511));
    SB_LUT4 position_1944_add_4_16_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[14] ), .I3(n50509), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_16 (.CI(n50509), .I0(direction_N_3832), 
            .I1(\encoder1_position[14] ), .CO(n50510));
    SB_LUT4 position_1944_add_4_15_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[13] ), .I3(n50508), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_15 (.CI(n50508), .I0(direction_N_3832), 
            .I1(\encoder1_position[13] ), .CO(n50509));
    SB_LUT4 position_1944_add_4_14_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[12] ), .I3(n50507), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_14 (.CI(n50507), .I0(direction_N_3832), 
            .I1(\encoder1_position[12] ), .CO(n50508));
    SB_LUT4 position_1944_add_4_13_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[11] ), .I3(n50506), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_DFFE position_1944__i30 (.Q(n1788), .C(n1779), .E(position_31__N_3827), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i29 (.Q(n1790), .C(n1779), .E(position_31__N_3827), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i28 (.Q(n1792), .C(n1779), .E(position_31__N_3827), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i27 (.Q(n1794), .C(n1779), .E(position_31__N_3827), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i26 (.Q(n1796), .C(n1779), .E(position_31__N_3827), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i25 (.Q(\encoder1_position[25] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i24 (.Q(\encoder1_position[24] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i23 (.Q(\encoder1_position[23] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i22 (.Q(\encoder1_position[22] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i21 (.Q(\encoder1_position[21] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i20 (.Q(\encoder1_position[20] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i19 (.Q(\encoder1_position[19] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i18 (.Q(\encoder1_position[18] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_CARRY position_1944_add_4_13 (.CI(n50506), .I0(direction_N_3832), 
            .I1(\encoder1_position[11] ), .CO(n50507));
    SB_DFFE position_1944__i17 (.Q(\encoder1_position[17] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i16 (.Q(\encoder1_position[16] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i15 (.Q(\encoder1_position[15] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i14 (.Q(\encoder1_position[14] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i13 (.Q(\encoder1_position[13] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i12 (.Q(\encoder1_position[12] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i11 (.Q(\encoder1_position[11] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i10 (.Q(\encoder1_position[10] ), .C(n1779), 
            .E(position_31__N_3827), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i9 (.Q(\encoder1_position[9] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i8 (.Q(\encoder1_position[8] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i7 (.Q(\encoder1_position[7] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i6 (.Q(\encoder1_position[6] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i5 (.Q(\encoder1_position[5] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i4 (.Q(\encoder1_position[4] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i3 (.Q(\encoder1_position[3] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i2 (.Q(\encoder1_position[2] ), .C(n1779), .E(position_31__N_3827), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_1944__i1 (.Q(n1822), .C(n1779), .E(position_31__N_3827), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 position_1944_add_4_12_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[10] ), .I3(n50505), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_12 (.CI(n50505), .I0(direction_N_3832), 
            .I1(\encoder1_position[10] ), .CO(n50506));
    SB_LUT4 position_1944_add_4_11_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[9] ), .I3(n50504), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_11 (.CI(n50504), .I0(direction_N_3832), 
            .I1(\encoder1_position[9] ), .CO(n50505));
    SB_LUT4 position_1944_add_4_10_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[8] ), .I3(n50503), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_10 (.CI(n50503), .I0(direction_N_3832), 
            .I1(\encoder1_position[8] ), .CO(n50504));
    SB_LUT4 position_1944_add_4_9_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[7] ), .I3(n50502), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_9 (.CI(n50502), .I0(direction_N_3832), 
            .I1(\encoder1_position[7] ), .CO(n50503));
    SB_LUT4 position_1944_add_4_8_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[6] ), .I3(n50501), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_8 (.CI(n50501), .I0(direction_N_3832), 
            .I1(\encoder1_position[6] ), .CO(n50502));
    SB_LUT4 position_1944_add_4_7_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[5] ), .I3(n50500), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_7 (.CI(n50500), .I0(direction_N_3832), 
            .I1(\encoder1_position[5] ), .CO(n50501));
    SB_LUT4 position_1944_add_4_6_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[4] ), .I3(n50499), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_6 (.CI(n50499), .I0(direction_N_3832), 
            .I1(\encoder1_position[4] ), .CO(n50500));
    SB_LUT4 position_1944_add_4_5_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[3] ), .I3(n50498), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_5 (.CI(n50498), .I0(direction_N_3832), 
            .I1(\encoder1_position[3] ), .CO(n50499));
    SB_LUT4 position_1944_add_4_4_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(\encoder1_position[2] ), .I3(n50497), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_4 (.CI(n50497), .I0(direction_N_3832), 
            .I1(\encoder1_position[2] ), .CO(n50498));
    SB_LUT4 position_1944_add_4_3_lut (.I0(GND_net), .I1(direction_N_3832), 
            .I2(n1822), .I3(n50496), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_3 (.CI(n50496), .I0(direction_N_3832), 
            .I1(n1822), .CO(n50497));
    SB_LUT4 position_1944_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1824), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1944_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1944_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(n1824), 
            .CO(n50496));
    SB_DFF b_prev_39 (.Q(b_prev), .C(n1779), .D(n29477));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i1 (.Q(a_new[1]), .C(n1779), .D(a_new_c[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1779), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 i15744_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3835), .I2(a_new[1]), 
            .I3(a_prev), .O(n29752));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15744_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15469_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3835), .I2(b_new[1]), 
            .I3(b_prev), .O(n29477));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i15469_3_lut_4_lut.LUT_INIT = 16'hf780;
    
endmodule
//
// Verilog Description of module coms
//

module coms (n29968, \data_in_frame[22] , clk16MHz, VCC_net, \data_in_frame[4] , 
            \FRAME_MATCHER.i_31__N_2509 , \data_out_frame[23] , neopxl_color, 
            \data_out_frame[25] , GND_net, \FRAME_MATCHER.state[3] , \data_out_frame[22] , 
            \current[7] , n51598, n3470, \current[6] , \current[5] , 
            n2873, \data_out_frame[8] , n56908, \current[4] , n56907, 
            \current[3] , \current[2] , \data_out_frame[18] , \current[1] , 
            \current[0] , \data_out_frame[21] , \current[15] , n52657, 
            \current[11] , n57377, n57350, \data_out_frame[20] , \current[10] , 
            \data_out_frame[24] , \current[9] , \current[8] , displacement, 
            n59466, n57295, \data_out_frame[19] , n51730, n51640, 
            \data_out_frame[15] , n51676, \data_out_frame[13] , n57232, 
            \data_out_frame[16] , n52803, n59193, n57398, \data_out_frame[17] , 
            n68335, \data_out_frame[14] , n68339, \data_out_frame[11] , 
            \data_out_frame[12] , \data_out_frame[6] , n29959, n51654, 
            n29956, n29953, n29663, n29949, n29946, n57741, \data_in_frame[3][6] , 
            \data_in_frame[3][5] , n25810, n65441, n65487, \data_in_frame[3][4] , 
            n29669, \data_in_frame[3][3] , \data_in_frame[3][2] , \data_in_frame[3][1] , 
            n57456, \data_in_frame[3][0] , \data_in_frame[2] , n29674, 
            n57131, n22726, \data_in_frame[11] , \data_in_frame[17] , 
            \data_in_frame[8] , \data_in_frame[9] , \data_out_frame[10] , 
            \data_in_frame[10] , \data_in_frame[1] , setpoint, \data_in_frame[6][5] , 
            \data_out_frame[5] , \data_out_frame[7] , n56906, n56905, 
            \data_out_frame[9] , n26524, \data_out_frame[4] , n56952, 
            \data_in_frame[6][4] , Kp_23__N_1748, reset, n59636, \data_in_frame[20] , 
            n56031, \data_in_frame[18] , \data_in_frame[21] , rx_data_ready, 
            rx_data, n57516, n56904, n56773, n56903, pwm_setpoint, 
            \data_in_frame[16] , n56902, n56901, n56900, n56899, n56898, 
            n56897, n56896, n56895, n56894, n56893, n56892, n56891, 
            n56890, n56889, n56888, n56887, n56886, n56885, n56884, 
            n56883, n56882, n56881, n56880, n56879, n56878, n56877, 
            n56876, n56875, n56874, n56873, n30569, n29046, n56872, 
            \data_in_frame[12] , n26482, n56871, n56870, \data_in_frame[13] , 
            \FRAME_MATCHER.rx_data_ready_prev , n57917, \data_in_frame[19] , 
            n56869, n56868, n56867, n28417, n29684, n8, n161, 
            n10, n10_adj_11, encoder0_position_scaled, \data_out_frame[26][2] , 
            \byte_transmit_counter[2] , n29889, n29687, \byte_transmit_counter[1] , 
            encoder1_position_scaled, n29885, n29881, n29878, n56866, 
            n56865, n56864, \data_in_frame[15][6] , \data_out_frame[27][2] , 
            n56027, n56863, n29874, n56862, n56861, n56860, n59242, 
            n56859, n56858, n30585, n29030, n56857, n56856, n56855, 
            n29870, n29867, n28387, \FRAME_MATCHER.i[5] , \FRAME_MATCHER.i[3] , 
            \byte_transmit_counter[0] , n376, n456, n11610, n27692, 
            n29853, deadband, n29849, n29848, n29847, n29846, n29845, 
            n29844, n29843, n29842, n29841, n29840, n29839, n29837, 
            n29836, n29835, n29834, n29833, n29832, n29831, n29830, 
            n29829, n29828, n29827, IntegralLimit, n29826, n29825, 
            n29824, n29823, n29822, n29821, n29820, n29819, n29818, 
            n29817, n29816, n29815, n29814, n29813, n29812, n29811, 
            n29810, n29809, n29808, n29807, n29806, n29805, n29804, 
            \Kp[1] , n29803, \Kp[2] , n29802, \Kp[3] , \pwm_counter[22] , 
            n45, \pwm_counter[21] , n43, n29801, \Kp[4] , n29800, 
            \Kp[5] , n29799, \Kp[6] , \Kp[7] , n29797, \Kp[8] , 
            n29796, \Kp[9] , n29795, \Kp[10] , n29794, \Kp[11] , 
            n29793, \Kp[12] , n29792, \Kp[13] , n29791, \Kp[14] , 
            n29790, \Kp[15] , n29789, \Ki[1] , n29788, \Ki[2] , 
            n29787, \Ki[3] , n29786, \Ki[4] , n29785, \Ki[5] , n29784, 
            \Ki[6] , n29783, \Ki[7] , n29782, \Ki[8] , n29781, \Ki[9] , 
            n29780, \Ki[10] , n29779, \Ki[11] , n29778, \Ki[12] , 
            n29777, \Ki[13] , \Ki[14] , n29775, \Ki[15] , n56854, 
            n56853, n56852, n56851, n56850, n56849, n56775, n56777, 
            n57044, n56778, n56779, n56780, n56781, n56783, n56784, 
            n56785, n56786, n56787, n56788, n29746, n56789, n56790, 
            n56791, n56792, n29736, n56793, n56774, n56794, n56795, 
            n56796, n29735, current_limit, n29734, control_mode, n29733, 
            n29732, n29731, n56797, n56798, n29727, n29726, n29725, 
            n29723, n29722, n29721, n29720, n29719, n29718, n29717, 
            n56799, n56800, n29716, n29712, n29711, n56801, n56802, 
            n29708, n29707, n56803, n29706, n29705, n29703, n29702, 
            n29698, n29694, n40973, n28438, n29691, Kp_23__N_1301, 
            n57039, \data_in_frame[15][7] , \data_in_frame[15][4] , n57780, 
            n29673, n29672, n29662, n29644, PWMLimit, n29639, n29638, 
            n29637, n29636, \Ki[0] , n29635, \Kp[0] , n29613, n56804, 
            n56805, n56806, n30647, n28989, n56807, n30649, n28987, 
            n56808, n56809, n56810, n56811, n56812, n30655, n28981, 
            n56813, n56814, n56815, n56816, n56817, n56818, n56819, 
            n56820, n56821, n56822, n56823, n56824, n56825, n8_adj_12, 
            n56826, n56827, n56828, n56829, n56830, n56831, \data_out_frame[0][2] , 
            n56951, \data_out_frame[0][3] , n56950, \data_out_frame[0][4] , 
            n56949, \data_out_frame[1][0] , n56948, \data_in_frame[16][7] , 
            \data_in_frame[19][3] , n57717, \data_out_frame[1][1] , n56947, 
            \data_out_frame[1][3] , n56946, \data_out_frame[1][5] , n56945, 
            \data_in_frame[15][1] , \data_in_frame[14] , n25864, n57720, 
            \data_out_frame[1][6] , n56944, \data_in_frame[19][4] , \data_out_frame[1][7] , 
            n56943, \data_out_frame[3][1] , n56942, \data_in_frame[15][3] , 
            n30519, n30518, n30517, n30515, n30514, n30513, n30512, 
            \data_in_frame[15][0] , \data_in_frame[15][2] , n30470, n30468, 
            n30467, n30466, n30465, n30464, n30444, n30398, n30396, 
            n30395, n30384, n30375, \data_out_frame[3][3] , n56941, 
            n25952, \data_out_frame[3][4] , n56940, n30350, n30349, 
            n30348, n30347, n29973, \data_in_frame[5] , n29976, n30343, 
            n29979, n29982, n56201, \data_in_frame[16][1] , n30339, 
            n56199, \data_in_frame[16][2] , n29490, n29493, n29496, 
            n29499, n56249, n56107, n56103, n56101, n56099, n56095, 
            n56091, \data_out_frame[3][6] , n56771, n29986, n29989, 
            n29992, n56087, n56083, n56079, n30305, n29995, \data_in_frame[6][0] , 
            \data_in_frame[6][1] , \data_in_frame[6][2] , \data_in_frame[6][3] , 
            n30299, \data_out_frame[3][7] , n56939, n30047, n30050, 
            n30054, n30057, n30282, n30281, n30280, n30063, n30066, 
            n30069, n30072, n30075, n30079, n30082, n30085, n30089, 
            n30092, n30095, \data_in_frame[10][1] , \data_in_frame[10][2] , 
            \data_in_frame[10][3] , \data_in_frame[10][5] , \data_in_frame[10][7] , 
            n30149, n30152, n30250, n30156, n56303, n56343, n30166, 
            n30169, n30172, n30176, n30179, n30182, n30186, n30189, 
            n30192, n30196, n56075, n56071, n30232, n29540, n29543, 
            n29546, n56065, n56061, n56057, \data_in_frame[19][0] , 
            n56053, \data_in_frame[19][1] , n56049, \data_in_frame[19][2] , 
            n30207, n56045, n56041, \data_in_frame[19][5] , n56037, 
            n29579, n29588, n29591, n29594, n30155, n57701, n29600, 
            n57361, n57467, n56938, n172, n33761, n30739, n29117, 
            n30740, n29116, n30741, n29115, n56937, n59574, n29509, 
            n10_adj_13, n56936, n56935, n57473, \FRAME_MATCHER.i_31__N_2513 , 
            n56934, n56933, n56932, n56931, n56930, n56929, n56928, 
            n56927, n56926, n56925, n56924, n56923, n56922, n56921, 
            n56920, n56919, n29480, n57125, n57680, n29478, n56832, 
            n56833, n56834, n56835, n56836, n56837, n56838, n56839, 
            n56840, n56772, n56782, n56841, n56842, n56843, n56844, 
            n56918, n56917, n56916, n56915, n56845, n56846, n56847, 
            n56848, n56776, LED_c, n56914, DE_c, n56913, n56912, 
            n56911, n56910, n29969, n56909, n92, ID, n33769, n27696, 
            n28383, n28379, n28434, n26, n21, tx_active, n57921, 
            n260, n8_adj_14, n130, n65436, n28428, n59230, n375, 
            n455, n37189, n15, n15_adj_15, n19, n28375, n56988, 
            n8_adj_16, n28381, n69525, n4, n4_adj_17, n30, n361, 
            n32, n69309, n25, n134, n20, n43_adj_18, n401, n4_adj_19, 
            n65432, n69489, n62711, n62712, n62859, n62858, n52677, 
            r_SM_Main, n57935, n6, tx_o, n29661, r_Clock_Count, 
            n4940, n27, tx_enable, \r_Bit_Index[0] , n4937, \o_Rx_DV_N_3488[8] , 
            n60724, baudrate, \r_SM_Main[2]_adj_20 , n25530, r_Rx_Data, 
            RX_N_2, \r_SM_Main[1]_adj_21 , n27966, n56959, n60740, 
            n29884, n60788, n60756, n29866, \o_Rx_DV_N_3488[7] , \o_Rx_DV_N_3488[6] , 
            \o_Rx_DV_N_3488[5] , \o_Rx_DV_N_3488[4] , \o_Rx_DV_N_3488[3] , 
            \o_Rx_DV_N_3488[2] , \o_Rx_DV_N_3488[1] , \o_Rx_DV_N_3488[0] , 
            n29774, n29773, n29772, r_Clock_Count_adj_30, n58000, 
            n30502, n52851, n30498, n30201, n30200, n60708, n60692, 
            n60804, n27724, n60772) /* synthesis syn_module_defined=1 */ ;
    input n29968;
    output [7:0]\data_in_frame[22] ;
    input clk16MHz;
    input VCC_net;
    output [7:0]\data_in_frame[4] ;
    output \FRAME_MATCHER.i_31__N_2509 ;
    output [7:0]\data_out_frame[23] ;
    output [23:0]neopxl_color;
    output [7:0]\data_out_frame[25] ;
    input GND_net;
    output \FRAME_MATCHER.state[3] ;
    output [7:0]\data_out_frame[22] ;
    input \current[7] ;
    input n51598;
    output n3470;
    input \current[6] ;
    input \current[5] ;
    input n2873;
    output [7:0]\data_out_frame[8] ;
    input n56908;
    input \current[4] ;
    input n56907;
    input \current[3] ;
    input \current[2] ;
    output [7:0]\data_out_frame[18] ;
    input \current[1] ;
    input \current[0] ;
    output [7:0]\data_out_frame[21] ;
    input \current[15] ;
    input n52657;
    input \current[11] ;
    output n57377;
    input n57350;
    output [7:0]\data_out_frame[20] ;
    input \current[10] ;
    output [7:0]\data_out_frame[24] ;
    input \current[9] ;
    input \current[8] ;
    input [23:0]displacement;
    output n59466;
    output n57295;
    output [7:0]\data_out_frame[19] ;
    output n51730;
    output n51640;
    output [7:0]\data_out_frame[15] ;
    output n51676;
    output [7:0]\data_out_frame[13] ;
    output n57232;
    output [7:0]\data_out_frame[16] ;
    output n52803;
    output n59193;
    output n57398;
    output [7:0]\data_out_frame[17] ;
    output n68335;
    output [7:0]\data_out_frame[14] ;
    output n68339;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[6] ;
    input n29959;
    output n51654;
    input n29956;
    input n29953;
    input n29663;
    input n29949;
    input n29946;
    input n57741;
    output \data_in_frame[3][6] ;
    output \data_in_frame[3][5] ;
    input n25810;
    input n65441;
    input n65487;
    output \data_in_frame[3][4] ;
    input n29669;
    output \data_in_frame[3][3] ;
    output \data_in_frame[3][2] ;
    output \data_in_frame[3][1] ;
    output n57456;
    output \data_in_frame[3][0] ;
    output [7:0]\data_in_frame[2] ;
    input n29674;
    output n57131;
    input n22726;
    output [7:0]\data_in_frame[11] ;
    output [7:0]\data_in_frame[17] ;
    output [7:0]\data_in_frame[8] ;
    output [7:0]\data_in_frame[9] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_in_frame[10] ;
    output [7:0]\data_in_frame[1] ;
    output [23:0]setpoint;
    output \data_in_frame[6][5] ;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[7] ;
    input n56906;
    input n56905;
    output [7:0]\data_out_frame[9] ;
    input n26524;
    output [7:0]\data_out_frame[4] ;
    input n56952;
    output \data_in_frame[6][4] ;
    output Kp_23__N_1748;
    input reset;
    input n59636;
    output [7:0]\data_in_frame[20] ;
    input n56031;
    output [7:0]\data_in_frame[18] ;
    output [7:0]\data_in_frame[21] ;
    output rx_data_ready;
    output [7:0]rx_data;
    input n57516;
    input n56904;
    input n56773;
    input n56903;
    input [23:0]pwm_setpoint;
    output [7:0]\data_in_frame[16] ;
    input n56902;
    input n56901;
    input n56900;
    input n56899;
    input n56898;
    input n56897;
    input n56896;
    input n56895;
    input n56894;
    input n56893;
    input n56892;
    input n56891;
    input n56890;
    input n56889;
    input n56888;
    input n56887;
    input n56886;
    input n56885;
    input n56884;
    input n56883;
    input n56882;
    input n56881;
    input n56880;
    input n56879;
    input n56878;
    input n56877;
    input n56876;
    input n56875;
    input n56874;
    input n56873;
    input n30569;
    input n29046;
    input n56872;
    output [7:0]\data_in_frame[12] ;
    output n26482;
    input n56871;
    input n56870;
    output [7:0]\data_in_frame[13] ;
    output \FRAME_MATCHER.rx_data_ready_prev ;
    output n57917;
    output [7:0]\data_in_frame[19] ;
    input n56869;
    input n56868;
    input n56867;
    input n28417;
    input n29684;
    output n8;
    output n161;
    output n10;
    output n10_adj_11;
    input [23:0]encoder0_position_scaled;
    output \data_out_frame[26][2] ;
    output \byte_transmit_counter[2] ;
    input n29889;
    input n29687;
    output \byte_transmit_counter[1] ;
    input [23:0]encoder1_position_scaled;
    input n29885;
    input n29881;
    input n29878;
    input n56866;
    input n56865;
    input n56864;
    output \data_in_frame[15][6] ;
    output \data_out_frame[27][2] ;
    input n56027;
    input n56863;
    input n29874;
    input n56862;
    input n56861;
    input n56860;
    output n59242;
    input n56859;
    input n56858;
    input n30585;
    input n29030;
    input n56857;
    input n56856;
    input n56855;
    input n29870;
    input n29867;
    output n28387;
    output \FRAME_MATCHER.i[5] ;
    output \FRAME_MATCHER.i[3] ;
    output \byte_transmit_counter[0] ;
    input n376;
    input n456;
    input n11610;
    output n27692;
    input n29853;
    output [23:0]deadband;
    input n29849;
    input n29848;
    input n29847;
    input n29846;
    input n29845;
    input n29844;
    input n29843;
    input n29842;
    input n29841;
    input n29840;
    input n29839;
    input n29837;
    input n29836;
    input n29835;
    input n29834;
    input n29833;
    input n29832;
    input n29831;
    input n29830;
    input n29829;
    input n29828;
    input n29827;
    output [23:0]IntegralLimit;
    input n29826;
    input n29825;
    input n29824;
    input n29823;
    input n29822;
    input n29821;
    input n29820;
    input n29819;
    input n29818;
    input n29817;
    input n29816;
    input n29815;
    input n29814;
    input n29813;
    input n29812;
    input n29811;
    input n29810;
    input n29809;
    input n29808;
    input n29807;
    input n29806;
    input n29805;
    input n29804;
    output \Kp[1] ;
    input n29803;
    output \Kp[2] ;
    input n29802;
    output \Kp[3] ;
    input \pwm_counter[22] ;
    output n45;
    input \pwm_counter[21] ;
    output n43;
    input n29801;
    output \Kp[4] ;
    input n29800;
    output \Kp[5] ;
    input n29799;
    output \Kp[6] ;
    output \Kp[7] ;
    input n29797;
    output \Kp[8] ;
    input n29796;
    output \Kp[9] ;
    input n29795;
    output \Kp[10] ;
    input n29794;
    output \Kp[11] ;
    input n29793;
    output \Kp[12] ;
    input n29792;
    output \Kp[13] ;
    input n29791;
    output \Kp[14] ;
    input n29790;
    output \Kp[15] ;
    input n29789;
    output \Ki[1] ;
    input n29788;
    output \Ki[2] ;
    input n29787;
    output \Ki[3] ;
    input n29786;
    output \Ki[4] ;
    input n29785;
    output \Ki[5] ;
    input n29784;
    output \Ki[6] ;
    input n29783;
    output \Ki[7] ;
    input n29782;
    output \Ki[8] ;
    input n29781;
    output \Ki[9] ;
    input n29780;
    output \Ki[10] ;
    input n29779;
    output \Ki[11] ;
    input n29778;
    output \Ki[12] ;
    input n29777;
    output \Ki[13] ;
    output \Ki[14] ;
    input n29775;
    output \Ki[15] ;
    input n56854;
    input n56853;
    input n56852;
    input n56851;
    input n56850;
    input n56849;
    input n56775;
    input n56777;
    output n57044;
    input n56778;
    input n56779;
    input n56780;
    input n56781;
    input n56783;
    input n56784;
    input n56785;
    input n56786;
    input n56787;
    input n56788;
    input n29746;
    input n56789;
    input n56790;
    input n56791;
    input n56792;
    input n29736;
    input n56793;
    input n56774;
    input n56794;
    input n56795;
    input n56796;
    input n29735;
    output [15:0]current_limit;
    input n29734;
    output [7:0]control_mode;
    input n29733;
    input n29732;
    input n29731;
    input n56797;
    input n56798;
    input n29727;
    input n29726;
    input n29725;
    input n29723;
    input n29722;
    input n29721;
    input n29720;
    input n29719;
    input n29718;
    input n29717;
    input n56799;
    input n56800;
    input n29716;
    input n29712;
    input n29711;
    input n56801;
    input n56802;
    input n29708;
    input n29707;
    input n56803;
    input n29706;
    input n29705;
    input n29703;
    input n29702;
    input n29698;
    input n29694;
    output n40973;
    output n28438;
    input n29691;
    input Kp_23__N_1301;
    output n57039;
    output \data_in_frame[15][7] ;
    output \data_in_frame[15][4] ;
    input n57780;
    input n29673;
    input n29672;
    input n29662;
    input n29644;
    output [23:0]PWMLimit;
    input n29639;
    input n29638;
    input n29637;
    input n29636;
    output \Ki[0] ;
    input n29635;
    output \Kp[0] ;
    input n29613;
    input n56804;
    input n56805;
    input n56806;
    input n30647;
    input n28989;
    input n56807;
    input n30649;
    input n28987;
    input n56808;
    input n56809;
    input n56810;
    input n56811;
    input n56812;
    input n30655;
    input n28981;
    input n56813;
    input n56814;
    input n56815;
    input n56816;
    input n56817;
    input n56818;
    input n56819;
    input n56820;
    input n56821;
    input n56822;
    input n56823;
    input n56824;
    input n56825;
    output n8_adj_12;
    input n56826;
    input n56827;
    input n56828;
    input n56829;
    input n56830;
    input n56831;
    output \data_out_frame[0][2] ;
    input n56951;
    output \data_out_frame[0][3] ;
    input n56950;
    output \data_out_frame[0][4] ;
    input n56949;
    output \data_out_frame[1][0] ;
    input n56948;
    output \data_in_frame[16][7] ;
    output \data_in_frame[19][3] ;
    input n57717;
    output \data_out_frame[1][1] ;
    input n56947;
    output \data_out_frame[1][3] ;
    input n56946;
    output \data_out_frame[1][5] ;
    input n56945;
    output \data_in_frame[15][1] ;
    output [7:0]\data_in_frame[14] ;
    output n25864;
    output n57720;
    output \data_out_frame[1][6] ;
    input n56944;
    output \data_in_frame[19][4] ;
    output \data_out_frame[1][7] ;
    input n56943;
    output \data_out_frame[3][1] ;
    input n56942;
    output \data_in_frame[15][3] ;
    input n30519;
    input n30518;
    input n30517;
    input n30515;
    input n30514;
    input n30513;
    input n30512;
    output \data_in_frame[15][0] ;
    output \data_in_frame[15][2] ;
    input n30470;
    input n30468;
    input n30467;
    input n30466;
    input n30465;
    input n30464;
    input n30444;
    input n30398;
    input n30396;
    input n30395;
    input n30384;
    input n30375;
    output \data_out_frame[3][3] ;
    input n56941;
    output n25952;
    output \data_out_frame[3][4] ;
    input n56940;
    input n30350;
    input n30349;
    input n30348;
    input n30347;
    input n29973;
    output [7:0]\data_in_frame[5] ;
    input n29976;
    input n30343;
    input n29979;
    input n29982;
    input n56201;
    output \data_in_frame[16][1] ;
    input n30339;
    input n56199;
    output \data_in_frame[16][2] ;
    input n29490;
    input n29493;
    input n29496;
    input n29499;
    input n56249;
    input n56107;
    input n56103;
    input n56101;
    input n56099;
    input n56095;
    input n56091;
    output \data_out_frame[3][6] ;
    input n56771;
    input n29986;
    input n29989;
    input n29992;
    input n56087;
    input n56083;
    input n56079;
    input n30305;
    input n29995;
    output \data_in_frame[6][0] ;
    output \data_in_frame[6][1] ;
    output \data_in_frame[6][2] ;
    output \data_in_frame[6][3] ;
    input n30299;
    output \data_out_frame[3][7] ;
    input n56939;
    input n30047;
    input n30050;
    input n30054;
    input n30057;
    input n30282;
    input n30281;
    input n30280;
    input n30063;
    input n30066;
    input n30069;
    input n30072;
    input n30075;
    input n30079;
    input n30082;
    input n30085;
    input n30089;
    input n30092;
    input n30095;
    output \data_in_frame[10][1] ;
    output \data_in_frame[10][2] ;
    output \data_in_frame[10][3] ;
    output \data_in_frame[10][5] ;
    output \data_in_frame[10][7] ;
    input n30149;
    input n30152;
    input n30250;
    input n30156;
    input n56303;
    input n56343;
    input n30166;
    input n30169;
    input n30172;
    input n30176;
    input n30179;
    input n30182;
    input n30186;
    input n30189;
    input n30192;
    input n30196;
    input n56075;
    input n56071;
    input n30232;
    input n29540;
    input n29543;
    input n29546;
    input n56065;
    input n56061;
    input n56057;
    output \data_in_frame[19][0] ;
    input n56053;
    output \data_in_frame[19][1] ;
    input n56049;
    output \data_in_frame[19][2] ;
    input n30207;
    input n56045;
    input n56041;
    output \data_in_frame[19][5] ;
    input n56037;
    input n29579;
    input n29588;
    input n29591;
    input n29594;
    input n30155;
    output n57701;
    input n29600;
    input n57361;
    output n57467;
    input n56938;
    output n172;
    output n33761;
    input n30739;
    input n29117;
    input n30740;
    input n29116;
    input n30741;
    input n29115;
    input n56937;
    input n59574;
    input n29509;
    input n10_adj_13;
    input n56936;
    input n56935;
    output n57473;
    output \FRAME_MATCHER.i_31__N_2513 ;
    input n56934;
    input n56933;
    input n56932;
    input n56931;
    input n56930;
    input n56929;
    input n56928;
    input n56927;
    input n56926;
    input n56925;
    input n56924;
    input n56923;
    input n56922;
    input n56921;
    input n56920;
    input n56919;
    input n29480;
    output n57125;
    output n57680;
    input n29478;
    input n56832;
    input n56833;
    input n56834;
    input n56835;
    input n56836;
    input n56837;
    input n56838;
    input n56839;
    input n56840;
    input n56772;
    input n56782;
    input n56841;
    input n56842;
    input n56843;
    input n56844;
    input n56918;
    input n56917;
    input n56916;
    input n56915;
    input n56845;
    input n56846;
    input n56847;
    input n56848;
    input n56776;
    output LED_c;
    input n56914;
    output DE_c;
    input n56913;
    input n56912;
    input n56911;
    input n56910;
    input n29969;
    input n56909;
    input n92;
    input [7:0]ID;
    output n33769;
    output n27696;
    output n28383;
    output n28379;
    input n28434;
    input n26;
    output n21;
    output tx_active;
    output n57921;
    output n260;
    output n8_adj_14;
    output n130;
    output n65436;
    output n28428;
    output n59230;
    input n375;
    input n455;
    output n37189;
    input n15;
    input n15_adj_15;
    output n19;
    output n28375;
    output n56988;
    output n8_adj_16;
    output n28381;
    output n69525;
    output n4;
    output n4_adj_17;
    input n30;
    input n361;
    output n32;
    input n69309;
    input n25;
    output n134;
    output n20;
    input n43_adj_18;
    input n401;
    output n4_adj_19;
    output n65432;
    output n69489;
    input n62711;
    input n62712;
    input n62859;
    input n62858;
    output n52677;
    output [2:0]r_SM_Main;
    input n57935;
    output n6;
    output tx_o;
    input n29661;
    output [8:0]r_Clock_Count;
    input n4940;
    output n27;
    output tx_enable;
    output \r_Bit_Index[0] ;
    input n4937;
    output \o_Rx_DV_N_3488[8] ;
    output n60724;
    input [31:0]baudrate;
    output \r_SM_Main[2]_adj_20 ;
    output n25530;
    output r_Rx_Data;
    input RX_N_2;
    output \r_SM_Main[1]_adj_21 ;
    output n27966;
    input n56959;
    output n60740;
    input n29884;
    output n60788;
    output n60756;
    input n29866;
    output \o_Rx_DV_N_3488[7] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[0] ;
    input n29774;
    input n29773;
    input n29772;
    output [7:0]r_Clock_Count_adj_30;
    output n58000;
    input n30502;
    input n52851;
    input n30498;
    input n30201;
    input n30200;
    output n60708;
    output n60692;
    output n60804;
    output n27724;
    output n60772;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n29967;
    wire [31:0]\FRAME_MATCHER.state_31__N_2612 ;
    
    wire n2, n51736, n57328, n57484, n57359, n3, n2_adj_4726, 
        n2_adj_4727, n2_adj_4728, n2_adj_4729, n2_adj_4730, n51658;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    wire [31:0]n133;
    
    wire \FRAME_MATCHER.i_31__N_2507 , n28050, n52789, n3_adj_4731, 
        n2_adj_4732, n29964, n2_adj_4733, n2_adj_4734, n2_adj_4735, 
        n2_adj_4736, n57245, n57392, n52665, n3_adj_4737, n57242, 
        n52576, n3_adj_4738, n2_adj_4739, n2_adj_4740, n57668, n2_adj_4741, 
        n2_adj_4742, n2_adj_4743, n2_adj_4744, n2_adj_4745, n2_adj_4746, 
        n51745, n14, n2_adj_4747, n9, n57626, n59922, n2_adj_4748, 
        n7, n52767, n2_adj_4749, n2_adj_4750, n2_adj_4751, n2_adj_4752, 
        n57609, n8_c, n2_adj_4753, n52735, n12, n2_adj_4754, n25071, 
        n3_adj_4755, n57325, n2_adj_4756, n3_adj_4757, n2_adj_4758, 
        n57065, n57412, n51784, n25716, n57659, n2_adj_4759, n57322, 
        n24, n2_adj_4760, n2_adj_4761, n51670, n57358, n52761, n22, 
        n2_adj_4762, n23668, n17, n59054, n26_c, n51672, n59736, 
        n57428, n24_adj_4763, n26_adj_4764, n57762, n25_c, n27_c, 
        n10_c, n14_adj_4765, n26374, n57283, n57395, n3_adj_4766, 
        n57633, n57487, n25158, n57216, n23709, n3_adj_4767, n57756, 
        n57647, n12_adj_4768, n57137, n8_adj_4769, n3_adj_4770, n51617, 
        n26825, n52130, n15_c, n51652, n14_adj_4771, n2217, n57641, 
        n57644, n10_adj_4772, n59521, n52581, n51837, n57419, n57422, 
        n10_adj_4773, n51832, n57460, n26693, n26394, n1699, n57450, 
        n23666, n6_c, n51605, n57305, n57416, n16, n771, \FRAME_MATCHER.i_31__N_2508 , 
        n1951, n1954, n25488, n25696, n57590, n51682, n26858, 
        n57689, n17_adj_4774, n60097, n4452, n1957, n59002, n26253, 
        n6_adj_4775, n57345, n25679, n1668, n51541, n26_adj_4776, 
        n57374, n57638, n24_adj_4777, n1191, n57692, n57596, n25_adj_4778, 
        n57729, n23, n58952, n52669, n18, n57587, n57200, n57553, 
        n24_adj_4779, n57570, n57185, n22_adj_4780, n57735, n25667, 
        n26_adj_4781, n57140, n62408, \FRAME_MATCHER.i_31__N_2514 , 
        n59835, n57386, n59591, n11, n56355;
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(99[12:25])
    
    wire n29666;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(99[12:25])
    
    wire n29939, n29936, n2076, n26241, n13, n52737, n51811, n16_adj_4782;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(105[12:33])
    
    wire n69177, n69480, n26626, n57413, n57235, n17_adj_4783, n69279, 
        n69315;
    wire [7:0]tx_data;   // verilog/coms.v(108[13:20])
    
    wire n57606, n69183, n65454, n69474, n69291, n7_adj_4784, n69189, 
        n65442, n69468, n69285, n7_adj_4785, n67511, n69462, n14_adj_4786, 
        n7_adj_4787, n29933, n29929, n29926, n59153, n10_adj_4788, 
        n10_adj_4789, n25095, n57446, n12_adj_4790, n52164, n29923, 
        n29920, n29917, n29913, n29910, n29678, n57560, n10_adj_4791, 
        n57747, n25734, n12_adj_4792, n6_adj_4793, n52327;
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(99[12:25])
    
    wire n29692, n29693, n51720, n10_adj_4794, n25128, n57404, n25853, 
        n59043, n57352, n6_adj_4795, Kp_23__N_1080, n57331, n25105, 
        n52618, n12_adj_4796, n8_adj_4797, n3_adj_4798, n57771, n26428, 
        n4_c, n57573, n26724, n62074, n57072, n57425, n12_adj_4799, 
        n2_adj_4800, n36, n57695, n26423, n26031, n2_adj_4801, n2_adj_4802, 
        n57732, n51619, n6_adj_4803, n26415, n25068, n26100, n25918, 
        n57280, n2_adj_4804, n2_adj_4805, n26257, n51753, n57171, 
        n25797, n57289, n26332, n26298, n57104, n57181, n2_adj_4806, 
        n57656, n57653, n57547, n59779, n1516, n26757, n57567, 
        n26363, n57108, n57111, n57622, n10_adj_4807, n57753, n57090, 
        n57759, Kp_23__N_872, n6_adj_4808, n25671, n57150, n2_adj_4809, 
        n6_adj_4810, n57154, n26066, n2_adj_4811, n10_adj_4812, n57265, 
        n1563, n14_adj_4813, n29906, n51805, n2_adj_4814, n26607, 
        n26335, n57157, n57160, n2_adj_4815, n57564, n57146, n6_adj_4816, 
        n51656, n57744, n14_adj_4817, n10_adj_4818, n57528, n57052, 
        n15_adj_4819, n14_adj_4820, n57248, n57613, n10_adj_4821, 
        n56737, n49184, n56736, n1720, n57203, n57178, n10_adj_4822, 
        n2_adj_4823, n57581, n26083, n10_adj_4824, Kp_23__N_878, n57271, 
        n57314, n57619, n26193, n57726, n2_adj_4825, n26662, n25893, 
        n35660, n57665, n2068, n29903;
    wire [23:0]n4762;
    
    wire n27737, n7_adj_4826, n57792, n57084, n2_adj_4827, n57441, 
        n8_adj_4828, n57789, n1130, n2_adj_4829, n28912, n4_adj_4830, 
        n62128;
    wire [7:0]\data_in[3] ;   // verilog/coms.v(98[12:19])
    
    wire n30351, n2_adj_4831, n56743, n49183, n22_adj_4832, n21_c, 
        n14_adj_4833, n23_adj_4834, n24_adj_4835, n2_adj_4836;
    wire [7:0]\data_in[1] ;   // verilog/coms.v(98[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(98[12:19])
    
    wire n29650, n2_adj_4837, n30382, n2_adj_4838, n29899, n18_adj_4839, 
        n30_c, n30381, n57342, n28, n32_c, n27_adj_4840, n8_adj_4841, 
        n7_adj_4842, n51588, n10_adj_4843, n59162, n2_adj_4844, n56742, 
        n49182, n57584, n2_adj_4845, n57175, n10_adj_4846, n30380, 
        n30379, n26780, n2_adj_4847, n29896, n2_adj_4848, n10_adj_4849, 
        n30378, n14_adj_4850, n2_adj_4851, n34, n30377, n24_adj_4852, 
        n38, n52624, n36_adj_4853, n30376, n2_adj_4854;
    wire [7:0]\data_in[2] ;   // verilog/coms.v(98[12:19])
    
    wire n30374, n22_adj_4855, n37, n2_adj_4856, n35, n12_adj_4857, 
        n59907, \FRAME_MATCHER.i_31__N_2511 , n33763, n6_adj_4858, n28901, 
        n57674, n57191, n30373, n2_adj_4859, n57786, n2_adj_4860, 
        n30372, n30371, n2_adj_4861, n2_adj_4862, n30370, n52017, 
        n52655, n51281, n57686, n52653, n8_adj_4863, n2_adj_4864, 
        n2_adj_4865, n2_adj_4866, n2_adj_4867, n2_adj_4868, n2_adj_4869, 
        n2_adj_4870, n2_adj_4871, n2_adj_4872, n2_adj_4873, n2_adj_4874, 
        n2_adj_4875, n2_adj_4876, n2_adj_4877, n2_adj_4878, n2_adj_4879, 
        n56741, n49181, n2_adj_4880, n30368, n30367, n30366, n6_adj_4881, 
        n57408, n30365, n30364, n25731, n6_adj_4882, n11_adj_4883, 
        n13_adj_4884, n28399, n56297, n30363, n6_adj_4885, n57317, 
        n2_adj_4886, n2_adj_4887, n2_adj_4888, n2_adj_4889, n2_adj_4890, 
        n2_adj_4891, n2_adj_4892, n2_adj_4893, n26272, n2_adj_4894, 
        n2_adj_4895, n2_adj_4896, n2_adj_4897, n2_adj_4898, n2_adj_4899, 
        n2_adj_4900, n2_adj_4901, n29893, n2_adj_4902, n30362, n6_adj_4903, 
        n14_adj_4904, n2_adj_4905, n2_adj_4906, n30361, n2_adj_4907, 
        n57068, n57534, n28415;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(99[12:25])
    
    wire n56157, n9_adj_4908, n68337, n2_adj_4909, n51646, n30360, 
        n30359, n30358, n2_adj_4910, n56163, n2_adj_4911, n56165, 
        n30357, n30356, n57671, n10_adj_4912, n3_adj_4913, n30355, 
        n2_adj_4914, n30354, n26449, n30353, n56740, n49180, n2_adj_4915, 
        n30352, n30369, n2_adj_4916, n2_adj_4917, n2_adj_4918;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    
    wire n56754, n2_adj_4919, n2_adj_4920, n59212, n59279, n51684, 
        n59284, n52615, n56369, n56755, n56367, n2_adj_4921, n28409, 
        n2_adj_4925, n56756, n62366, n2_adj_4926, Kp_23__N_748, n24_adj_4927, 
        n2_adj_4928, n26652, n2_adj_4929, n56752, n57519, n56739, 
        n49179, n56757, n56750, n56758, n56738, n49178, n56759;
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    
    wire n56760, n2_adj_4930, n28391;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(99[12:25])
    
    wire n56197, n2_adj_4931, n2_adj_4932, n56153, n2_adj_4933, n2_adj_4934, 
        n56761, n2_adj_4935, n56762, n56753, n56749, n2_adj_4936, 
        n2_adj_4937, n2_adj_4938, n2_adj_4939, n57041, n2_adj_4940, 
        n2_adj_4941, n2_adj_4942, n2_adj_4943, n56751, n2_adj_4944, 
        n2_adj_4945, n29699;
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(99[12:25])
    
    wire n56763, n56764, n40970, n7_adj_4946, n29713, n29728, n56744, 
        tx_transmit_N_3416, n29737, n29740, n56361, n29756, n29759, 
        n29762, n29765, n29768, n29850, n29838, n29798, n29776, 
        n43293, n145, n57016, n25991;
    wire [7:0]\data_in_frame[19]_c ;   // verilog/coms.v(99[12:25])
    
    wire n62126, n52651, n57463, n62134, n52695, n57497, n62140, 
        n57389, n57494, n62146, n2_adj_4947, n23898, n57371, n62152, 
        n57372, n57783, n57168, n57292, n25987, n57635, n57037, 
        n52594, n62014, n57433, n62018, n52337, n59955, n51926, 
        n57476, n62036;
    wire [7:0]\data_in_frame[16]_c ;   // verilog/coms.v(99[12:25])
    
    wire n62042, Kp_23__N_1389, n62046, n57774, Kp_23__N_1067, n62052, 
        n29640, n57143, n57355, n62058, n52825, n59802, n62064, 
        n57479, n52637, n26406, n57713, n25899, n57062, n62026, 
        n2_adj_4948, n2_adj_4949, n57490, n62160, n62164, n2_adj_4950, 
        n2_adj_4952, n28052, n28054, n28056, n28058, n28060, n28062, 
        n28064, n28066, n28068, n28070, n28072, n28074, n28076, 
        n28078, n28080, n28082, n28084, n28086, n28088, n28090, 
        n28092, n28094, n28096, n28098, n28100, n28102, n28104, 
        n28106, n28108, n28110, n28112, n59141, n2_adj_4953, n2_adj_4954, 
        n2_adj_4955, n2_adj_4956, n28374, n50464, n65365, n50463, 
        n65362, n50462, n65361, n50461, n65360, n50460, n65359, 
        n50459, n65355, n50458, n65313, n50457, n65312, n50456, 
        n65311, n50455, n65307, n50454, n65297, n2_adj_4957, n50453, 
        n65290, n50452, n65286, n50451, n65284, n50450, n65282, 
        n50449, n65279, n50448, n65277, n50447, n65276, n50446, 
        n65275, n50445, n65268, n50444, n65267, n50443, n65266, 
        n59980, n57238, n50442, n65265, n50441, n65264, n50440, 
        n65263, n50439, n65262, n50438, n65261, n50437, n65260, 
        n2_adj_4958, n50436, n65259, n50435, n65258, n50434, n65257, 
        n2_adj_4959, n2_adj_4960, n52406, n57128, n2_adj_4961, n2_adj_4962, 
        n2_adj_4963, n62098, n57512, n62104, n57723, n52705, n57698, 
        n62090, n2_adj_4964, n52626, n51755, n2_adj_4965, n2_adj_4966, 
        n57223, n57401, n57442, n25938, n60027, n52572, n51706, 
        n58909, n25971, n29441, n29444, n30503, n29447, n29450, 
        n30482, n29453, n29456, n29459, n30476, n29462, n30472, 
        n29465, n30420, n29474, n2_adj_4967, n57683, n2_adj_4968, 
        n62174, n2_adj_4969, n2_adj_4970, n56177, n2_adj_4971, n30312, 
        n29998, n30001, n30004, n30007, n30010, n30013, n30016, 
        n2_adj_4972, n30019, n30025, n30028, n30031, n30034, n30037, 
        n30098;
    wire [7:0]\data_in_frame[10]_c ;   // verilog/coms.v(99[12:25])
    
    wire n30102, n30105, n30108, n30111, n30114, n30118, n30121, 
        n56257, n56273, n56283, n30136, n30139, n30142, n30146, 
        n56067, n30199, n30195, n57101, n57550, n57777, n57302, 
        n29609, n107, n51613, n26286, n29614, n6_adj_4973, n29618, 
        n26683, n61924, n29621, n61926, n57765, n57259, n61932, 
        n29629, n57738, n61938, n25820, n62012, n57134, n57707, 
        n61944, n59504, n59380, n57274, n6_adj_4974, n29632, n26266, 
        n57750, n10_adj_4975, n2_adj_4976, n40837, n2_adj_4977, n2_adj_4978, 
        n2_adj_4979, n51826, n2_adj_4980, n59024, n29651, n7_adj_4982, 
        n29505, n52745, n2_adj_4983, n52747, n2_adj_4984, n57188, 
        n57593, n12_adj_4985, n57616, n2_adj_4986, n57226, n69553, 
        n27011, n2048, n2049, n20371, n55927, \FRAME_MATCHER.i_31__N_2512 , 
        n2060, n27014, n2_adj_4987, n57474, n52234, n26815, n25889, 
        n2_adj_4988, n52607, n57576, n4_adj_4989, n57482, n25746, 
        n62292, n2_adj_4990, n57437, n2_adj_4991, n2_adj_4992, n2_adj_4993, 
        n57662, n6_adj_4994, n23938, n57229, n68333, n51600, n57209, 
        n25762, n12_adj_4995, n57602, n2_adj_4996, n2_adj_4997, n2_adj_4998, 
        n2_adj_4999, n2_adj_5000, n2_adj_5001, n2_adj_5002, n2_adj_5003, 
        n2_adj_5004, n2_adj_5005, n2_adj_5006, n2_adj_5007, n2_adj_5008, 
        n25169, n57704, Kp_23__N_1271, n25707, n26458, n57367, n10_adj_5009, 
        n18_adj_5010, n24_adj_5011, n25868, n22_adj_5012, n26_adj_5013, 
        n57522, n57262, n26_adj_5014, n57058, n24_adj_5015, n57163, 
        n57650, n25_adj_5016, n23_adj_5017, n6_adj_5018, n3_adj_5019, 
        n2_adj_5020, Kp_23__N_974, n57097, n57333, n62190, n57531, 
        n68329, n25903, n56625, n57599, n57115, n62248, n61990, 
        n61988, n61994, Kp_23__N_760, n57118, n57557, n62254, n57311, 
        n62000, n62256, n62002, n26329, Kp_23__N_799, n23942, n4_adj_5021, 
        n57206, n25804, n6_adj_5022, n26390, n25906, n57253, n14_adj_5023, 
        n57122, n15_adj_5024, n25915, n57055, n25924, n6_adj_5025, 
        Kp_23__N_869, n29655, n62080, n52662, n26470, n3_adj_5026, 
        n3_adj_5027, n3_adj_5028, n1;
    wire [2:0]r_SM_Main_2__N_3545;
    
    wire n2_adj_5029, n5, n28911, n3_adj_5030, n1_adj_5031, n1_adj_5032, 
        n1_adj_5033, n1_adj_5034, n1_adj_5035, n1_adj_5036, n1_adj_5037, 
        n2_adj_5038, n26912, n52688, n1_adj_5039, n2_adj_5040, n2_adj_5041, 
        n69207, n65479, n69336, n2_adj_5042, n62268, n2_adj_5043, 
        n2_adj_5044, n57710, n10_adj_5045, n59238, n58846, n58857, 
        n69267, n7_adj_5046, n59777, n61950, n61952, n57500, n61954, 
        n59473, n61958, n62202, n62206, n62214, n62220, n61960, 
        n59377, n62232, n59440, n61964, n59860, n59259, n62110, 
        n61970, n62170, n62116, n61974, n69213, n65421, n69330, 
        n69201, n69219, n66928, n69237, n62400, n20366, n15_adj_5047, 
        n22702, n52467, n16_adj_5048, n15_adj_5049, n62406, n8_adj_5050, 
        n14_adj_5051, n59689, n7_adj_5052, n3303, n62323, n1955, 
        n25483, n6_adj_5053, n6_adj_5054, n25401, n25580, n27585, 
        n59226, n16_adj_5055, n17_adj_5056, n25577, n10_adj_5057, 
        n25574, n14_adj_5058, n15_adj_5059, n25427, n10_adj_5060, 
        n14_adj_5061, n25513, n20_c, n19_c, n62506, n18_adj_5062, 
        n20_adj_5063, n15_adj_5064, n16_adj_5065, n17_adj_5066, n28_adj_5067, 
        n43466, n59359, n42668, n6_adj_5068, n38_adj_5069, n59867, 
        n36_adj_5070, n42, n40, n41, n39, n62846, n62847, n62844, 
        n62843, n62855, n62856, n62625, n62624, n62831, n62832, 
        n62706, n62705, n62819, n62820, n62769, n62768, n62798, 
        n62799, n62802, n62801, n62720, n62721, n62724, n62723, 
        n62729, n62867, n62868, n62709, n62708, n106, n40807, 
        n62714, n62715, n40852, n62727, n62726, n62786, n62787, 
        n62790, n62789, n62807, n62808, n62754, n28175, n62755, 
        n62753, n62829, n62828, n69303, n65477, n62825, n62826, 
        n62718, n62717, n62621, n62622, n62877, n62876, n57007, 
        n1_adj_5071, n65394, n5_adj_5072, n4_adj_5073, n28125, n62778, 
        n62779, n62777, n69531, n5_adj_5076, n69249, n7_adj_5077, 
        n65396, n27274, n4_adj_5079, n4_adj_5080, n57019, n40783, 
        n57046, n62763, n62764, n62762, n69507, n69231, n69243, 
        n69255, n28117, n62757, n62758, n62756, n69195, n28115, 
        n62748, n62749, n62747, n69225, n65497, n62772, n62773, 
        n62771, n69318, n62730, n6_adj_5084, n69312, n69528, n12_adj_5086, 
        n10_adj_5087, n11_adj_5088, n9_adj_5089, n69522, n57308, n10_adj_5090, 
        n22_adj_5091, n27_adj_5092, n26_adj_5093, n29, n31, n40822, 
        n69300, n69516, n62815, n69510, n7_adj_5096, n69288, n62818, 
        n69504, n69282, n69171, n69498, n69276, n69261, n69264, 
        n69258, n69252, n69246, n69240, n69234, n69228, n69222, 
        n69216, n69210, n69204, n69198, n69192, n69186, n69180, 
        n69486, n69174, n51364, n69168, n23_adj_5103, n33766;
    wire [2:0]r_SM_Main_2__N_3536;
    
    wire n58550, n29_adj_5105, n23_adj_5106;
    wire [24:0]o_Rx_DV_N_3488;
    
    SB_DFF data_in_frame_0___i177 (.Q(\data_in_frame[22] [0]), .C(clk16MHz), 
           .D(n29968));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i39 (.Q(\data_in_frame[4] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29967));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[23] [4]), 
            .I2(neopxl_color[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut (.I0(\data_out_frame[25] [5]), .I1(n51736), .I2(GND_net), 
            .I3(GND_net), .O(n57328));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 select_777_Select_222_i3_4_lut (.I0(n57328), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n57484), .I3(n57359), .O(n3));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_222_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 select_777_Select_187_i2_4_lut (.I0(\data_out_frame[23] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4726));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_187_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_186_i2_4_lut (.I0(\data_out_frame[23] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4727));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_186_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_185_i2_4_lut (.I0(\data_out_frame[23] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4728));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_185_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_184_i2_4_lut (.I0(\data_out_frame[23] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4729));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_184_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_183_i2_4_lut (.I0(\data_out_frame[22] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4730));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_183_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1090 (.I0(\data_out_frame[25] [3]), .I1(n51598), 
            .I2(GND_net), .I3(GND_net), .O(n51658));
    defparam i1_2_lut_adj_1090.LUT_INIT = 16'h6666;
    SB_LUT4 i14043_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n133[0]), .I2(n3470), 
            .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n28050));   // verilog/coms.v(158[12:15])
    defparam i14043_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 select_777_Select_220_i3_4_lut (.I0(n52789), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\data_out_frame[25] [2]), .I3(n51658), .O(n3_adj_4731));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_220_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 select_777_Select_182_i2_4_lut (.I0(\data_out_frame[22] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4732));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_182_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i38 (.Q(\data_in_frame[4] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29964));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_181_i2_4_lut (.I0(\data_out_frame[22] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4733));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_181_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4734), .S(n56908));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_180_i2_4_lut (.I0(\data_out_frame[22] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[4] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4735));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_180_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4736), .S(n56907));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_219_i3_4_lut (.I0(n57245), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n57392), .I3(n52665), .O(n3_adj_4737));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_219_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 select_777_Select_218_i3_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n57242), .I3(n52576), .O(n3_adj_4738));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_218_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 select_777_Select_179_i2_4_lut (.I0(\data_out_frame[22] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[3] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4739));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_179_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_178_i2_4_lut (.I0(\data_out_frame[22] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[2] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4740));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_178_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1091 (.I0(\data_out_frame[23] [1]), .I1(\data_out_frame[18] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n57668));
    defparam i1_2_lut_adj_1091.LUT_INIT = 16'h6666;
    SB_LUT4 select_777_Select_177_i2_4_lut (.I0(\data_out_frame[22] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[1] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4741));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_177_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_176_i2_4_lut (.I0(\data_out_frame[22] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[0] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4742));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_176_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_175_i2_4_lut (.I0(\data_out_frame[21] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4743));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_175_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_174_i2_4_lut (.I0(\data_out_frame[21] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4744));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_174_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1092 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[21] [5]), 
            .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4745));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1092.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1093 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[21] [4]), 
            .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4746));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1093.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_adj_1094 (.I0(\data_out_frame[23] [0]), .I1(n52657), 
            .I2(GND_net), .I3(GND_net), .O(n52576));
    defparam i1_2_lut_adj_1094.LUT_INIT = 16'h9999;
    SB_LUT4 i6_4_lut (.I0(n57668), .I1(n51745), .I2(\data_out_frame[23] [0]), 
            .I3(n52657), .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1095 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[21] [3]), 
            .I2(\current[11] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4747));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1095.LUT_INIT = 16'ha088;
    SB_LUT4 i7_4_lut (.I0(n9), .I1(n14), .I2(n57377), .I3(n57350), .O(n52789));
    defparam i7_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut (.I0(n57626), .I1(n59922), .I2(\data_out_frame[23] [3]), 
            .I3(\data_out_frame[20] [7]), .O(n51736));
    defparam i3_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 select_777_Select_170_i2_4_lut (.I0(\data_out_frame[21] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[10] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4748));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_170_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_2_lut (.I0(\data_out_frame[22] [6]), .I1(\data_out_frame[24] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n7));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(n7), .I1(n52789), .I2(n52576), .I3(n52767), 
            .O(n57392));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_169_i2_4_lut (.I0(\data_out_frame[21] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[9] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4749));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_169_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_168_i2_4_lut (.I0(\data_out_frame[21] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[8] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4750));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_168_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_167_i2_4_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4751));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_167_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1096 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20] [6]), 
            .I2(displacement[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4752));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1096.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_adj_1097 (.I0(n57609), .I1(n51598), .I2(GND_net), 
            .I3(GND_net), .O(n8_c));
    defparam i1_2_lut_adj_1097.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1098 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20] [5]), 
            .I2(displacement[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4753));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1098.LUT_INIT = 16'ha088;
    SB_LUT4 i5_4_lut (.I0(n52665), .I1(n57392), .I2(n51736), .I3(n52735), 
            .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 select_777_Select_164_i2_4_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4754));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_164_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_217_i3_4_lut (.I0(n25071), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n12), .I3(n8_c), .O(n3_adj_4755));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_217_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i3_4_lut_adj_1099 (.I0(\data_out_frame[25] [0]), .I1(n52735), 
            .I2(\data_out_frame[24] [6]), .I3(n57325), .O(n57242));
    defparam i3_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1100 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20] [3]), 
            .I2(displacement[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4756));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1100.LUT_INIT = 16'ha088;
    SB_LUT4 select_777_Select_216_i3_3_lut (.I0(n57242), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n57609), .I3(GND_net), .O(n3_adj_4757));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_216_i3_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 select_777_Select_162_i2_4_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4758));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_162_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut (.I0(n52735), .I1(\data_out_frame[25] [2]), .I2(\data_out_frame[25] [1]), 
            .I3(GND_net), .O(n57245));
    defparam i2_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1101 (.I0(n57065), .I1(n57412), .I2(n51784), 
            .I3(GND_net), .O(n25716));
    defparam i2_3_lut_adj_1101.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1102 (.I0(n59466), .I1(\data_out_frame[21] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n57295));
    defparam i1_2_lut_adj_1102.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1103 (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[23] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n57659));
    defparam i1_2_lut_adj_1103.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1104 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20] [1]), 
            .I2(displacement[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4759));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1104.LUT_INIT = 16'ha088;
    SB_LUT4 i10_4_lut (.I0(n57626), .I1(\data_out_frame[22] [5]), .I2(n57322), 
            .I3(n57350), .O(n24));
    defparam i10_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 select_777_Select_160_i2_4_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4760));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_160_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_159_i2_4_lut (.I0(\data_out_frame[19] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4761));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_159_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i8_4_lut (.I0(\data_out_frame[24] [5]), .I1(n51670), .I2(n57358), 
            .I3(n52761), .O(n22));
    defparam i8_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 select_777_Select_158_i2_4_lut (.I0(\data_out_frame[19] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4762));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_158_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut (.I0(n23668), .I1(\data_out_frame[20] [3]), .I2(n51730), 
            .I3(\data_out_frame[22] [5]), .O(n52735));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut (.I0(n17), .I1(n24), .I2(\data_out_frame[20] [1]), 
            .I3(n59054), .O(n26_c));
    defparam i12_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i13_4_lut (.I0(\data_out_frame[22] [7]), .I1(n26_c), .I2(n22), 
            .I3(n51672), .O(n59736));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n57428), .I1(n57659), .I2(\data_out_frame[24] [3]), 
            .I3(\data_out_frame[23] [0]), .O(n24_adj_4763));
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut (.I0(\data_out_frame[24] [2]), .I1(\data_out_frame[23] [1]), 
            .I2(\data_out_frame[23] [7]), .I3(\data_out_frame[24] [7]), 
            .O(n26_adj_4764));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1105 (.I0(\data_out_frame[24] [4]), .I1(n57762), 
            .I2(\data_out_frame[23] [4]), .I3(n52735), .O(n25_c));
    defparam i10_4_lut_adj_1105.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1106 (.I0(\data_out_frame[23] [5]), .I1(n24_adj_4763), 
            .I2(\data_out_frame[24] [6]), .I3(n59736), .O(n27_c));
    defparam i12_4_lut_adj_1106.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut (.I0(\data_out_frame[25] [3]), .I1(n27_c), .I2(n25_c), 
            .I3(n26_adj_4764), .O(n10_c));
    defparam i2_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1107 (.I0(\data_out_frame[25] [4]), .I1(\data_out_frame[25] [5]), 
            .I2(n57245), .I3(\data_out_frame[25] [6]), .O(n14_adj_4765));
    defparam i6_4_lut_adj_1107.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1108 (.I0(n26374), .I1(n14_adj_4765), .I2(n10_c), 
            .I3(n57283), .O(n57609));
    defparam i7_4_lut_adj_1108.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_215_i3_4_lut (.I0(n57395), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n57609), .I3(\data_out_frame[25] [0]), .O(n3_adj_4766));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_215_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i1_2_lut_adj_1109 (.I0(\data_out_frame[24] [3]), .I1(n57633), 
            .I2(GND_net), .I3(GND_net), .O(n57487));
    defparam i1_2_lut_adj_1109.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1110 (.I0(\data_out_frame[24] [2]), .I1(n25158), 
            .I2(GND_net), .I3(GND_net), .O(n57216));
    defparam i1_2_lut_adj_1110.LUT_INIT = 16'h6666;
    SB_LUT4 select_777_Select_211_i3_4_lut (.I0(n23709), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n57216), .I3(\data_out_frame[24] [1]), .O(n3_adj_4767));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_211_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_adj_1111 (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[23] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n57762));
    defparam i1_2_lut_adj_1111.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1112 (.I0(n57756), .I1(n57762), .I2(\data_out_frame[24] [0]), 
            .I3(n57647), .O(n12_adj_4768));
    defparam i5_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_210_i3_4_lut (.I0(n57137), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n12_adj_4768), .I3(n8_adj_4769), .O(n3_adj_4770));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_210_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i2_3_lut_adj_1113 (.I0(n51617), .I1(n51672), .I2(\data_out_frame[23] [5]), 
            .I3(GND_net), .O(n26374));
    defparam i2_3_lut_adj_1113.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1114 (.I0(n51640), .I1(\data_out_frame[21] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n57647));
    defparam i1_2_lut_adj_1114.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1115 (.I0(n57322), .I1(n52761), .I2(n26825), 
            .I3(n52130), .O(n15_c));
    defparam i6_4_lut_adj_1115.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1116 (.I0(n15_c), .I1(n51652), .I2(n14_adj_4771), 
            .I3(n2217), .O(n25158));
    defparam i8_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1117 (.I0(\data_out_frame[21] [7]), .I1(n52761), 
            .I2(\data_out_frame[21] [5]), .I3(GND_net), .O(n57756));
    defparam i2_3_lut_adj_1117.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1118 (.I0(n57641), .I1(\data_out_frame[23] [7]), 
            .I2(n57756), .I3(n57644), .O(n10_adj_4772));
    defparam i4_4_lut_adj_1118.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(n59521), .I1(n10_adj_4772), .I2(n52581), .I3(GND_net), 
            .O(n23709));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1119 (.I0(\data_out_frame[22] [4]), .I1(n51837), 
            .I2(GND_net), .I3(GND_net), .O(n57325));
    defparam i1_2_lut_adj_1119.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1120 (.I0(n57419), .I1(\data_out_frame[15] [6]), 
            .I2(n51676), .I3(n57422), .O(n10_adj_4773));
    defparam i4_4_lut_adj_1120.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1121 (.I0(\data_out_frame[13] [7]), .I1(n51832), 
            .I2(GND_net), .I3(GND_net), .O(n57419));
    defparam i1_2_lut_adj_1121.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1122 (.I0(n57232), .I1(\data_out_frame[20] [2]), 
            .I2(\data_out_frame[20] [4]), .I3(n57460), .O(n2217));   // verilog/coms.v(100[12:26])
    defparam i3_4_lut_adj_1122.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1123 (.I0(n51784), .I1(n26693), .I2(n26394), 
            .I3(n1699), .O(n57450));
    defparam i3_4_lut_adj_1123.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1124 (.I0(\data_out_frame[16] [2]), .I1(n57450), 
            .I2(n52803), .I3(GND_net), .O(n59193));
    defparam i2_3_lut_adj_1124.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1125 (.I0(n59193), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n57398));
    defparam i1_2_lut_adj_1125.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1126 (.I0(n2217), .I1(n52581), .I2(n23666), .I3(n6_c), 
            .O(n51670));
    defparam i4_4_lut_adj_1126.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1127 (.I0(n52767), .I1(n51670), .I2(GND_net), 
            .I3(GND_net), .O(n51605));
    defparam i1_2_lut_adj_1127.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1128 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[18] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n57305));
    defparam i1_2_lut_adj_1128.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1129 (.I0(\data_out_frame[17] [2]), .I1(\data_out_frame[17] [3]), 
            .I2(n57416), .I3(\data_out_frame[17] [1]), .O(n16));
    defparam i6_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n1951), .I3(n1954), .O(n25488));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i1_3_lut_4_lut_adj_1130 (.I0(n25696), .I1(n57590), .I2(n51682), 
            .I3(\data_out_frame[19] [5]), .O(n52581));
    defparam i1_3_lut_4_lut_adj_1130.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1131 (.I0(\data_out_frame[17] [5]), .I1(n26858), 
            .I2(n57689), .I3(\data_out_frame[16] [5]), .O(n17_adj_4774));
    defparam i7_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1132 (.I0(n17_adj_4774), .I1(\data_out_frame[17] [4]), 
            .I2(n16), .I3(n68335), .O(n60097));
    defparam i9_4_lut_adj_1132.LUT_INIT = 16'h9669;
    SB_LUT4 i52653_4_lut (.I0(n60097), .I1(\data_out_frame[14] [4]), .I2(n57305), 
            .I3(\data_out_frame[18] [5]), .O(n68339));
    defparam i52653_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1133 (.I0(n1951), .I1(n4452), .I2(n1954), 
            .I3(n1957), .O(n59002));   // verilog/coms.v(145[4] 147[7])
    defparam i2_3_lut_4_lut_adj_1133.LUT_INIT = 16'h2000;
    SB_LUT4 i4_4_lut_adj_1134 (.I0(n25696), .I1(n26253), .I2(\data_out_frame[15] [3]), 
            .I3(n6_adj_4775), .O(n51640));
    defparam i4_4_lut_adj_1134.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1135 (.I0(\data_out_frame[19] [3]), .I1(n51640), 
            .I2(GND_net), .I3(GND_net), .O(n57641));
    defparam i1_2_lut_adj_1135.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_1136 (.I0(n57345), .I1(n25679), .I2(n1668), 
            .I3(n51541), .O(n26_adj_4776));
    defparam i11_4_lut_adj_1136.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1137 (.I0(n57374), .I1(n57638), .I2(\data_out_frame[11] [0]), 
            .I3(\data_out_frame[12] [1]), .O(n24_adj_4777));
    defparam i9_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1138 (.I0(n1191), .I1(n57692), .I2(\data_out_frame[12] [2]), 
            .I3(n57596), .O(n25_adj_4778));
    defparam i10_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 i8_3_lut (.I0(\data_out_frame[12] [0]), .I1(n57729), .I2(\data_out_frame[12] [3]), 
            .I3(GND_net), .O(n23));
    defparam i8_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i14_4_lut (.I0(n23), .I1(n25_adj_4778), .I2(n24_adj_4777), 
            .I3(n26_adj_4776), .O(n58952));
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut (.I0(\data_out_frame[11] [7]), .I1(n52669), .I2(GND_net), 
            .I3(GND_net), .O(n18));
    defparam i4_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1139 (.I0(n57587), .I1(n57200), .I2(n57553), 
            .I3(\data_out_frame[6] [0]), .O(n24_adj_4779));
    defparam i10_4_lut_adj_1139.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1140 (.I0(\data_out_frame[14] [1]), .I1(n58952), 
            .I2(n57570), .I3(n57185), .O(n22_adj_4780));
    defparam i8_4_lut_adj_1140.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut_adj_1141 (.I0(n57735), .I1(n24_adj_4779), .I2(n18), 
            .I3(n25667), .O(n26_adj_4781));
    defparam i12_4_lut_adj_1141.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1142 (.I0(n25696), .I1(n57590), .I2(\data_out_frame[22] [0]), 
            .I3(\data_out_frame[19] [6]), .O(n52761));
    defparam i2_3_lut_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1143 (.I0(n25679), .I1(n26_adj_4781), .I2(n22_adj_4780), 
            .I3(\data_out_frame[13] [7]), .O(n51784));
    defparam i13_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1144 (.I0(n57140), .I1(\data_out_frame[16] [3]), 
            .I2(n51784), .I3(GND_net), .O(n52803));
    defparam i2_3_lut_adj_1144.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_4_lut (.I0(n1951), .I1(n4452), .I2(n62408), .I3(\FRAME_MATCHER.i_31__N_2514 ), 
            .O(n59835));   // verilog/coms.v(145[4] 147[7])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'ha2a0;
    SB_DFFE data_in_frame_0___i37 (.Q(\data_in_frame[4] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29959));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1145 (.I0(\data_out_frame[18] [6]), .I1(n57386), 
            .I2(n59591), .I3(\data_out_frame[18] [5]), .O(n51654));
    defparam i3_4_lut_adj_1145.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i36 (.Q(\data_in_frame[4] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29956));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i35 (.Q(\data_in_frame[4] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29953));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i178 (.Q(\data_in_frame[22] [1]), .C(clk16MHz), 
           .D(n29663));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i34 (.Q(\data_in_frame[4] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29949));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i33 (.Q(\data_in_frame[4] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29946));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_2_lut (.I0(n57741), .I1(n57412), .I2(GND_net), .I3(GND_net), 
            .O(n11));
    defparam i3_2_lut.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i32 (.Q(\data_in_frame[3] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n56355));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i2 (.Q(\data_in_frame[0] [1]), .C(clk16MHz), 
           .D(n29666));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i31 (.Q(\data_in_frame[3][6] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29939));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i30 (.Q(\data_in_frame[3][5] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29936));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_4_lut_adj_1146 (.I0(n2076), .I1(n57641), .I2(n26241), .I3(\data_out_frame[16] [5]), 
            .O(n13));
    defparam i5_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1147 (.I0(n13), .I1(n11), .I2(n52737), .I3(n25810), 
            .O(n51811));
    defparam i7_4_lut_adj_1147.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1148 (.I0(n51811), .I1(n51654), .I2(\data_out_frame[19] [5]), 
            .I3(\data_out_frame[16] [6]), .O(n16_adj_4782));
    defparam i6_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_53751 (.I0(byte_transmit_counter[3]), 
            .I1(n69177), .I2(n65441), .I3(byte_transmit_counter[4]), .O(n69480));
    defparam byte_transmit_counter_3__bdd_4_lut_53751.LUT_INIT = 16'he4aa;
    SB_LUT4 i7_4_lut_adj_1149 (.I0(n52803), .I1(n26626), .I2(n57413), 
            .I3(n57235), .O(n17_adj_4783));
    defparam i7_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 n69480_bdd_4_lut (.I0(n69480), .I1(n69279), .I2(n69315), .I3(byte_transmit_counter[4]), 
            .O(tx_data[3]));
    defparam n69480_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9_4_lut_adj_1150 (.I0(n17_adj_4783), .I1(n57606), .I2(n16_adj_4782), 
            .I3(n57065), .O(n23666));
    defparam i9_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_53736 (.I0(byte_transmit_counter[3]), 
            .I1(n69183), .I2(n65454), .I3(byte_transmit_counter[4]), .O(n69474));
    defparam byte_transmit_counter_3__bdd_4_lut_53736.LUT_INIT = 16'he4aa;
    SB_LUT4 n69474_bdd_4_lut (.I0(n69474), .I1(n69291), .I2(n7_adj_4784), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n69474_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_53731 (.I0(byte_transmit_counter[3]), 
            .I1(n69189), .I2(n65442), .I3(byte_transmit_counter[4]), .O(n69468));
    defparam byte_transmit_counter_3__bdd_4_lut_53731.LUT_INIT = 16'he4aa;
    SB_LUT4 n69468_bdd_4_lut (.I0(n69468), .I1(n69285), .I2(n7_adj_4785), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n69468_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1151 (.I0(n23666), .I1(\data_out_frame[22] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26825));
    defparam i1_2_lut_adj_1151.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_53726 (.I0(byte_transmit_counter[3]), 
            .I1(n67511), .I2(n65487), .I3(byte_transmit_counter[4]), .O(n69462));
    defparam byte_transmit_counter_3__bdd_4_lut_53726.LUT_INIT = 16'he4aa;
    SB_LUT4 n69462_bdd_4_lut (.I0(n69462), .I1(n14_adj_4786), .I2(n7_adj_4787), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n69462_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFE data_in_frame_0___i29 (.Q(\data_in_frame[3][4] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29933));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1152 (.I0(\data_out_frame[20] [5]), .I1(n51730), 
            .I2(GND_net), .I3(GND_net), .O(n52665));
    defparam i1_2_lut_adj_1152.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i179 (.Q(\data_in_frame[22] [2]), .C(clk16MHz), 
           .D(n29669));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i28 (.Q(\data_in_frame[3][3] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29929));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i27 (.Q(\data_in_frame[3][2] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29926));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1153 (.I0(n52665), .I1(n59153), .I2(n51837), 
            .I3(n26825), .O(n10_adj_4788));
    defparam i4_4_lut_adj_1153.LUT_INIT = 16'h9669;
    SB_LUT4 i3_2_lut_adj_1154 (.I0(n57422), .I1(\data_out_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4789));
    defparam i3_2_lut_adj_1154.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1155 (.I0(n25095), .I1(n10_adj_4789), .I2(n52737), 
            .I3(n57446), .O(n12_adj_4790));
    defparam i5_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1156 (.I0(\data_out_frame[13] [5]), .I1(n12_adj_4790), 
            .I2(n57446), .I3(\data_out_frame[17] [7]), .O(n52164));
    defparam i6_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i26 (.Q(\data_in_frame[3][1] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29923));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1157 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[18] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n57456));
    defparam i1_2_lut_adj_1157.LUT_INIT = 16'h6666;
    SB_DFFE data_in_frame_0___i25 (.Q(\data_in_frame[3][0] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29920));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i24 (.Q(\data_in_frame[2] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29917));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i180 (.Q(\data_in_frame[22] [3]), .C(clk16MHz), 
           .D(n29674));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i23 (.Q(\data_in_frame[2] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29913));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i22 (.Q(\data_in_frame[2] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29910));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i3 (.Q(\data_in_frame[0] [2]), .C(clk16MHz), 
           .D(n29678));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1158 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n57689));
    defparam i1_2_lut_adj_1158.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1159 (.I0(n57456), .I1(n51676), .I2(n52164), 
            .I3(n57560), .O(n10_adj_4791));
    defparam i4_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1160 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n57747));
    defparam i1_2_lut_adj_1160.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1161 (.I0(n51676), .I1(n57590), .I2(\data_out_frame[22] [2]), 
            .I3(n25734), .O(n12_adj_4792));
    defparam i5_4_lut_adj_1161.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1162 (.I0(\data_out_frame[20] [0]), .I1(n12_adj_4792), 
            .I2(n57747), .I3(\data_out_frame[17] [6]), .O(n59153));
    defparam i6_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1163 (.I0(\data_out_frame[15] [3]), .I1(n26253), 
            .I2(n25734), .I3(\data_out_frame[17] [5]), .O(n57131));
    defparam i3_4_lut_adj_1163.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1164 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[19] [7]), 
            .I2(n57131), .I3(n6_adj_4793), .O(n52130));
    defparam i4_4_lut_adj_1164.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1165 (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[22] [3]), 
            .I2(n52130), .I3(GND_net), .O(n59054));
    defparam i2_3_lut_adj_1165.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1166 (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[20] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n57460));
    defparam i1_2_lut_adj_1166.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1167 (.I0(n52164), .I1(\data_out_frame[18] [1]), 
            .I2(n52327), .I3(GND_net), .O(n23668));
    defparam i2_3_lut_adj_1167.LUT_INIT = 16'h9696;
    SB_LUT4 i24102_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n22726), .I3(GND_net), .O(n29692));
    defparam i24102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24103_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n22726), .I3(GND_net), .O(n29693));
    defparam i24103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[11] [1]), .I1(n51720), .I2(\data_in_frame[17] [7]), 
            .I3(n10_adj_4794), .O(n25128));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1168 (.I0(\data_out_frame[25] [7]), .I1(n26374), 
            .I2(\data_out_frame[24] [0]), .I3(GND_net), .O(n57283));
    defparam i2_3_lut_adj_1168.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_in_frame[11] [1]), .I1(n51720), .I2(\data_in_frame[8] [6]), 
            .I3(GND_net), .O(n57404));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_4_lut (.I0(n25853), .I1(n59043), .I2(\data_in_frame[9] [0]), 
            .I3(n57352), .O(n6_adj_4795));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut (.I0(n25853), .I1(n59043), .I2(\data_in_frame[9] [0]), 
            .I3(Kp_23__N_1080), .O(n57331));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1169 (.I0(n57633), .I1(n57283), .I2(n25105), 
            .I3(n52618), .O(n12_adj_4796));
    defparam i5_4_lut_adj_1169.LUT_INIT = 16'h9669;
    SB_LUT4 select_777_Select_209_i3_4_lut (.I0(n25158), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n12_adj_4796), .I3(n8_adj_4797), .O(n3_adj_4798));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_209_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_adj_1170 (.I0(\data_out_frame[21] [4]), .I1(n26626), 
            .I2(GND_net), .I3(GND_net), .O(n57771));
    defparam i1_2_lut_adj_1170.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1171 (.I0(n26428), .I1(n4_c), .I2(n57573), 
            .I3(n26724), .O(n62074));   // verilog/coms.v(77[16:43])
    defparam i1_3_lut_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1172 (.I0(n57072), .I1(n57425), .I2(\data_out_frame[12] [7]), 
            .I3(\data_out_frame[10] [7]), .O(n12_adj_4799));   // verilog/coms.v(77[16:43])
    defparam i5_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_157_i2_4_lut (.I0(\data_out_frame[19] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4800));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_157_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i6_4_lut_adj_1173 (.I0(n36), .I1(n12_adj_4799), .I2(n57695), 
            .I3(n26423), .O(n26253));   // verilog/coms.v(77[16:43])
    defparam i6_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1174 (.I0(n26428), .I1(n4_c), .I2(\data_in_frame[10] [4]), 
            .I3(GND_net), .O(n26031));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1174.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_156_i2_4_lut (.I0(\data_out_frame[19] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4801));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_156_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1175 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[19] [3]), 
            .I2(displacement[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4802));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1175.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[1] [7]), .O(n57732));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1176 (.I0(n51619), .I1(n26253), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4803));
    defparam i1_2_lut_adj_1176.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1177 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[3][5] ), .I3(GND_net), .O(n26415));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut_adj_1177.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1178 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(\data_out_frame[15] [1]), .I3(n6_adj_4803), .O(n51682));
    defparam i4_4_lut_adj_1178.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1179 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[19] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n57386));
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1180 (.I0(n25068), .I1(\data_out_frame[14] [3]), 
            .I2(\data_out_frame[12] [1]), .I3(GND_net), .O(n57412));
    defparam i2_3_lut_adj_1180.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1181 (.I0(\data_out_frame[16] [3]), .I1(n26100), 
            .I2(\data_out_frame[16] [5]), .I3(\data_out_frame[16] [7]), 
            .O(n25918));   // verilog/coms.v(88[17:28])
    defparam i3_4_lut_adj_1181.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1182 (.I0(\data_out_frame[16] [6]), .I1(n25918), 
            .I2(n57280), .I3(\data_out_frame[16] [4]), .O(n57446));   // verilog/coms.v(88[17:28])
    defparam i3_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_154_i2_4_lut (.I0(\data_out_frame[19] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4804));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_154_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_153_i2_4_lut (.I0(\data_out_frame[19] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4805));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_153_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1183 (.I0(\data_out_frame[15] [5]), .I1(n26257), 
            .I2(n51676), .I3(GND_net), .O(n57416));
    defparam i2_3_lut_adj_1183.LUT_INIT = 16'h9696;
    SB_LUT4 i52649_4_lut (.I0(n52737), .I1(n57413), .I2(n57446), .I3(n51753), 
            .O(n68335));
    defparam i52649_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1184 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26100));
    defparam i1_2_lut_adj_1184.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1185 (.I0(n52737), .I1(n68335), .I2(GND_net), 
            .I3(GND_net), .O(n57171));
    defparam i1_2_lut_adj_1185.LUT_INIT = 16'h6666;
    SB_LUT4 i1288_2_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n2076));   // verilog/coms.v(88[17:28])
    defparam i1288_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1186 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[15] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n25734));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1186.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1187 (.I0(\data_in_frame[6] [7]), .I1(n25797), 
            .I2(n57289), .I3(n26332), .O(n26298));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_4_lut_adj_1187.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1188 (.I0(\data_out_frame[15] [1]), .I1(\data_out_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n57104));
    defparam i1_2_lut_adj_1188.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1189 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n57181));
    defparam i1_2_lut_adj_1189.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1190 (.I0(\data_out_frame[14] [4]), .I1(n26241), 
            .I2(GND_net), .I3(GND_net), .O(n57235));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1190.LUT_INIT = 16'h6666;
    SB_LUT4 select_777_Select_110_i2_4_lut (.I0(\data_out_frame[13] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4806));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_110_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1191 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n25679));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1191.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1192 (.I0(\data_out_frame[10] [4]), .I1(n57656), 
            .I2(n57653), .I3(n57547), .O(n59779));   // verilog/coms.v(75[16:27])
    defparam i3_4_lut_adj_1192.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1193 (.I0(\data_out_frame[14] [6]), .I1(n1516), 
            .I2(n59779), .I3(n25679), .O(n26757));
    defparam i3_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1194 (.I0(\data_in_frame[2] [0]), .I1(n57567), 
            .I2(n26363), .I3(\data_in_frame[6][5] ), .O(n57108));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_4_lut_adj_1194.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1195 (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n57553));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1195.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1196 (.I0(n57111), .I1(\data_out_frame[8] [0]), 
            .I2(n57622), .I3(n57553), .O(n10_adj_4807));   // verilog/coms.v(77[16:27])
    defparam i4_4_lut_adj_1196.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1197 (.I0(\data_out_frame[10] [0]), .I1(n10_adj_4807), 
            .I2(\data_out_frame[10] [1]), .I3(GND_net), .O(n57753));   // verilog/coms.v(77[16:27])
    defparam i5_3_lut_adj_1197.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1198 (.I0(n57090), .I1(n57759), .I2(\data_out_frame[6] [0]), 
            .I3(GND_net), .O(n57547));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1198.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1199 (.I0(\data_in_frame[2] [0]), .I1(n57567), 
            .I2(n26363), .I3(Kp_23__N_872), .O(n6_adj_4808));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_4_lut_adj_1199.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1200 (.I0(n57596), .I1(\data_out_frame[11] [0]), 
            .I2(n25671), .I3(GND_net), .O(n57425));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1200.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1201 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[12] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n57200));
    defparam i1_2_lut_adj_1201.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1202 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[4] [2]), .I3(GND_net), .O(n57150));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1202.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_109_i2_4_lut (.I0(\data_out_frame[13] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4809));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_109_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1203 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4810));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1203.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1204 (.I0(n57154), .I1(n26066), .I2(\data_out_frame[11] [7]), 
            .I3(n6_adj_4810), .O(n25068));   // verilog/coms.v(79[16:43])
    defparam i4_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_108_i2_4_lut (.I0(\data_out_frame[13] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4811));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_108_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_2_lut_adj_1205 (.I0(n25068), .I1(n57200), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4812));
    defparam i2_2_lut_adj_1205.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1206 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[12] [0]), 
            .I2(n57265), .I3(n1563), .O(n14_adj_4813));
    defparam i6_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i21 (.Q(\data_in_frame[2] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29906));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i7_4_lut_adj_1207 (.I0(\data_out_frame[14] [2]), .I1(n14_adj_4813), 
            .I2(n10_adj_4812), .I3(n57622), .O(n57140));
    defparam i7_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1208 (.I0(\data_out_frame[14] [4]), .I1(n57140), 
            .I2(GND_net), .I3(GND_net), .O(n51805));
    defparam i1_2_lut_adj_1208.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4814), .S(n56906));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1209 (.I0(\data_out_frame[14] [0]), .I1(n57265), 
            .I2(\data_out_frame[11] [6]), .I3(n26066), .O(n26693));
    defparam i3_4_lut_adj_1209.LUT_INIT = 16'h6996;
    SB_LUT4 i880_2_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1668));   // verilog/coms.v(88[17:28])
    defparam i880_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1210 (.I0(\data_out_frame[8] [2]), .I1(n1668), 
            .I2(\data_out_frame[10] [4]), .I3(\data_out_frame[8] [3]), .O(n57735));   // verilog/coms.v(77[16:27])
    defparam i3_4_lut_adj_1210.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1211 (.I0(n26607), .I1(\data_out_frame[13] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n57695));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1211.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1212 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(n26335), .I3(GND_net), .O(n57157));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut_adj_1212.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[4] [1]), .I3(\data_in_frame[3] [7]), .O(n57160));   // verilog/coms.v(73[16:69])
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4815), .S(n56905));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1213 (.I0(n57564), .I1(n57146), .I2(n57735), 
            .I3(n6_adj_4816), .O(n51656));   // verilog/coms.v(77[16:27])
    defparam i4_4_lut_adj_1213.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1214 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n57374));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1214.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1215 (.I0(n57744), .I1(\data_out_frame[6] [7]), 
            .I2(n57374), .I3(n36), .O(n14_adj_4817));   // verilog/coms.v(88[17:28])
    defparam i6_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1216 (.I0(\data_out_frame[13] [3]), .I1(n14_adj_4817), 
            .I2(n10_adj_4818), .I3(\data_out_frame[8] [7]), .O(n26257));   // verilog/coms.v(88[17:28])
    defparam i7_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1217 (.I0(n57528), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[11] [1]), .I3(n57052), .O(n15_adj_4819));   // verilog/coms.v(100[12:26])
    defparam i6_4_lut_adj_1217.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1218 (.I0(n15_adj_4819), .I1(\data_out_frame[9] [0]), 
            .I2(n14_adj_4820), .I3(\data_out_frame[8] [7]), .O(n25696));   // verilog/coms.v(100[12:26])
    defparam i8_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1219 (.I0(\data_out_frame[8] [6]), .I1(n57146), 
            .I2(GND_net), .I3(GND_net), .O(n36));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1219.LUT_INIT = 16'h6666;
    SB_LUT4 i911_2_lut (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1699));   // verilog/coms.v(74[16:27])
    defparam i911_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1220 (.I0(n57248), .I1(n36), .I2(\data_out_frame[13] [4]), 
            .I3(n57613), .O(n10_adj_4821));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_LUT4 add_1099_9_lut (.I0(n56736), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n49184), .O(n56737)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1099_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1221 (.I0(n25696), .I1(n26257), .I2(GND_net), 
            .I3(GND_net), .O(n1720));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1221.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1222 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n57528));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1222.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1223 (.I0(n57203), .I1(n57178), .I2(n26524), 
            .I3(\data_out_frame[7] [1]), .O(n10_adj_4822));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1223.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1224 (.I0(\data_out_frame[6] [7]), .I1(n10_adj_4822), 
            .I2(\data_out_frame[4] [7]), .I3(GND_net), .O(n51541));   // verilog/coms.v(88[17:70])
    defparam i5_3_lut_adj_1224.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1225 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n57203));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1225.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4823), .S(n56952));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1226 (.I0(n57581), .I1(n26083), .I2(\data_out_frame[9] [2]), 
            .I3(n57744), .O(n10_adj_4824));
    defparam i4_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1227 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6][5] ), 
            .I2(n26332), .I3(Kp_23__N_878), .O(n57271));   // verilog/coms.v(80[16:43])
    defparam i2_3_lut_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1228 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[10] [3]), 
            .I2(\data_out_frame[10] [4]), .I3(GND_net), .O(n57314));   // verilog/coms.v(88[17:63])
    defparam i2_3_lut_adj_1228.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1229 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6][5] ), 
            .I2(\data_in_frame[6][4] ), .I3(GND_net), .O(n57619));   // verilog/coms.v(80[16:43])
    defparam i1_2_lut_3_lut_adj_1229.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1230 (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n57638));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1230.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1231 (.I0(\data_in_frame[1] [5]), .I1(n57732), 
            .I2(n26193), .I3(GND_net), .O(n57726));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_3_lut_adj_1231.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_152_i2_4_lut (.I0(\data_out_frame[19] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4825));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_152_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1232 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26662));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1232.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1233 (.I0(\data_in_frame[1] [5]), .I1(n57732), 
            .I2(\data_in_frame[1] [0]), .I3(n25893), .O(n35660));   // verilog/coms.v(73[16:69])
    defparam i1_3_lut_4_lut_adj_1233.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1234 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[4] [3]), .I3(GND_net), .O(n57146));   // verilog/coms.v(100[12:26])
    defparam i2_3_lut_adj_1234.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1235 (.I0(n25671), .I1(n57146), .I2(\data_out_frame[8] [5]), 
            .I3(GND_net), .O(n26423));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1235.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1236 (.I0(\data_out_frame[9] [1]), .I1(n26423), 
            .I2(GND_net), .I3(GND_net), .O(n57665));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1236.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1237 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n57613));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1237.LUT_INIT = 16'h6666;
    SB_LUT4 i775_2_lut (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1563));   // verilog/coms.v(74[16:27])
    defparam i775_2_lut.LUT_INIT = 16'h6666;
    SB_DFFR \FRAME_MATCHER.state_FSM_i1  (.Q(Kp_23__N_1748), .C(clk16MHz), 
            .D(n2068), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFE data_in_frame_0___i20 (.Q(\data_in_frame[2] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29903));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i0 (.Q(setpoint[0]), .C(clk16MHz), .E(n27737), 
            .D(n4762[0]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1238 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n57759));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_adj_1238.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_in_frame[4] [5]), .I1(n57271), .I2(\data_in_frame[8] [7]), 
            .I3(GND_net), .O(n7_adj_4826));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1239 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[7] [1]), 
            .I2(\data_out_frame[8] [7]), .I3(GND_net), .O(n57792));   // verilog/coms.v(74[16:62])
    defparam i2_3_lut_adj_1239.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1240 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n57656));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_adj_1240.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1241 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n57084));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_adj_1241.LUT_INIT = 16'h6666;
    SB_LUT4 select_777_Select_151_i2_4_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4827));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_151_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_3_lut_4_lut_adj_1242 (.I0(n59636), .I1(n57441), .I2(\data_in_frame[22] [6]), 
            .I3(\data_in_frame[20] [4]), .O(n8_adj_4828));
    defparam i3_3_lut_4_lut_adj_1242.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1243 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n57581));
    defparam i1_2_lut_adj_1243.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1244 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n57789));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_adj_1244.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1245 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n57248));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1245.LUT_INIT = 16'h6666;
    SB_LUT4 i342_2_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1130));   // verilog/coms.v(79[16:27])
    defparam i342_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1246 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n57178));
    defparam i1_2_lut_adj_1246.LUT_INIT = 16'h6666;
    SB_LUT4 select_777_Select_107_i2_4_lut (.I0(\data_out_frame[13] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4829));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_107_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14904_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n28912));   // verilog/coms.v(130[12] 305[6])
    defparam i14904_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_DFF data_in_frame_0___i181 (.Q(\data_in_frame[22] [4]), .C(clk16MHz), 
           .D(n56031));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1247 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[20] [7]), 
            .I2(\data_in_frame[18] [4]), .I3(GND_net), .O(n4_adj_4830));
    defparam i1_2_lut_3_lut_adj_1247.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1248 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[20] [7]), 
            .I2(\data_in_frame[21] [6]), .I3(\data_in_frame[21] [7]), .O(n62128));
    defparam i1_2_lut_3_lut_4_lut_adj_1248.LUT_INIT = 16'h6996;
    SB_LUT4 i16343_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in[3] [7]), .O(n30351));   // verilog/coms.v(130[12] 305[6])
    defparam i16343_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_777_Select_106_i2_4_lut (.I0(\data_out_frame[13] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4831));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_106_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 add_1099_8_lut (.I0(n56736), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n49183), .O(n56743)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1099_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i9_4_lut_adj_1249 (.I0(n1130), .I1(n57516), .I2(n57564), .I3(n57248), 
            .O(n22_adj_4832));
    defparam i9_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1250 (.I0(n57581), .I1(n25667), .I2(\data_out_frame[4] [4]), 
            .I3(n57084), .O(n21_c));
    defparam i8_4_lut_adj_1250.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1251 (.I0(\data_out_frame[6] [4]), .I1(n26607), 
            .I2(\data_out_frame[6] [1]), .I3(n14_adj_4833), .O(n23_adj_4834));
    defparam i10_4_lut_adj_1251.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1252 (.I0(n23_adj_4834), .I1(n57789), .I2(n21_c), 
            .I3(n22_adj_4832), .O(n24_adj_4835));   // verilog/coms.v(74[16:62])
    defparam i7_4_lut_adj_1252.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1253 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [6]), 
            .I2(displacement[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4836));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1253.LUT_INIT = 16'ha088;
    SB_LUT4 i15642_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [0]), 
            .I3(\data_in[0] [0]), .O(n29650));   // verilog/coms.v(130[12] 305[6])
    defparam i15642_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_777_Select_149_i2_4_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4837));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_149_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16374_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [1]), 
            .I3(\data_in[0] [1]), .O(n30382));   // verilog/coms.v(130[12] 305[6])
    defparam i16374_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_777_Select_148_i2_4_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4838));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_148_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i19 (.Q(\data_in_frame[2] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29899));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13_4_lut_adj_1254 (.I0(n57656), .I1(\data_out_frame[7] [4]), 
            .I2(n57084), .I3(n18_adj_4839), .O(n30_c));   // verilog/coms.v(74[16:62])
    defparam i13_4_lut_adj_1254.LUT_INIT = 16'h6996;
    SB_LUT4 i16373_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [2]), 
            .I3(\data_in[0] [2]), .O(n30381));   // verilog/coms.v(130[12] 305[6])
    defparam i16373_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11_4_lut_adj_1255 (.I0(\data_out_frame[7] [5]), .I1(n57792), 
            .I2(n57342), .I3(\data_out_frame[7] [2]), .O(n28));   // verilog/coms.v(74[16:62])
    defparam i11_4_lut_adj_1255.LUT_INIT = 16'h6996;
    SB_CARRY add_1099_8 (.CI(n49183), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n49184));
    SB_LUT4 i15_4_lut (.I0(n57759), .I1(n30_c), .I2(n24_adj_4835), .I3(\data_out_frame[8] [6]), 
            .O(n32_c));   // verilog/coms.v(74[16:62])
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1256 (.I0(n57613), .I1(n57665), .I2(\data_out_frame[9] [7]), 
            .I3(n57587), .O(n27_adj_4840));   // verilog/coms.v(74[16:62])
    defparam i10_4_lut_adj_1256.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1257 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4841));
    defparam i2_2_lut_adj_1257.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1258 (.I0(n27_adj_4840), .I1(n1563), .I2(n32_c), 
            .I3(n28), .O(n7_adj_4842));
    defparam i1_4_lut_adj_1258.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_4_lut_adj_1259 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[20] [7]), 
            .I2(n51588), .I3(n10_adj_4843), .O(n59162));
    defparam i5_3_lut_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1260 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [3]), 
            .I2(displacement[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4844));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1260.LUT_INIT = 16'ha088;
    SB_LUT4 add_1099_7_lut (.I0(n56736), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n49182), .O(n56742)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1099_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i5_4_lut_adj_1261 (.I0(n26662), .I1(n7_adj_4842), .I2(n26423), 
            .I3(n8_adj_4841), .O(n57692));
    defparam i5_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_CARRY add_1099_7 (.CI(n49182), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n49183));
    SB_LUT4 i1_2_lut_adj_1262 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n57584));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1262.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4845), .S(n56904));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1263 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n26607));
    defparam i2_3_lut_adj_1263.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1264 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n57175));
    defparam i1_2_lut_adj_1264.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1265 (.I0(n57175), .I1(n26607), .I2(\data_out_frame[9] [1]), 
            .I3(n57584), .O(n10_adj_4846));   // verilog/coms.v(88[17:28])
    defparam i4_4_lut_adj_1265.LUT_INIT = 16'h6996;
    SB_LUT4 i16372_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [3]), 
            .I3(\data_in[0] [3]), .O(n30380));   // verilog/coms.v(130[12] 305[6])
    defparam i16372_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16371_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [4]), 
            .I3(\data_in[0] [4]), .O(n30379));   // verilog/coms.v(130[12] 305[6])
    defparam i16371_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1266 (.I0(\data_out_frame[13] [5]), .I1(n25095), 
            .I2(GND_net), .I3(GND_net), .O(n26780));
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4847), .S(n56773));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i18 (.Q(\data_in_frame[2] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29896));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4848), .S(n56903));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_2_lut_adj_1267 (.I0(\data_out_frame[8] [3]), .I1(n57692), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4849));   // verilog/coms.v(88[17:63])
    defparam i2_2_lut_adj_1267.LUT_INIT = 16'h6666;
    SB_LUT4 i16370_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [5]), 
            .I3(\data_in[0] [5]), .O(n30378));   // verilog/coms.v(130[12] 305[6])
    defparam i16370_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_1268 (.I0(n57638), .I1(\data_out_frame[10] [2]), 
            .I2(\data_out_frame[11] [5]), .I3(n57314), .O(n14_adj_4850));   // verilog/coms.v(88[17:63])
    defparam i6_4_lut_adj_1268.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1269 (.I0(n57425), .I1(n14_adj_4850), .I2(n10_adj_4849), 
            .I3(\data_out_frame[11] [1]), .O(n52669));   // verilog/coms.v(88[17:63])
    defparam i7_4_lut_adj_1269.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_146_i2_4_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4851));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_146_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13_4_lut_adj_1270 (.I0(n57528), .I1(n1720), .I2(n51676), 
            .I3(n1699), .O(n34));
    defparam i13_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 i16369_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [6]), 
            .I3(\data_in[0] [6]), .O(n30377));   // verilog/coms.v(130[12] 305[6])
    defparam i16369_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i17_4_lut (.I0(n51832), .I1(n34), .I2(n24_adj_4852), .I3(\data_out_frame[8] [5]), 
            .O(n38));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1271 (.I0(\data_out_frame[10] [5]), .I1(n52624), 
            .I2(n52669), .I3(n26780), .O(n36_adj_4853));
    defparam i15_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i16368_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [7]), 
            .I3(\data_in[0] [7]), .O(n30376));   // verilog/coms.v(130[12] 305[6])
    defparam i16368_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_777_Select_145_i2_4_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4854));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_145_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16366_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [0]), 
            .I3(\data_in[1] [0]), .O(n30374));   // verilog/coms.v(130[12] 305[6])
    defparam i16366_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16_4_lut (.I0(\data_out_frame[14] [6]), .I1(n51805), .I2(n57280), 
            .I3(n22_adj_4855), .O(n37));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_144_i2_4_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4856));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_144_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14_4_lut_adj_1272 (.I0(\data_out_frame[14] [3]), .I1(n57547), 
            .I2(n57753), .I3(n57314), .O(n35));
    defparam i14_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1273 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[13] [5]), 
            .I2(n25095), .I3(\data_out_frame[15] [6]), .O(n6_adj_4793));
    defparam i1_2_lut_3_lut_4_lut_adj_1273.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1274 (.I0(n57181), .I1(n57280), .I2(\data_out_frame[15] [7]), 
            .I3(n57104), .O(n12_adj_4857));
    defparam i5_4_lut_adj_1274.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(n35), .I1(n37), .I2(n36_adj_4853), .I3(n38), 
            .O(n59907));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1275 (.I0(n59907), .I1(n12_adj_4857), .I2(n57560), 
            .I3(n25734), .O(n51753));
    defparam i6_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1276 (.I0(n26858), .I1(n26757), .I2(GND_net), 
            .I3(GND_net), .O(n57137));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1276.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_4_lut_adj_1277 (.I0(\FRAME_MATCHER.i_31__N_2511 ), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(n33763), .O(n6_adj_4858));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_4_lut_adj_1277.LUT_INIT = 16'hfffe;
    SB_LUT4 i14893_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(GND_net), .I3(GND_net), .O(n28901));   // verilog/coms.v(130[12] 305[6])
    defparam i14893_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3_4_lut_adj_1278 (.I0(\data_out_frame[16] [4]), .I1(n51753), 
            .I2(\data_out_frame[18] [7]), .I3(\data_out_frame[19] [1]), 
            .O(n57674));
    defparam i3_4_lut_adj_1278.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1279 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[5] [7]), .I3(GND_net), .O(n57191));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1279.LUT_INIT = 16'h9696;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(74[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16365_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [1]), 
            .I3(\data_in[1] [1]), .O(n30373));   // verilog/coms.v(130[12] 305[6])
    defparam i16365_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_777_Select_143_i2_4_lut (.I0(\data_out_frame[17] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4859));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_143_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1280 (.I0(\data_out_frame[14] [7]), .I1(n57191), 
            .I2(\data_out_frame[12] [5]), .I3(GND_net), .O(n57786));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1280.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_142_i2_4_lut (.I0(\data_out_frame[17] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4860));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_142_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1281 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n57111));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1281.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1282 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n57072));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1282.LUT_INIT = 16'h6666;
    SB_LUT4 i16364_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [2]), .O(n30372));   // verilog/coms.v(130[12] 305[6])
    defparam i16364_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16363_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [3]), 
            .I3(\data_in[1] [3]), .O(n30371));   // verilog/coms.v(130[12] 305[6])
    defparam i16363_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_777_Select_141_i2_4_lut (.I0(\data_out_frame[17] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4861));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_141_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_140_i2_4_lut (.I0(\data_out_frame[17] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4862));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_140_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16362_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [4]), .O(n30370));   // verilog/coms.v(130[12] 305[6])
    defparam i16362_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1283 (.I0(n52017), .I1(\data_in_frame[16] [5]), 
            .I2(n52655), .I3(\data_in_frame[16] [4]), .O(n51281));
    defparam i2_3_lut_4_lut_adj_1283.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_adj_1284 (.I0(n52017), .I1(\data_in_frame[16] [5]), 
            .I2(n57686), .I3(n52653), .O(n8_adj_4863));
    defparam i3_3_lut_4_lut_adj_1284.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4864), .S(n56902));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4865), .S(n56901));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4866), .S(n56900));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4867), .S(n56899));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4868), .S(n56898));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4869), .S(n56897));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4870), .S(n56896));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4871), .S(n56895));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4872), .S(n56894));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4873), .S(n56893));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4874), .S(n56892));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4875), .S(n56891));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4876), .S(n56890));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4877), .S(n56889));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4878), .S(n56888));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1285 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n57090));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1285.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4879), .S(n56887));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 add_1099_6_lut (.I0(n56736), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n49181), .O(n56741)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1099_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1286 (.I0(n25667), .I1(n25671), .I2(\data_out_frame[8] [2]), 
            .I3(\data_out_frame[10] [3]), .O(n57729));   // verilog/coms.v(75[16:27])
    defparam i3_4_lut_adj_1286.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1287 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n57345));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1287.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1288 (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n57570));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1288.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1289 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[8] [0]), 
            .I2(\data_out_frame[8] [2]), .I3(GND_net), .O(n57342));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1289.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_139_i2_4_lut (.I0(\data_out_frame[17] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4880));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_139_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1290 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n57653));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1290.LUT_INIT = 16'h6666;
    SB_LUT4 i16360_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [6]), 
            .I3(\data_in[1] [6]), .O(n30368));   // verilog/coms.v(130[12] 305[6])
    defparam i16360_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16359_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [7]), 
            .I3(\data_in[1] [7]), .O(n30367));   // verilog/coms.v(130[12] 305[6])
    defparam i16359_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16358_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [0]), 
            .I3(\data_in[2] [0]), .O(n30366));   // verilog/coms.v(130[12] 305[6])
    defparam i16358_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1291 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [4]), 
            .I2(n57342), .I3(n6_adj_4881), .O(n1516));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1291.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1292 (.I0(n52017), .I1(\data_in_frame[16] [5]), 
            .I2(n57408), .I3(GND_net), .O(n51588));
    defparam i2_2_lut_3_lut_adj_1292.LUT_INIT = 16'h9696;
    SB_LUT4 i16357_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [1]), 
            .I3(\data_in[2] [1]), .O(n30365));   // verilog/coms.v(130[12] 305[6])
    defparam i16357_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16356_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [2]), 
            .I3(\data_in[2] [2]), .O(n30364));   // verilog/coms.v(130[12] 305[6])
    defparam i16356_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1293 (.I0(\data_out_frame[8] [1]), .I1(n25731), 
            .I2(n57154), .I3(n6_adj_4882), .O(n26241));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1293.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1294 (.I0(\data_out_frame[14] [5]), .I1(n26241), 
            .I2(n1516), .I3(\data_out_frame[12] [4]), .O(n57280));
    defparam i1_4_lut_adj_1294.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut (.I0(n57786), .I1(\data_out_frame[5] [5]), .I2(n1191), 
            .I3(GND_net), .O(n11_adj_4883));   // verilog/coms.v(75[16:27])
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1295 (.I0(\data_out_frame[12] [6]), .I1(n57729), 
            .I2(n57090), .I3(\data_out_frame[7] [7]), .O(n13_adj_4884));   // verilog/coms.v(75[16:27])
    defparam i5_4_lut_adj_1295.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_4_lut_4_lut (.I0(n28399), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n56297));
    defparam i1_4_lut_4_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1296 (.I0(n13_adj_4884), .I1(n11_adj_4883), .I2(n57072), 
            .I3(\data_out_frame[8] [1]), .O(n51619));   // verilog/coms.v(75[16:27])
    defparam i7_4_lut_adj_1296.LUT_INIT = 16'h6996;
    SB_LUT4 i16355_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [3]), 
            .I3(\data_in[2] [3]), .O(n30363));   // verilog/coms.v(130[12] 305[6])
    defparam i16355_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1297 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4885));
    defparam i1_2_lut_adj_1297.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1298 (.I0(n51619), .I1(\data_out_frame[15] [0]), 
            .I2(n57280), .I3(n6_adj_4885), .O(n57317));
    defparam i4_4_lut_adj_1298.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_138_i2_4_lut (.I0(\data_out_frame[17] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4886));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_138_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4887), .S(n56886));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4888), .S(n56885));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4889), .S(n56884));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4890), .S(n56883));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4891), .S(n56882));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4892), .S(n56881));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4893), .S(n56880));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1299 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26272));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1299.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4894), .S(n56879));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4895), .S(n56878));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4896), .S(n56877));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4897), .S(n56876));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4898), .S(n56875));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4899), .S(n56874));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4900), .S(n56873));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk16MHz), 
            .E(n30569), .D(n2_adj_4901), .S(n29046));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i17 (.Q(\data_in_frame[2] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29893));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4902), .S(n56872));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i16354_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [4]), 
            .I3(\data_in[2] [4]), .O(n30362));   // verilog/coms.v(130[12] 305[6])
    defparam i16354_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1300 (.I0(\data_out_frame[16] [3]), .I1(n57606), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4903));
    defparam i1_2_lut_adj_1300.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1301 (.I0(\data_out_frame[21] [3]), .I1(n26272), 
            .I2(n57317), .I3(n6_adj_4903), .O(n51617));
    defparam i4_4_lut_adj_1301.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1302 (.I0(\data_out_frame[16] [6]), .I1(n57674), 
            .I2(n57137), .I3(\data_out_frame[16] [7]), .O(n14_adj_4904));
    defparam i6_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_137_i2_4_lut (.I0(\data_out_frame[17] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4905));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_137_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1303 (.I0(\data_out_frame[13] [0]), .I1(\data_out_frame[10] [6]), 
            .I2(\data_out_frame[8] [5]), .I3(\data_out_frame[8] [4]), .O(n6_adj_4816));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1303.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_136_i2_4_lut (.I0(\data_out_frame[17] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4906));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_136_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16353_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [5]), 
            .I3(\data_in[2] [5]), .O(n30361));   // verilog/coms.v(130[12] 305[6])
    defparam i16353_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_777_Select_135_i2_4_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4907));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_135_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1304 (.I0(\data_in_frame[12] [5]), .I1(n26031), 
            .I2(n57068), .I3(n26482), .O(n57534));
    defparam i2_3_lut_4_lut_adj_1304.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1305 (.I0(n28415), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n56157));
    defparam i1_4_lut_4_lut_4_lut_adj_1305.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1306 (.I0(n9_adj_4908), .I1(n14_adj_4904), .I2(n59466), 
            .I3(n68337), .O(n59922));
    defparam i7_4_lut_adj_1306.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_134_i2_4_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4909));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_134_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1307 (.I0(\data_in_frame[12] [5]), .I1(n26031), 
            .I2(\data_in_frame[12] [4]), .I3(n51646), .O(n52653));
    defparam i2_3_lut_4_lut_adj_1307.LUT_INIT = 16'h6996;
    SB_LUT4 i16352_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [6]), 
            .I3(\data_in[2] [6]), .O(n30360));   // verilog/coms.v(130[12] 305[6])
    defparam i16352_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16351_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [7]), 
            .I3(\data_in[2] [7]), .O(n30359));   // verilog/coms.v(130[12] 305[6])
    defparam i16351_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16350_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in[3] [0]), .O(n30358));   // verilog/coms.v(130[12] 305[6])
    defparam i16350_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_777_Select_133_i2_4_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4910));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_133_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1308 (.I0(n28415), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n56163));
    defparam i1_4_lut_4_lut_4_lut_adj_1308.LUT_INIT = 16'hfe10;
    SB_LUT4 select_777_Select_132_i2_4_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4911));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_132_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1309 (.I0(n28415), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n56165));
    defparam i1_4_lut_4_lut_4_lut_adj_1309.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1310 (.I0(n59922), .I1(n51617), .I2(GND_net), 
            .I3(GND_net), .O(n57358));
    defparam i1_2_lut_adj_1310.LUT_INIT = 16'h9999;
    SB_LUT4 i2_4_lut_adj_1311 (.I0(n59521), .I1(\data_out_frame[19] [3]), 
            .I2(\data_out_frame[21] [5]), .I3(n57644), .O(n57428));
    defparam i2_4_lut_adj_1311.LUT_INIT = 16'h6996;
    SB_CARRY add_1099_6 (.CI(n49181), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n49182));
    SB_LUT4 i16349_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in[3] [1]), .O(n30357));   // verilog/coms.v(130[12] 305[6])
    defparam i16349_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16348_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in[3] [2]), .O(n30356));   // verilog/coms.v(130[12] 305[6])
    defparam i16348_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFESS data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4831), .S(n56871));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1312 (.I0(\data_out_frame[19] [3]), .I1(n57771), 
            .I2(n57671), .I3(n26858), .O(n51672));
    defparam i3_4_lut_adj_1312.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1313 (.I0(n51672), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[23] [6]), .I3(\data_out_frame[25] [7]), 
            .O(n10_adj_4912));
    defparam i4_4_lut_adj_1313.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_208_i3_4_lut (.I0(n57359), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n10_adj_4912), .I3(n57428), .O(n3_adj_4913));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_208_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i16347_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in[3] [3]), .O(n30355));   // verilog/coms.v(130[12] 305[6])
    defparam i16347_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_777_Select_131_i2_4_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4914));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_131_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i16346_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in[3] [4]), .O(n30354));   // verilog/coms.v(130[12] 305[6])
    defparam i16346_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFESS data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4829), .S(n56870));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1314 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(\data_in_frame[13] [1]), .I3(GND_net), .O(n26449));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1314.LUT_INIT = 16'h9696;
    SB_LUT4 i16345_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in[3] [5]), .O(n30353));   // verilog/coms.v(130[12] 305[6])
    defparam i16345_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 add_1099_5_lut (.I0(n56736), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n49180), .O(n56740)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1099_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1315 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25] [7]), 
            .I2(neopxl_color[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4915));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1315.LUT_INIT = 16'ha088;
    SB_LUT4 i16344_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in[3] [6]), .O(n30352));   // verilog/coms.v(130[12] 305[6])
    defparam i16344_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16361_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [5]), 
            .I3(\data_in[1] [5]), .O(n30369));   // verilog/coms.v(130[12] 305[6])
    defparam i16361_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_777_Select_130_i2_4_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4916));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_130_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i42280_2_lut_3_lut (.I0(n3470), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n57917));
    defparam i42280_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1316 (.I0(\data_out_frame[15] [4]), .I1(n25696), 
            .I2(n26257), .I3(\data_out_frame[17] [5]), .O(n6_adj_4775));
    defparam i1_2_lut_3_lut_4_lut_adj_1316.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_129_i2_4_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4917));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_129_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_128_i2_4_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4918));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_128_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_105_i2_4_lut (.I0(\data_out_frame[13] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4902));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_105_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [0]), 
            .O(n56754));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h5100;
    SB_LUT4 select_777_Select_206_i2_4_lut (.I0(\data_out_frame[25] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4919));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_206_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1317 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[13] [0]), 
            .I2(setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4901));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1317.LUT_INIT = 16'ha088;
    SB_LUT4 select_777_Select_205_i2_4_lut (.I0(\data_out_frame[25] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4920));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_205_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1318 (.I0(n59212), .I1(n59279), .I2(\data_in_frame[19] [6]), 
            .I3(GND_net), .O(n51684));
    defparam i1_2_lut_3_lut_adj_1318.LUT_INIT = 16'h6969;
    SB_DFFESS data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4811), .S(n56869));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_103_i2_4_lut (.I0(\data_out_frame[12] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4900));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_103_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1319 (.I0(n59212), .I1(n59279), .I2(n59284), 
            .I3(GND_net), .O(n52615));
    defparam i1_2_lut_3_lut_adj_1319.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_102_i2_4_lut (.I0(\data_out_frame[12] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4899));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_102_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4809), .S(n56868));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4806), .S(n56867));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1320 (.I0(n28417), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n56369));
    defparam i1_4_lut_4_lut_4_lut_adj_1320.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1321 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [1]), 
            .O(n56755));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1321.LUT_INIT = 16'h5100;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1322 (.I0(n28417), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n56367));
    defparam i1_4_lut_4_lut_4_lut_adj_1322.LUT_INIT = 16'hfe10;
    SB_LUT4 select_777_Select_204_i2_4_lut (.I0(\data_out_frame[25] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4921));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_204_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_101_i2_4_lut (.I0(\data_out_frame[12] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4898));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_101_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i182 (.Q(\data_in_frame[22] [5]), .C(clk16MHz), 
           .D(n29684));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1099_5 (.CI(n49180), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n49181));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1323 (.I0(n8), .I1(n3470), .I2(n161), 
            .I3(n10), .O(n28409));
    defparam i1_2_lut_3_lut_4_lut_adj_1323.LUT_INIT = 16'hffbf;
    SB_LUT4 select_777_Select_100_i2_4_lut (.I0(\data_out_frame[12] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4897));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_100_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1324 (.I0(n8), .I1(n3470), .I2(n161), 
            .I3(n10_adj_11), .O(n28399));
    defparam i1_2_lut_3_lut_4_lut_adj_1324.LUT_INIT = 16'hffbf;
    SB_LUT4 select_777_Select_58_i2_4_lut (.I0(\data_out_frame[7] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4925));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_58_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1325 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26][2] ), 
            .O(n56756));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1325.LUT_INIT = 16'h5100;
    SB_LUT4 i46695_3_lut_4_lut (.I0(n26335), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[2] [7]), .O(n62366));
    defparam i46695_3_lut_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 select_777_Select_57_i2_4_lut (.I0(\data_out_frame[7] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4926));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_57_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_99_i2_4_lut (.I0(\data_out_frame[12] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4896));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_99_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i7_3_lut_4_lut (.I0(\data_in_frame[1] [7]), .I1(n25797), .I2(\data_in_frame[0] [0]), 
            .I3(Kp_23__N_748), .O(n24_adj_4927));
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h2112;
    SB_LUT4 i1_2_lut_3_lut_adj_1326 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n25797));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_3_lut_adj_1326.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_56_i2_4_lut (.I0(\data_out_frame[7] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4928));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_56_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1327 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[2] [6]), .I3(GND_net), .O(n26652));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_3_lut_adj_1327.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_127_i2_4_lut (.I0(\data_out_frame[15] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4929));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_127_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_98_i2_4_lut (.I0(\data_out_frame[12] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4895));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_98_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1328 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [3]), 
            .O(n56752));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1328.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_3_lut_adj_1329 (.I0(\data_in_frame[21] [7]), .I1(\data_in_frame[21] [6]), 
            .I2(n51684), .I3(GND_net), .O(n57519));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1329.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_97_i2_4_lut (.I0(\data_out_frame[12] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4894));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_97_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 add_1099_4_lut (.I0(n56736), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(n49179), .O(n56739)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1099_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1330 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [4]), 
            .O(n56757));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1330.LUT_INIT = 16'h5100;
    SB_DFFE data_in_frame_0___i16 (.Q(\data_in_frame[1] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29889));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i183 (.Q(\data_in_frame[22] [6]), .C(clk16MHz), 
           .D(n29687));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1331 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [5]), 
            .O(n56750));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1331.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1332 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [6]), 
            .O(n56758));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1332.LUT_INIT = 16'h5100;
    SB_CARRY add_1099_4 (.CI(n49179), .I0(\byte_transmit_counter[2] ), .I1(GND_net), 
            .CO(n49180));
    SB_LUT4 add_1099_3_lut (.I0(n56736), .I1(\byte_transmit_counter[1] ), 
            .I2(GND_net), .I3(n49178), .O(n56738)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1099_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1333 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [7]), 
            .O(n56759));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1333.LUT_INIT = 16'h5100;
    SB_LUT4 select_777_Select_96_i2_4_lut (.I0(\data_out_frame[12] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4893));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_96_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_95_i2_4_lut (.I0(\data_out_frame[11] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4892));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_95_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1334 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [0]), 
            .O(n56760));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1334.LUT_INIT = 16'h5100;
    SB_LUT4 i1_4_lut_adj_1335 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[11] [6]), 
            .I2(encoder1_position_scaled[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4891));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1335.LUT_INIT = 16'ha088;
    SB_DFFE data_in_frame_0___i15 (.Q(\data_in_frame[1] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29885));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i14 (.Q(\data_in_frame[1] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29881));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i13 (.Q(\data_in_frame[1] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29878));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4930), .S(n56866));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1099_3 (.CI(n49178), .I0(\byte_transmit_counter[1] ), .I1(GND_net), 
            .CO(n49179));
    SB_LUT4 select_777_Select_93_i2_4_lut (.I0(\data_out_frame[11] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4890));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_93_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1336 (.I0(n28391), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n56197));
    defparam i1_4_lut_4_lut_4_lut_adj_1336.LUT_INIT = 16'hfe10;
    SB_LUT4 select_777_Select_92_i2_4_lut (.I0(\data_out_frame[11] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4889));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_92_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4931), .S(n56865));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4932), .S(n56864));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_4_lut_4_lut_adj_1337 (.I0(n28391), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[15][6] ), .O(n56153));
    defparam i1_4_lut_4_lut_4_lut_adj_1337.LUT_INIT = 16'hfe10;
    SB_LUT4 select_777_Select_91_i2_4_lut (.I0(\data_out_frame[11] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4888));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_91_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_90_i2_4_lut (.I0(\data_out_frame[11] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4887));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_90_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_126_i2_4_lut (.I0(\data_out_frame[15] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4933));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_126_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_125_i2_4_lut (.I0(\data_out_frame[15] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4934));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_125_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1338 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [1]), 
            .O(n56761));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1338.LUT_INIT = 16'h5100;
    SB_LUT4 select_777_Select_124_i2_4_lut (.I0(\data_out_frame[15] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4935));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_124_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1339 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27][2] ), 
            .O(n56762));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1339.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1340 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [3]), 
            .O(n56753));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1340.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1341 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [4]), 
            .O(n56749));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1341.LUT_INIT = 16'h5100;
    SB_DFF data_in_frame_0___i184 (.Q(\data_in_frame[22] [7]), .C(clk16MHz), 
           .D(n56027));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4936), .S(n56863));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i12 (.Q(\data_in_frame[1] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29874));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4937), .S(n56862));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4938), .S(n56861));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4939), .S(n56860));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1342 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n57041), .O(n59242));   // verilog/coms.v(156[9:50])
    defparam i2_3_lut_4_lut_adj_1342.LUT_INIT = 16'hffbf;
    SB_DFFESS data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4940), .S(n56859));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4941), .S(n56858));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk16MHz), 
            .E(n30585), .D(n2_adj_4942), .S(n29030));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4943), .S(n56857));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1343 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [5]), 
            .O(n56751));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1343.LUT_INIT = 16'h5100;
    SB_DFFESS data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4944), .S(n56856));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4945), .S(n56855));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i185 (.Q(\data_in_frame[23] [0]), .C(clk16MHz), 
           .D(n29699));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i11 (.Q(\data_in_frame[1] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29870));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i10 (.Q(\data_in_frame[1] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29867));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1344 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [6]), 
            .O(n56763));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1344.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1345 (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [7]), 
            .O(n56764));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1345.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1346 (.I0(n40970), .I1(n57917), .I2(n7_adj_4946), 
            .I3(\FRAME_MATCHER.i [0]), .O(n28387));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_4_lut_adj_1346.LUT_INIT = 16'hf7ff;
    SB_DFF data_in_frame_0___i4 (.Q(\data_in_frame[0] [3]), .C(clk16MHz), 
           .D(n29713));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 equal_310_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i[5] ), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(GND_net), .O(n10));   // verilog/coms.v(158[12:15])
    defparam equal_310_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 select_777_Select_89_i2_4_lut (.I0(\data_out_frame[11] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4879));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_89_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i186 (.Q(\data_in_frame[23] [1]), .C(clk16MHz), 
           .D(n29728));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_88_i2_4_lut (.I0(\data_out_frame[11] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4878));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_88_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 equal_302_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i[5] ), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(GND_net), .O(n10_adj_11));   // verilog/coms.v(158[12:15])
    defparam equal_302_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 select_777_Select_87_i2_4_lut (.I0(\data_out_frame[10] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4877));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_87_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_86_i2_4_lut (.I0(\data_out_frame[10] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4876));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_86_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 add_1099_2_lut (.I0(n56736), .I1(\byte_transmit_counter[0] ), 
            .I2(tx_transmit_N_3416), .I3(GND_net), .O(n56744)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1099_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 select_777_Select_85_i2_4_lut (.I0(\data_out_frame[10] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4875));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_85_i2_4_lut.LUT_INIT = 16'hc088;
    SB_CARRY add_1099_2 (.CI(GND_net), .I0(\byte_transmit_counter[0] ), 
            .I1(tx_transmit_N_3416), .CO(n49178));
    SB_DFF data_in_frame_0___i187 (.Q(\data_in_frame[23] [2]), .C(clk16MHz), 
           .D(n29737));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_84_i2_4_lut (.I0(\data_out_frame[10] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4874));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_84_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i188 (.Q(\data_in_frame[23] [3]), .C(clk16MHz), 
           .D(n29740));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i5 (.Q(\data_in_frame[0] [4]), .C(clk16MHz), 
           .D(n56361));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_83_i2_4_lut (.I0(\data_out_frame[10] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4873));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_83_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_82_i2_4_lut (.I0(\data_out_frame[10] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4872));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_82_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_81_i2_4_lut (.I0(\data_out_frame[10] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4871));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_81_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_80_i2_4_lut (.I0(\data_out_frame[10] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4870));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_80_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i23225_3_lut (.I0(n376), .I1(n456), .I2(n11610), .I3(GND_net), 
            .O(n27692));
    defparam i23225_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0___i6 (.Q(\data_in_frame[0] [5]), .C(clk16MHz), 
           .D(n56369));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i7 (.Q(\data_in_frame[0] [6]), .C(clk16MHz), 
           .D(n56367));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_79_i2_4_lut (.I0(\data_out_frame[9] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4869));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_79_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i189 (.Q(\data_in_frame[23] [4]), .C(clk16MHz), 
           .D(n29756));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_78_i2_4_lut (.I0(\data_out_frame[9] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4868));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_78_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_77_i2_4_lut (.I0(\data_out_frame[9] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4867));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_77_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_76_i2_4_lut (.I0(\data_out_frame[9] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4866));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_76_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_75_i2_4_lut (.I0(\data_out_frame[9] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4865));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_75_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_74_i2_4_lut (.I0(\data_out_frame[9] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4864));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_74_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i190 (.Q(\data_in_frame[23] [5]), .C(clk16MHz), 
           .D(n29759));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i8 (.Q(\data_in_frame[0] [7]), .C(clk16MHz), 
           .D(n29762));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_73_i2_4_lut (.I0(\data_out_frame[9] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4848));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_73_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFE data_in_frame_0___i9 (.Q(\data_in_frame[1] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29853));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i191 (.Q(\data_in_frame[23] [6]), .C(clk16MHz), 
           .D(n29765));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i192 (.Q(\data_in_frame[23] [7]), .C(clk16MHz), 
           .D(n29768));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i1 (.Q(deadband[1]), .C(clk16MHz), .D(n29850), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i2 (.Q(deadband[2]), .C(clk16MHz), .D(n29849), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i3 (.Q(deadband[3]), .C(clk16MHz), .D(n29848), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i4 (.Q(deadband[4]), .C(clk16MHz), .D(n29847), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i5 (.Q(deadband[5]), .C(clk16MHz), .D(n29846), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i6 (.Q(deadband[6]), .C(clk16MHz), .D(n29845), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i7 (.Q(deadband[7]), .C(clk16MHz), .D(n29844), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i8 (.Q(deadband[8]), .C(clk16MHz), .D(n29843), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i9 (.Q(deadband[9]), .C(clk16MHz), .D(n29842), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i10 (.Q(deadband[10]), .C(clk16MHz), .D(n29841), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i11 (.Q(deadband[11]), .C(clk16MHz), .D(n29840), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i12 (.Q(deadband[12]), .C(clk16MHz), .D(n29839), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i13 (.Q(deadband[13]), .C(clk16MHz), .D(n29838), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i14 (.Q(deadband[14]), .C(clk16MHz), .D(n29837), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i15 (.Q(deadband[15]), .C(clk16MHz), .D(n29836), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i16 (.Q(deadband[16]), .C(clk16MHz), .D(n29835), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i17 (.Q(deadband[17]), .C(clk16MHz), .D(n29834), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i18 (.Q(deadband[18]), .C(clk16MHz), .D(n29833), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i19 (.Q(deadband[19]), .C(clk16MHz), .D(n29832), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i20 (.Q(deadband[20]), .C(clk16MHz), .D(n29831), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i21 (.Q(deadband[21]), .C(clk16MHz), .D(n29830), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i22 (.Q(deadband[22]), .C(clk16MHz), .D(n29829), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i23 (.Q(deadband[23]), .C(clk16MHz), .D(n29828), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk16MHz), .D(n29827), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk16MHz), .D(n29826), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk16MHz), .D(n29825), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk16MHz), .D(n29824), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk16MHz), .D(n29823), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk16MHz), .D(n29822), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk16MHz), .D(n29821), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk16MHz), .D(n29820), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk16MHz), .D(n29819), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk16MHz), .D(n29818), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk16MHz), .D(n29817), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk16MHz), .D(n29816), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk16MHz), .D(n29815), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk16MHz), .D(n29814), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk16MHz), .D(n29813), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk16MHz), .D(n29812), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1347 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[9] [0]), 
            .I2(encoder1_position_scaled[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4847));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1347.LUT_INIT = 16'ha088;
    SB_DFFR IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk16MHz), .D(n29811), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk16MHz), .D(n29810), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk16MHz), .D(n29809), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk16MHz), .D(n29808), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_71_i2_4_lut (.I0(\data_out_frame[8] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4845));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_71_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFR IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk16MHz), .D(n29807), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk16MHz), .D(n29806), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk16MHz), .D(n29805), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i1 (.Q(\Kp[1] ), .C(clk16MHz), .D(n29804), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i2 (.Q(\Kp[2] ), .C(clk16MHz), .D(n29803), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i3 (.Q(\Kp[3] ), .C(clk16MHz), .D(n29802), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13_2_lut (.I0(pwm_setpoint[22]), .I1(\pwm_counter[22] ), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/pwm.v(11[19:30])
    defparam i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15_2_lut (.I0(pwm_setpoint[21]), .I1(\pwm_counter[21] ), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/pwm.v(11[19:30])
    defparam i15_2_lut.LUT_INIT = 16'h6666;
    SB_DFFR Kp_i4 (.Q(\Kp[4] ), .C(clk16MHz), .D(n29801), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i5 (.Q(\Kp[5] ), .C(clk16MHz), .D(n29800), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i6 (.Q(\Kp[6] ), .C(clk16MHz), .D(n29799), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i7 (.Q(\Kp[7] ), .C(clk16MHz), .D(n29798), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i8 (.Q(\Kp[8] ), .C(clk16MHz), .D(n29797), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i9 (.Q(\Kp[9] ), .C(clk16MHz), .D(n29796), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i10 (.Q(\Kp[10] ), .C(clk16MHz), .D(n29795), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i11 (.Q(\Kp[11] ), .C(clk16MHz), .D(n29794), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i12 (.Q(\Kp[12] ), .C(clk16MHz), .D(n29793), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i13 (.Q(\Kp[13] ), .C(clk16MHz), .D(n29792), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i14 (.Q(\Kp[14] ), .C(clk16MHz), .D(n29791), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i15 (.Q(\Kp[15] ), .C(clk16MHz), .D(n29790), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i1 (.Q(\Ki[1] ), .C(clk16MHz), .D(n29789), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i2 (.Q(\Ki[2] ), .C(clk16MHz), .D(n29788), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i3 (.Q(\Ki[3] ), .C(clk16MHz), .D(n29787), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i4 (.Q(\Ki[4] ), .C(clk16MHz), .D(n29786), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i5 (.Q(\Ki[5] ), .C(clk16MHz), .D(n29785), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i6 (.Q(\Ki[6] ), .C(clk16MHz), .D(n29784), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i7 (.Q(\Ki[7] ), .C(clk16MHz), .D(n29783), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i8 (.Q(\Ki[8] ), .C(clk16MHz), .D(n29782), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i9 (.Q(\Ki[9] ), .C(clk16MHz), .D(n29781), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i10 (.Q(\Ki[10] ), .C(clk16MHz), .D(n29780), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i11 (.Q(\Ki[11] ), .C(clk16MHz), .D(n29779), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i12 (.Q(\Ki[12] ), .C(clk16MHz), .D(n29778), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i13 (.Q(\Ki[13] ), .C(clk16MHz), .D(n29777), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i14 (.Q(\Ki[14] ), .C(clk16MHz), .D(n29776), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i15 (.Q(\Ki[15] ), .C(clk16MHz), .D(n29775), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4935), .S(n56854));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4934), .S(n56853));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4933), .S(n56852));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4929), .S(n56851));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4918), .S(n56850));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4917), .S(n56849));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4916), .S(n56775));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4914), .S(n56777));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1348 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(n3470), .I3(n43293), .O(n145));
    defparam i4_4_lut_adj_1348.LUT_INIT = 16'h1000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1349 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n57041), .O(n57044));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1349.LUT_INIT = 16'hfffd;
    SB_DFFESS data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4911), .S(n56778));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4910), .S(n56779));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4909), .S(n56780));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4907), .S(n56781));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4906), .S(n56783));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4905), .S(n56784));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4886), .S(n56785));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4880), .S(n56786));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4862), .S(n56787));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4861), .S(n56788));   // verilog/coms.v(130[12] 305[6])
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_4012  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk16MHz), .D(n29746));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4860), .S(n56789));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4859), .S(n56790));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4856), .S(n56791));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4854), .S(n56792));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk16MHz), .D(n29736));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4851), .S(n56793));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4844), .S(n56774));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4838), .S(n56794));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4837), .S(n56795));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4836), .S(n56796));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i7 (.Q(current_limit[7]), .C(clk16MHz), .D(n29735));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk16MHz), .D(n29734));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk16MHz), .D(n29733));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk16MHz), .D(n29732));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk16MHz), .D(n29731));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4827), .S(n56797));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4825), .S(n56798));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk16MHz), .D(n29727));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk16MHz), .D(n29726));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk16MHz), .D(n29725));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk16MHz), .D(n29723));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk16MHz), .D(n29722));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk16MHz), .D(n29721));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk16MHz), .D(n29720));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk16MHz), .D(n29719));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk16MHz), .D(n29718));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i8 (.Q(current_limit[8]), .C(clk16MHz), .D(n29717));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4805), .S(n56799));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4804), .S(n56800));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i9 (.Q(current_limit[9]), .C(clk16MHz), .D(n29716));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i10 (.Q(current_limit[10]), .C(clk16MHz), .D(n29712));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk16MHz), .D(n29711));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4802), .S(n56801));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4801), .S(n56802));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i11 (.Q(current_limit[11]), .C(clk16MHz), .D(n29708));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i12 (.Q(current_limit[12]), .C(clk16MHz), .D(n29707));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4800), .S(n56803));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i13 (.Q(current_limit[13]), .C(clk16MHz), .D(n29706));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i14 (.Q(current_limit[14]), .C(clk16MHz), .D(n29705));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk16MHz), .D(n29703));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk16MHz), .D(n29702));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk16MHz), .D(n29698));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk16MHz), .D(n29694));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1350 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n40973), .O(n28438));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1350.LUT_INIT = 16'h0200;
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk16MHz), .D(n29693));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk16MHz), .D(n29692));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk16MHz), .D(n29691));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1351 (.I0(\FRAME_MATCHER.i [0]), .I1(n3470), .I2(GND_net), 
            .I3(GND_net), .O(n57016));
    defparam i1_2_lut_adj_1351.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_4_lut_adj_1352 (.I0(n25991), .I1(\data_in_frame[19]_c [7]), 
            .I2(\data_in_frame[16] [3]), .I3(\data_in_frame[20] [5]), .O(n62126));
    defparam i1_4_lut_adj_1352.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1353 (.I0(n52651), .I1(n57463), .I2(n62128), 
            .I3(n62126), .O(n62134));
    defparam i1_4_lut_adj_1353.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1354 (.I0(n52695), .I1(n57497), .I2(n59162), 
            .I3(n62134), .O(n62140));
    defparam i1_4_lut_adj_1354.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1355 (.I0(n57389), .I1(n51684), .I2(n62140), 
            .I3(n57494), .O(n62146));
    defparam i1_4_lut_adj_1355.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_55_i2_4_lut (.I0(\data_out_frame[6] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4947));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_55_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1356 (.I0(n23898), .I1(n57371), .I2(n62146), 
            .I3(n52615), .O(n62152));
    defparam i1_4_lut_adj_1356.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1357 (.I0(n57372), .I1(n57783), .I2(n57168), 
            .I3(n62152), .O(n57292));
    defparam i1_4_lut_adj_1357.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1358 (.I0(\data_in_frame[15][6] ), .I1(\data_in_frame[13] [4]), 
            .I2(Kp_23__N_1301), .I3(n25987), .O(n57635));
    defparam i3_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1359 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n57037), .O(n57039));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1359.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_4_lut_adj_1360 (.I0(n25128), .I1(n52594), .I2(n62014), 
            .I3(n57433), .O(n62018));
    defparam i1_4_lut_adj_1360.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1361 (.I0(n52337), .I1(n59955), .I2(n62018), 
            .I3(n51926), .O(n57476));
    defparam i1_4_lut_adj_1361.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1362 (.I0(\data_in_frame[16] [6]), .I1(\data_in_frame[15][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n62036));
    defparam i1_2_lut_adj_1362.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1363 (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[15][4] ), 
            .I2(\data_in_frame[13] [0]), .I3(\data_in_frame[16]_c [0]), 
            .O(n62042));
    defparam i1_4_lut_adj_1363.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1364 (.I0(n62042), .I1(Kp_23__N_1389), .I2(n62036), 
            .I3(\data_in_frame[10] [6]), .O(n62046));
    defparam i1_4_lut_adj_1364.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1365 (.I0(n57774), .I1(Kp_23__N_1067), .I2(n62046), 
            .I3(n57780), .O(n62052));
    defparam i1_4_lut_adj_1365.LUT_INIT = 16'h6996;
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk16MHz), .D(n29673));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk16MHz), .D(n29672));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i15 (.Q(current_limit[15]), .C(clk16MHz), .D(n29662));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk16MHz), .D(n29650));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk16MHz), .D(n29644), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk16MHz), .D(n29640), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i0 (.Q(current_limit[0]), .C(clk16MHz), .D(n29639));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk16MHz), .D(n29638));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk16MHz), .D(n29637));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i0 (.Q(\Ki[0] ), .C(clk16MHz), .D(n29636), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i0 (.Q(\Kp[0] ), .C(clk16MHz), .D(n29635), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk16MHz), .D(n29613), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1366 (.I0(n57686), .I1(n57143), .I2(n57355), 
            .I3(n62052), .O(n62058));
    defparam i1_4_lut_adj_1366.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4762), .S(n56804));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1367 (.I0(n52825), .I1(n52651), .I2(n59802), 
            .I3(n62058), .O(n62064));
    defparam i1_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1368 (.I0(n52615), .I1(n57479), .I2(n52637), 
            .I3(n62064), .O(n52337));
    defparam i1_4_lut_adj_1368.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4761), .S(n56805));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4760), .S(n56806));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk16MHz), 
            .E(n30647), .D(n2_adj_4759), .S(n28989));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4758), .S(n56807));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk16MHz), 
            .E(n30649), .D(n2_adj_4756), .S(n28987));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4754), .S(n56808));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4753), .S(n56809));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4752), .S(n56810));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4751), .S(n56811));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4750), .S(n56812));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk16MHz), 
            .E(n30655), .D(n2_adj_4749), .S(n28981));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4748), .S(n56813));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4747), .S(n56814));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4746), .S(n56815));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4745), .S(n56816));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4744), .S(n56817));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4743), .S(n56818));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4742), .S(n56819));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4741), .S(n56820));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4740), .S(n56821));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4739), .S(n56822));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4735), .S(n56823));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4733), .S(n56824));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4732), .S(n56825));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1369 (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26406));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1369.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1370 (.I0(\data_in_frame[18] [5]), .I1(n57713), 
            .I2(n25899), .I3(n26406), .O(n57062));
    defparam i3_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut (.I0(n51281), .I1(n57062), .I2(\data_in_frame[18] [0]), 
            .I3(GND_net), .O(n62026));
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_203_i2_4_lut (.I0(\data_out_frame[25] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4948));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_203_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1371 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[25] [2]), 
            .I2(neopxl_color[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4949));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1371.LUT_INIT = 16'ha088;
    SB_DFFR \FRAME_MATCHER.i_1942__i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk16MHz), 
            .D(n28050), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 i1_4_lut_adj_1372 (.I0(n59279), .I1(n52337), .I2(n51588), 
            .I3(n62026), .O(n59955));
    defparam i1_4_lut_adj_1372.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1373 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[18] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n57713));
    defparam i1_2_lut_adj_1373.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1374 (.I0(n57490), .I1(n62160), .I2(\data_in_frame[20] [1]), 
            .I3(\data_in_frame[20] [2]), .O(n62164));
    defparam i1_4_lut_adj_1374.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1375 (.I0(n59279), .I1(n59955), .I2(n51281), 
            .I3(n62164), .O(n57783));
    defparam i1_4_lut_adj_1375.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_201_i2_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4950));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_201_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 equal_293_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [1]), .I3(GND_net), .O(n8_adj_12));   // verilog/coms.v(157[7:23])
    defparam equal_293_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 select_777_Select_200_i2_4_lut (.I0(\data_out_frame[25] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4952));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_200_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4730), .S(n56826));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4729), .S(n56827));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4728), .S(n56828));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4727), .S(n56829));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4726), .S(n56830));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR \FRAME_MATCHER.i_1942__i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk16MHz), 
            .D(n28052), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk16MHz), 
            .D(n28054), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk16MHz), 
            .D(n28056), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk16MHz), 
            .D(n28058), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk16MHz), 
            .D(n28060), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk16MHz), 
            .D(n28062), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk16MHz), 
            .D(n28064), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk16MHz), 
            .D(n28066), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk16MHz), 
            .D(n28068), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk16MHz), 
            .D(n28070), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk16MHz), 
            .D(n28072), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk16MHz), 
            .D(n28074), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk16MHz), 
            .D(n28076), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk16MHz), 
            .D(n28078), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk16MHz), 
            .D(n28080), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk16MHz), 
            .D(n28082), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk16MHz), 
            .D(n28084), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk16MHz), 
            .D(n28086), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk16MHz), 
            .D(n28088), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk16MHz), 
            .D(n28090), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk16MHz), 
            .D(n28092), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFESS data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2), .S(n56831));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR \FRAME_MATCHER.i_1942__i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk16MHz), 
            .D(n28094), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk16MHz), 
            .D(n28096), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk16MHz), 
            .D(n28098), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk16MHz), 
            .D(n28100), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk16MHz), 
            .D(n28102), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i5  (.Q(\FRAME_MATCHER.i[5] ), .C(clk16MHz), 
            .D(n28104), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk16MHz), 
            .D(n28106), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i3  (.Q(\FRAME_MATCHER.i[3] ), .C(clk16MHz), 
            .D(n28108), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk16MHz), 
            .D(n28110), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_1942__i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk16MHz), 
            .D(n28112), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 i1_3_lut_adj_1376 (.I0(n59284), .I1(n59141), .I2(n59212), 
            .I3(GND_net), .O(n57371));
    defparam i1_3_lut_adj_1376.LUT_INIT = 16'h6969;
    SB_LUT4 select_777_Select_199_i2_4_lut (.I0(\data_out_frame[24] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4953));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_199_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1377 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[24] [6]), 
            .I2(neopxl_color[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4954));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1377.LUT_INIT = 16'ha088;
    SB_LUT4 select_777_Select_197_i2_4_lut (.I0(\data_out_frame[24] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4955));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_197_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_196_i2_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4956));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_196_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_33_lut  (.I0(n65365), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [31]), .I3(n50464), .O(n28052)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_33_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_32_lut  (.I0(n65362), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [30]), .I3(n50463), .O(n28054)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_32_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_32  (.CI(n50463), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [30]), .CO(n50464));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_31_lut  (.I0(n65361), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [29]), .I3(n50462), .O(n28056)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_31_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_31  (.CI(n50462), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [29]), .CO(n50463));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_30_lut  (.I0(n65360), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [28]), .I3(n50461), .O(n28058)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_30_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_30  (.CI(n50461), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [28]), .CO(n50462));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_29_lut  (.I0(n65359), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [27]), .I3(n50460), .O(n28060)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_29_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_29  (.CI(n50460), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [27]), .CO(n50461));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_28_lut  (.I0(n65355), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [26]), .I3(n50459), .O(n28062)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_28_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_28  (.CI(n50459), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [26]), .CO(n50460));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_27_lut  (.I0(n65313), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [25]), .I3(n50458), .O(n28064)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_27_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_27  (.CI(n50458), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [25]), .CO(n50459));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_26_lut  (.I0(n65312), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [24]), .I3(n50457), .O(n28066)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_26_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_26  (.CI(n50457), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [24]), .CO(n50458));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_25_lut  (.I0(n65311), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [23]), .I3(n50456), .O(n28068)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_25_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_25  (.CI(n50456), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [23]), .CO(n50457));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_24_lut  (.I0(n65307), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [22]), .I3(n50455), .O(n28070)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_24_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_24  (.CI(n50455), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [22]), .CO(n50456));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_23_lut  (.I0(n65297), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [21]), .I3(n50454), .O(n28072)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_23_lut .LUT_INIT = 16'h8BB8;
    SB_DFFESS data_out_frame_0___i3 (.Q(\data_out_frame[0][2] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4957), .S(n56951));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_23  (.CI(n50454), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [21]), .CO(n50455));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_22_lut  (.I0(n65290), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [20]), .I3(n50453), .O(n28074)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_22_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_22  (.CI(n50453), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [20]), .CO(n50454));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_21_lut  (.I0(n65286), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [19]), .I3(n50452), .O(n28076)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_21_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_21  (.CI(n50452), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [19]), .CO(n50453));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_20_lut  (.I0(n65284), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [18]), .I3(n50451), .O(n28078)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_20_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_20  (.CI(n50451), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [18]), .CO(n50452));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_19_lut  (.I0(n65282), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [17]), .I3(n50450), .O(n28080)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_19_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_19  (.CI(n50450), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [17]), .CO(n50451));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_18_lut  (.I0(n65279), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [16]), .I3(n50449), .O(n28082)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_18_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_18  (.CI(n50449), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [16]), .CO(n50450));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_17_lut  (.I0(n65277), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [15]), .I3(n50448), .O(n28084)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_17_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_17  (.CI(n50448), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [15]), .CO(n50449));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_16_lut  (.I0(n65276), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [14]), .I3(n50447), .O(n28086)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_16_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_16  (.CI(n50447), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [14]), .CO(n50448));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_15_lut  (.I0(n65275), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [13]), .I3(n50446), .O(n28088)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_15_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_15  (.CI(n50446), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [13]), .CO(n50447));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_14_lut  (.I0(n65268), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [12]), .I3(n50445), .O(n28090)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_14_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_14  (.CI(n50445), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [12]), .CO(n50446));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_13_lut  (.I0(n65267), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [11]), .I3(n50444), .O(n28092)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_13_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_13  (.CI(n50444), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [11]), .CO(n50445));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_12_lut  (.I0(n65266), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [10]), .I3(n50443), .O(n28094)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_12_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_12  (.CI(n50443), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [10]), .CO(n50444));
    SB_LUT4 i1_3_lut_adj_1378 (.I0(n59141), .I1(n59980), .I2(\data_in_frame[21] [5]), 
            .I3(GND_net), .O(n57238));
    defparam i1_3_lut_adj_1378.LUT_INIT = 16'h9696;
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_11_lut  (.I0(n65265), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [9]), .I3(n50442), .O(n28096)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_11_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_11  (.CI(n50442), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [9]), .CO(n50443));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_10_lut  (.I0(n65264), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [8]), .I3(n50441), .O(n28098)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_10_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_10  (.CI(n50441), .I0(n28374), 
            .I1(\FRAME_MATCHER.i [8]), .CO(n50442));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_9_lut  (.I0(n65263), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [7]), .I3(n50440), .O(n28100)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_9_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_9  (.CI(n50440), .I0(n28374), .I1(\FRAME_MATCHER.i [7]), 
            .CO(n50441));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_8_lut  (.I0(n65262), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [6]), .I3(n50439), .O(n28102)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_8_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_8  (.CI(n50439), .I0(n28374), .I1(\FRAME_MATCHER.i [6]), 
            .CO(n50440));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_7_lut  (.I0(n65261), .I1(n28374), 
            .I2(\FRAME_MATCHER.i[5] ), .I3(n50438), .O(n28104)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_7_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_7  (.CI(n50438), .I0(n28374), .I1(\FRAME_MATCHER.i[5] ), 
            .CO(n50439));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_6_lut  (.I0(n65260), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [4]), .I3(n50437), .O(n28106)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_6_lut .LUT_INIT = 16'h8BB8;
    SB_DFFESS data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4958), .S(n56950));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_6  (.CI(n50437), .I0(n28374), .I1(\FRAME_MATCHER.i [4]), 
            .CO(n50438));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_5_lut  (.I0(n65259), .I1(n28374), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(n50436), .O(n28108)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_5_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_5  (.CI(n50436), .I0(n28374), .I1(\FRAME_MATCHER.i[3] ), 
            .CO(n50437));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_4_lut  (.I0(n65258), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n50435), .O(n28110)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_4_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_4  (.CI(n50435), .I0(n28374), .I1(\FRAME_MATCHER.i [2]), 
            .CO(n50436));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_3_lut  (.I0(n65257), .I1(n28374), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n50434), .O(n28112)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_3_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_3  (.CI(n50434), .I0(n28374), .I1(\FRAME_MATCHER.i [1]), 
            .CO(n50435));
    SB_LUT4 \FRAME_MATCHER.i_1942_add_4_2_lut  (.I0(GND_net), .I1(n161), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_1942_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \FRAME_MATCHER.i_1942_add_4_2  (.CI(GND_net), .I0(n161), .I1(\FRAME_MATCHER.i [0]), 
            .CO(n50434));
    SB_DFFESS data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4959), .S(n56949));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i9 (.Q(\data_out_frame[1][0] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4960), .S(n56948));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1379 (.I0(\data_in_frame[17] [1]), .I1(n52406), 
            .I2(GND_net), .I3(GND_net), .O(n57479));
    defparam i1_2_lut_adj_1379.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1380 (.I0(\data_in_frame[16][7] ), .I1(n57479), 
            .I2(\data_in_frame[19][3] ), .I3(n57717), .O(n59980));
    defparam i1_4_lut_adj_1380.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1381 (.I0(n59980), .I1(n57128), .I2(GND_net), 
            .I3(GND_net), .O(n23898));
    defparam i1_2_lut_adj_1381.LUT_INIT = 16'h9999;
    SB_DFFESS data_out_frame_0___i10 (.Q(\data_out_frame[1][1] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4961), .S(n56947));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i12 (.Q(\data_out_frame[1][3] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4962), .S(n56946));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i14 (.Q(\data_out_frame[1][5] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4963), .S(n56945));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_adj_1382 (.I0(\data_in_frame[15][1] ), .I1(\data_in_frame[14] [6]), 
            .I2(\data_in_frame[17] [2]), .I3(GND_net), .O(n62098));
    defparam i1_3_lut_adj_1382.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1383 (.I0(n57512), .I1(n25864), .I2(n57720), 
            .I3(n62098), .O(n62104));
    defparam i1_4_lut_adj_1383.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1384 (.I0(n57723), .I1(n52705), .I2(n57698), 
            .I3(n25987), .O(n62090));
    defparam i1_4_lut_adj_1384.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i15 (.Q(\data_out_frame[1][6] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4964), .S(n56944));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1385 (.I0(n52626), .I1(n62090), .I2(n62104), 
            .I3(n51755), .O(n52406));
    defparam i1_4_lut_adj_1385.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1386 (.I0(n59284), .I1(n52406), .I2(\data_in_frame[19][4] ), 
            .I3(GND_net), .O(n59141));
    defparam i1_3_lut_adj_1386.LUT_INIT = 16'h6969;
    SB_DFFESS data_out_frame_0___i16 (.Q(\data_out_frame[1][7] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4965), .S(n56943));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i26 (.Q(\data_out_frame[3][1] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4966), .S(n56942));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1387 (.I0(\data_in_frame[21] [3]), .I1(\data_in_frame[21] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n57223));
    defparam i1_2_lut_adj_1387.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1388 (.I0(\data_in_frame[15] [5]), .I1(n57401), 
            .I2(GND_net), .I3(GND_net), .O(n52695));
    defparam i1_2_lut_adj_1388.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1389 (.I0(n51720), .I1(n57442), .I2(n25938), 
            .I3(\data_in_frame[13] [2]), .O(n57698));
    defparam i3_4_lut_adj_1389.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1390 (.I0(n57698), .I1(\data_in_frame[15][3] ), 
            .I2(\data_in_frame[13] [1]), .I3(GND_net), .O(n59802));
    defparam i2_3_lut_adj_1390.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1391 (.I0(n59802), .I1(n60027), .I2(\data_in_frame[17] [5]), 
            .I3(GND_net), .O(n59279));
    defparam i1_3_lut_adj_1391.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1392 (.I0(\data_in_frame[15][3] ), .I1(n52572), 
            .I2(\data_in_frame[17] [4]), .I3(GND_net), .O(n59212));
    defparam i1_3_lut_adj_1392.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1393 (.I0(n51706), .I1(n58909), .I2(n25971), 
            .I3(\data_in_frame[14] [7]), .O(n51755));
    defparam i1_4_lut_adj_1393.LUT_INIT = 16'h9669;
    SB_DFFS PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk16MHz), .D(n30519), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk16MHz), .D(n30518), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk16MHz), .D(n30517), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i117 (.Q(\data_in_frame[14] [4]), .C(clk16MHz), 
           .D(n29441));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk16MHz), .D(n30515), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk16MHz), .D(n30514), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk16MHz), .D(n30513), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk16MHz), .D(n30512), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i118 (.Q(\data_in_frame[14] [5]), .C(clk16MHz), 
           .D(n29444));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i1 (.Q(\data_in_frame[0] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30503));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i119 (.Q(\data_in_frame[14] [6]), .C(clk16MHz), 
           .D(n29447));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i120 (.Q(\data_in_frame[14] [7]), .C(clk16MHz), 
           .D(n29450));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i116 (.Q(\data_in_frame[14] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n30482));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i121 (.Q(\data_in_frame[15][0] ), .C(clk16MHz), 
           .D(n29453));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i122 (.Q(\data_in_frame[15][1] ), .C(clk16MHz), 
           .D(n29456));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i123 (.Q(\data_in_frame[15][2] ), .C(clk16MHz), 
           .D(n29459));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i115 (.Q(\data_in_frame[14] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n30476));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i124 (.Q(\data_in_frame[15][3] ), .C(clk16MHz), 
           .D(n29462));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i114 (.Q(\data_in_frame[14] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n30472));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i125 (.Q(\data_in_frame[15][4] ), .C(clk16MHz), 
           .D(n29465));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk16MHz), .D(n30470), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i126 (.Q(\data_in_frame[15] [5]), .C(clk16MHz), 
           .D(n56197));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk16MHz), .D(n30468), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk16MHz), .D(n30467));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk16MHz), .D(n30466), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk16MHz), .D(n30465), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk16MHz), .D(n30464), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i127 (.Q(\data_in_frame[15][6] ), .C(clk16MHz), 
           .D(n56153));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk16MHz), .D(n30444), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk16MHz), .D(n30420), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk16MHz), .D(n30398), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i128 (.Q(\data_in_frame[15][7] ), .C(clk16MHz), 
           .D(n29474));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk16MHz), .D(n30396), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk16MHz), .D(n30395), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk16MHz), .D(n30384), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk16MHz), .D(n30382));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk16MHz), .D(n30381));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk16MHz), .D(n30380));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk16MHz), .D(n30379));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk16MHz), .D(n30378));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk16MHz), .D(n30377));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk16MHz), .D(n30376));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk16MHz), .D(n30375));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk16MHz), .D(n30374));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk16MHz), .D(n30373));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i28 (.Q(\data_out_frame[3][3] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4967), .S(n56941));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1394 (.I0(\data_in_frame[12] [6]), .I1(n26031), 
            .I2(GND_net), .I3(GND_net), .O(n57512));
    defparam i1_2_lut_adj_1394.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk16MHz), .D(n30372));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk16MHz), .D(n30371));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk16MHz), .D(n30370));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk16MHz), .D(n30369));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk16MHz), .D(n30368));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk16MHz), .D(n30367));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk16MHz), .D(n30366));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk16MHz), .D(n30365));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1395 (.I0(n25952), .I1(n25971), .I2(\data_in_frame[13] [5]), 
            .I3(GND_net), .O(n25987));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1395.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk16MHz), .D(n30364));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk16MHz), .D(n30363));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk16MHz), .D(n30362));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1396 (.I0(n25987), .I1(\data_in_frame[15][1] ), 
            .I2(GND_net), .I3(GND_net), .O(n57355));
    defparam i1_2_lut_adj_1396.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk16MHz), .D(n30361));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1397 (.I0(n57774), .I1(n57683), .I2(n25853), 
            .I3(n57068), .O(n52572));
    defparam i1_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk16MHz), .D(n30360));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk16MHz), .D(n30359));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk16MHz), .D(n30358));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk16MHz), .D(n30357));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk16MHz), .D(n30356));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk16MHz), .D(n30355));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk16MHz), .D(n30354));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i29 (.Q(\data_out_frame[3][4] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4968), .S(n56940));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk16MHz), .D(n30353));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk16MHz), .D(n30352));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk16MHz), .D(n30351));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_adj_1398 (.I0(n52572), .I1(n57355), .I2(\data_in_frame[17] [3]), 
            .I3(GND_net), .O(n62174));
    defparam i1_3_lut_adj_1398.LUT_INIT = 16'h9696;
    SB_DFFR PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk16MHz), .D(n30350), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk16MHz), .D(n30349), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk16MHz), .D(n30348));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk16MHz), .D(n30347), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_195_i2_4_lut (.I0(\data_out_frame[24] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4969));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_195_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i41 (.Q(\data_in_frame[5] [0]), .C(clk16MHz), 
           .D(n29973));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_194_i2_4_lut (.I0(\data_out_frame[24] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4970));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_194_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFF data_in_frame_0___i129 (.Q(\data_in_frame[16]_c [0]), .C(clk16MHz), 
           .D(n56177));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i42 (.Q(\data_in_frame[5] [1]), .C(clk16MHz), 
           .D(n29976));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk16MHz), .D(n30343), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i43 (.Q(\data_in_frame[5] [2]), .C(clk16MHz), 
           .D(n29979));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i44 (.Q(\data_in_frame[5] [3]), .C(clk16MHz), 
           .D(n29982));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1399 (.I0(n57401), .I1(n51755), .I2(n52825), 
            .I3(n62174), .O(n59284));
    defparam i1_4_lut_adj_1399.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0___i130 (.Q(\data_in_frame[16][1] ), .C(clk16MHz), 
           .D(n56201));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i1 (.Q(current_limit[1]), .C(clk16MHz), .D(n30339));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i131 (.Q(\data_in_frame[16][2] ), .C(clk16MHz), 
           .D(n56199));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i132 (.Q(\data_in_frame[16] [3]), .C(clk16MHz), 
           .D(n29490));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i133 (.Q(\data_in_frame[16] [4]), .C(clk16MHz), 
           .D(n29493));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i134 (.Q(\data_in_frame[16] [5]), .C(clk16MHz), 
           .D(n29496));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i135 (.Q(\data_in_frame[16] [6]), .C(clk16MHz), 
           .D(n29499));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i136 (.Q(\data_in_frame[16][7] ), .C(clk16MHz), 
           .D(n56249));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i137 (.Q(\data_in_frame[17] [0]), .C(clk16MHz), 
           .D(n56107));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i138 (.Q(\data_in_frame[17] [1]), .C(clk16MHz), 
           .D(n56103));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i139 (.Q(\data_in_frame[17] [2]), .C(clk16MHz), 
           .D(n56101));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i140 (.Q(\data_in_frame[17] [3]), .C(clk16MHz), 
           .D(n56099));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i141 (.Q(\data_in_frame[17] [4]), .C(clk16MHz), 
           .D(n56095));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i142 (.Q(\data_in_frame[17] [5]), .C(clk16MHz), 
           .D(n56091));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i31 (.Q(\data_out_frame[3][6] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4971), .S(n56771));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i45 (.Q(\data_in_frame[5] [4]), .C(clk16MHz), 
           .D(n29986));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i46 (.Q(\data_in_frame[5] [5]), .C(clk16MHz), 
           .D(n29989));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i47 (.Q(\data_in_frame[5] [6]), .C(clk16MHz), 
           .D(n29992));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i113 (.Q(\data_in_frame[14] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n30312));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i143 (.Q(\data_in_frame[17] [6]), .C(clk16MHz), 
           .D(n56087));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i144 (.Q(\data_in_frame[17] [7]), .C(clk16MHz), 
           .D(n56083));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i145 (.Q(\data_in_frame[18] [0]), .C(clk16MHz), 
           .D(n56079));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i112 (.Q(\data_in_frame[13] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n30305));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i48 (.Q(\data_in_frame[5] [7]), .C(clk16MHz), 
           .D(n29995));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i49 (.Q(\data_in_frame[6][0] ), .C(clk16MHz), 
           .D(n29998));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i50 (.Q(\data_in_frame[6][1] ), .C(clk16MHz), 
           .D(n30001));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i51 (.Q(\data_in_frame[6][2] ), .C(clk16MHz), 
           .D(n30004));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i52 (.Q(\data_in_frame[6][3] ), .C(clk16MHz), 
           .D(n30007));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i2 (.Q(current_limit[2]), .C(clk16MHz), .D(n30299));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i53 (.Q(\data_in_frame[6][4] ), .C(clk16MHz), 
           .D(n30010));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i54 (.Q(\data_in_frame[6][5] ), .C(clk16MHz), 
           .D(n30013));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i55 (.Q(\data_in_frame[6] [6]), .C(clk16MHz), 
           .D(n30016));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i32 (.Q(\data_out_frame[3][7] ), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4972), .S(n56939));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i56 (.Q(\data_in_frame[6] [7]), .C(clk16MHz), 
           .D(n30019));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i57 (.Q(\data_in_frame[7] [0]), .C(clk16MHz), 
           .D(n56157));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i58 (.Q(\data_in_frame[7] [1]), .C(clk16MHz), 
           .D(n30025));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i59 (.Q(\data_in_frame[7] [2]), .C(clk16MHz), 
           .D(n30028));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i60 (.Q(\data_in_frame[7] [3]), .C(clk16MHz), 
           .D(n30031));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i61 (.Q(\data_in_frame[7] [4]), .C(clk16MHz), 
           .D(n30034));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i62 (.Q(\data_in_frame[7] [5]), .C(clk16MHz), 
           .D(n30037));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i63 (.Q(\data_in_frame[7] [6]), .C(clk16MHz), 
           .D(n56163));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i64 (.Q(\data_in_frame[7] [7]), .C(clk16MHz), 
           .D(n56165));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i65 (.Q(\data_in_frame[8] [0]), .C(clk16MHz), 
           .D(n30047));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i66 (.Q(\data_in_frame[8] [1]), .C(clk16MHz), 
           .D(n30050));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i67 (.Q(\data_in_frame[8] [2]), .C(clk16MHz), 
           .D(n30054));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i68 (.Q(\data_in_frame[8] [3]), .C(clk16MHz), 
           .D(n30057));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i3 (.Q(current_limit[3]), .C(clk16MHz), .D(n30282));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i4 (.Q(current_limit[4]), .C(clk16MHz), .D(n30281));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i69 (.Q(\data_in_frame[8] [4]), .C(clk16MHz), 
           .D(n30280));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i70 (.Q(\data_in_frame[8] [5]), .C(clk16MHz), 
           .D(n30063));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i71 (.Q(\data_in_frame[8] [6]), .C(clk16MHz), 
           .D(n30066));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i72 (.Q(\data_in_frame[8] [7]), .C(clk16MHz), 
           .D(n30069));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i73 (.Q(\data_in_frame[9] [0]), .C(clk16MHz), 
           .D(n30072));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i74 (.Q(\data_in_frame[9] [1]), .C(clk16MHz), 
           .D(n30075));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i75 (.Q(\data_in_frame[9] [2]), .C(clk16MHz), 
           .D(n30079));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i76 (.Q(\data_in_frame[9] [3]), .C(clk16MHz), 
           .D(n30082));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i77 (.Q(\data_in_frame[9] [4]), .C(clk16MHz), 
           .D(n30085));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i78 (.Q(\data_in_frame[9] [5]), .C(clk16MHz), 
           .D(n30089));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i79 (.Q(\data_in_frame[9] [6]), .C(clk16MHz), 
           .D(n30092));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i80 (.Q(\data_in_frame[9] [7]), .C(clk16MHz), 
           .D(n30095));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i81 (.Q(\data_in_frame[10]_c [0]), .C(clk16MHz), 
           .D(n30098));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i82 (.Q(\data_in_frame[10][1] ), .C(clk16MHz), 
           .D(n30102));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i83 (.Q(\data_in_frame[10][2] ), .C(clk16MHz), 
           .D(n30105));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i84 (.Q(\data_in_frame[10][3] ), .C(clk16MHz), 
           .D(n30108));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i85 (.Q(\data_in_frame[10] [4]), .C(clk16MHz), 
           .D(n30111));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i86 (.Q(\data_in_frame[10][5] ), .C(clk16MHz), 
           .D(n30114));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i87 (.Q(\data_in_frame[10] [6]), .C(clk16MHz), 
           .D(n30118));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i88 (.Q(\data_in_frame[10][7] ), .C(clk16MHz), 
           .D(n30121));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i89 (.Q(\data_in_frame[11] [0]), .C(clk16MHz), 
           .D(n56297));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i90 (.Q(\data_in_frame[11] [1]), .C(clk16MHz), 
           .D(n56257));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i91 (.Q(\data_in_frame[11] [2]), .C(clk16MHz), 
           .D(n56273));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i92 (.Q(\data_in_frame[11] [3]), .C(clk16MHz), 
           .D(n56283));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i93 (.Q(\data_in_frame[11] [4]), .C(clk16MHz), 
           .D(n30136));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i94 (.Q(\data_in_frame[11] [5]), .C(clk16MHz), 
           .D(n30139));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i95 (.Q(\data_in_frame[11] [6]), .C(clk16MHz), 
           .D(n30142));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i96 (.Q(\data_in_frame[11] [7]), .C(clk16MHz), 
           .D(n30146));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i97 (.Q(\data_in_frame[12] [0]), .C(clk16MHz), 
           .D(n30149));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i98 (.Q(\data_in_frame[12] [1]), .C(clk16MHz), 
           .D(n30152));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i5 (.Q(current_limit[5]), .C(clk16MHz), .D(n30250));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i99 (.Q(\data_in_frame[12] [2]), .C(clk16MHz), 
           .D(n30156));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i100 (.Q(\data_in_frame[12] [3]), .C(clk16MHz), 
           .D(n56303));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i101 (.Q(\data_in_frame[12] [4]), .C(clk16MHz), 
           .D(n56343));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i102 (.Q(\data_in_frame[12] [5]), .C(clk16MHz), 
           .D(n30166));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i103 (.Q(\data_in_frame[12] [6]), .C(clk16MHz), 
           .D(n30169));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i104 (.Q(\data_in_frame[12] [7]), .C(clk16MHz), 
           .D(n30172));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i105 (.Q(\data_in_frame[13] [0]), .C(clk16MHz), 
           .D(n30176));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i106 (.Q(\data_in_frame[13] [1]), .C(clk16MHz), 
           .D(n30179));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i107 (.Q(\data_in_frame[13] [2]), .C(clk16MHz), 
           .D(n30182));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i108 (.Q(\data_in_frame[13] [3]), .C(clk16MHz), 
           .D(n30186));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i109 (.Q(\data_in_frame[13] [4]), .C(clk16MHz), 
           .D(n30189));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i110 (.Q(\data_in_frame[13] [5]), .C(clk16MHz), 
           .D(n30192));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i111 (.Q(\data_in_frame[13] [6]), .C(clk16MHz), 
           .D(n30196));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i146 (.Q(\data_in_frame[18] [1]), .C(clk16MHz), 
           .D(n56075));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i147 (.Q(\data_in_frame[18] [2]), .C(clk16MHz), 
           .D(n56071));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i6 (.Q(current_limit[6]), .C(clk16MHz), .D(n30232));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i148 (.Q(\data_in_frame[18] [3]), .C(clk16MHz), 
           .D(n29540));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i149 (.Q(\data_in_frame[18] [4]), .C(clk16MHz), 
           .D(n29543));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i150 (.Q(\data_in_frame[18] [5]), .C(clk16MHz), 
           .D(n29546));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i151 (.Q(\data_in_frame[18] [6]), .C(clk16MHz), 
           .D(n56065));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i152 (.Q(\data_in_frame[18] [7]), .C(clk16MHz), 
           .D(n56061));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i153 (.Q(\data_in_frame[19][0] ), .C(clk16MHz), 
           .D(n56057));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i154 (.Q(\data_in_frame[19][1] ), .C(clk16MHz), 
           .D(n56053));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i155 (.Q(\data_in_frame[19][2] ), .C(clk16MHz), 
           .D(n56049));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i156 (.Q(\data_in_frame[19][3] ), .C(clk16MHz), 
           .D(n30207));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i157 (.Q(\data_in_frame[19][4] ), .C(clk16MHz), 
           .D(n56045));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i158 (.Q(\data_in_frame[19][5] ), .C(clk16MHz), 
           .D(n56041));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i159 (.Q(\data_in_frame[19] [6]), .C(clk16MHz), 
           .D(n56037));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i160 (.Q(\data_in_frame[19]_c [7]), .C(clk16MHz), 
           .D(n56067));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i161 (.Q(\data_in_frame[20] [0]), .C(clk16MHz), 
           .D(n29579));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i162 (.Q(\data_in_frame[20] [1]), .C(clk16MHz), 
           .D(n30199));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i163 (.Q(\data_in_frame[20] [2]), .C(clk16MHz), 
           .D(n30195));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i164 (.Q(\data_in_frame[20] [3]), .C(clk16MHz), 
           .D(n29588));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i165 (.Q(\data_in_frame[20] [4]), .C(clk16MHz), 
           .D(n29591));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1400 (.I0(n52637), .I1(\data_in_frame[17] [6]), 
            .I2(\data_in_frame[20] [0]), .I3(GND_net), .O(n57101));
    defparam i2_3_lut_adj_1400.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i166 (.Q(\data_in_frame[20] [5]), .C(clk16MHz), 
           .D(n29594));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i167 (.Q(\data_in_frame[20] [6]), .C(clk16MHz), 
           .D(n30155));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1401 (.I0(n52615), .I1(\data_in_frame[19][5] ), 
            .I2(\data_in_frame[19]_c [7]), .I3(GND_net), .O(n57550));
    defparam i2_3_lut_adj_1401.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1402 (.I0(n57701), .I1(\data_in_frame[13] [1]), 
            .I2(\data_in_frame[15] [5]), .I3(n57777), .O(n10_adj_4794));
    defparam i4_4_lut_adj_1402.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1403 (.I0(\data_in_frame[18] [1]), .I1(n25128), 
            .I2(GND_net), .I3(GND_net), .O(n57302));
    defparam i1_2_lut_adj_1403.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i168 (.Q(\data_in_frame[20] [7]), .C(clk16MHz), 
           .D(n29600));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i169 (.Q(\data_in_frame[21] [0]), .C(clk16MHz), 
           .D(n29609));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1404 (.I0(n10), .I1(n145), .I2(GND_net), .I3(GND_net), 
            .O(n107));
    defparam i1_2_lut_adj_1404.LUT_INIT = 16'h4444;
    SB_LUT4 i2_3_lut_adj_1405 (.I0(n51613), .I1(n26286), .I2(\data_in_frame[11] [5]), 
            .I3(GND_net), .O(n51706));
    defparam i2_3_lut_adj_1405.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i170 (.Q(\data_in_frame[21] [1]), .C(clk16MHz), 
           .D(n29614));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1406 (.I0(\data_in_frame[12] [7]), .I1(n25853), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4973));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1406.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i171 (.Q(\data_in_frame[21] [2]), .C(clk16MHz), 
           .D(n29618));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1407 (.I0(\data_in_frame[10] [6]), .I1(n26683), 
            .I2(\data_in_frame[11] [1]), .I3(n6_adj_4973), .O(n57442));   // verilog/coms.v(74[16:27])
    defparam i4_4_lut_adj_1407.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1408 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n57068));
    defparam i1_2_lut_adj_1408.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1409 (.I0(n26482), .I1(n51646), .I2(GND_net), 
            .I3(GND_net), .O(n52626));
    defparam i1_2_lut_adj_1409.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1410 (.I0(\data_in_frame[12] [0]), .I1(\data_in_frame[11] [4]), 
            .I2(\data_in_frame[7] [3]), .I3(\data_in_frame[11] [3]), .O(n61924));
    defparam i1_4_lut_adj_1410.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i172 (.Q(\data_in_frame[21] [3]), .C(clk16MHz), 
           .D(n29621));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1411 (.I0(\data_in_frame[11] [2]), .I1(n61924), 
            .I2(\data_in_frame[11] [0]), .I3(\data_in_frame[11] [7]), .O(n61926));
    defparam i1_4_lut_adj_1411.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1412 (.I0(n57352), .I1(n57765), .I2(n61926), 
            .I3(n57259), .O(n61932));
    defparam i1_4_lut_adj_1412.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i173 (.Q(\data_in_frame[21] [4]), .C(clk16MHz), 
           .D(n29629));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1413 (.I0(n57738), .I1(n57361), .I2(n57442), 
            .I3(n61932), .O(n61938));
    defparam i1_4_lut_adj_1413.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1414 (.I0(n52626), .I1(n25820), .I2(n26031), 
            .I3(n26683), .O(n62012));
    defparam i1_4_lut_adj_1414.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1415 (.I0(n57134), .I1(n57707), .I2(n57467), 
            .I3(n61938), .O(n61944));
    defparam i1_4_lut_adj_1415.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1416 (.I0(n61944), .I1(n59504), .I2(n62012), 
            .I3(n57331), .O(n59380));
    defparam i1_4_lut_adj_1416.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1417 (.I0(n51706), .I1(n57723), .I2(n57534), 
            .I3(\data_in_frame[13] [5]), .O(n58909));
    defparam i1_4_lut_adj_1417.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1418 (.I0(n58909), .I1(\data_in_frame[15][7] ), 
            .I2(n57534), .I3(n59380), .O(n57777));
    defparam i1_4_lut_adj_1418.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_4_lut_adj_1419 (.I0(n51745), .I1(n52327), .I2(n23668), 
            .I3(n51605), .O(n14_adj_4771));
    defparam i5_3_lut_4_lut_adj_1419.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1420 (.I0(\data_in_frame[8] [7]), .I1(n57274), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4974));
    defparam i1_2_lut_adj_1420.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i174 (.Q(\data_in_frame[21] [5]), .C(clk16MHz), 
           .D(n29632));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1421 (.I0(\data_in_frame[11] [3]), .I1(n26266), 
            .I2(n57271), .I3(n6_adj_4974), .O(n25952));
    defparam i4_4_lut_adj_1421.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1422 (.I0(n57750), .I1(n26449), .I2(\data_in_frame[16][2] ), 
            .I3(n57777), .O(n10_adj_4975));
    defparam i4_4_lut_adj_1422.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1423 (.I0(n25952), .I1(n10_adj_4975), .I2(\data_in_frame[16][1] ), 
            .I3(GND_net), .O(n51926));
    defparam i5_3_lut_adj_1423.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4976), .S(n56938));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i26903_4_lut (.I0(n172), .I1(n107), .I2(rx_data[6]), .I3(\data_in_frame[4] [6]), 
            .O(n40837));   // verilog/coms.v(94[13:20])
    defparam i26903_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i21016_3_lut_4_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n30420));
    defparam i21016_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_DFFESS data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk16MHz), 
            .E(n30739), .D(n2_adj_4977), .S(n29117));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk16MHz), 
            .E(n30740), .D(n2_adj_4978), .S(n29116));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk16MHz), 
            .E(n30741), .D(n2_adj_4979), .S(n29115));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_adj_1424 (.I0(n51826), .I1(\data_in_frame[18] [3]), 
            .I2(n51926), .I3(GND_net), .O(n57389));
    defparam i1_3_lut_adj_1424.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1425 (.I0(\data_in_frame[21] [1]), .I1(\data_in_frame[21] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n25991));
    defparam i1_2_lut_adj_1425.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4980), .S(n56937));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1426 (.I0(\data_in_frame[19][0] ), .I1(n59024), 
            .I2(GND_net), .I3(GND_net), .O(n57497));
    defparam i1_2_lut_adj_1426.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1427 (.I0(n59574), .I1(\data_in_frame[16][7] ), 
            .I2(\data_in_frame[17] [0]), .I3(GND_net), .O(n57686));
    defparam i2_3_lut_adj_1427.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1428 (.I0(n25938), .I1(n26428), .I2(\data_in_frame[10][5] ), 
            .I3(GND_net), .O(n26683));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1428.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i175 (.Q(\data_in_frame[21] [6]), .C(clk16MHz), 
           .D(n29651));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1429 (.I0(\data_in_frame[12] [4]), .I1(n26683), 
            .I2(GND_net), .I3(GND_net), .O(n25864));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1429.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1430 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[15][0] ), 
            .I2(GND_net), .I3(GND_net), .O(n57720));
    defparam i1_2_lut_adj_1430.LUT_INIT = 16'h6666;
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk16MHz), .D(n29509));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1431 (.I0(\data_in_frame[19][2] ), .I1(n52653), 
            .I2(n10_adj_13), .I3(\data_in_frame[17] [0]), .O(n57128));
    defparam i1_4_lut_adj_1431.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_adj_1432 (.I0(\data_in_frame[14] [6]), .I1(n57408), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4982));
    defparam i2_2_lut_adj_1432.LUT_INIT = 16'h6666;
    SB_DFFR deadband_i0_i0 (.Q(deadband[0]), .C(clk16MHz), .D(n29505), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_4_lut_adj_1433 (.I0(\data_in_frame[18] [7]), .I1(n7_adj_4982), 
            .I2(\data_in_frame[19][1] ), .I3(n8_adj_4863), .O(n59024));
    defparam i2_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1434 (.I0(n59024), .I1(n57128), .I2(GND_net), 
            .I3(GND_net), .O(n52745));
    defparam i1_2_lut_adj_1434.LUT_INIT = 16'h9999;
    SB_DFFESS data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4983), .S(n56936));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1435 (.I0(n52747), .I1(\data_in_frame[21] [3]), 
            .I2(n52745), .I3(GND_net), .O(n57494));
    defparam i2_3_lut_adj_1435.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1436 (.I0(n52655), .I1(n57408), .I2(\data_in_frame[16] [4]), 
            .I3(GND_net), .O(n52594));
    defparam i2_3_lut_adj_1436.LUT_INIT = 16'h6969;
    SB_DFFESS data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4984), .S(n56935));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i23 (.Q(setpoint[23]), .C(clk16MHz), .E(n27737), 
            .D(n4762[23]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1437 (.I0(n59380), .I1(\data_in_frame[13] [7]), 
            .I2(\data_in_frame[13] [6]), .I3(n26449), .O(n57723));
    defparam i1_2_lut_3_lut_4_lut_adj_1437.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1438 (.I0(n57188), .I1(n57593), .I2(\data_in_frame[10][3] ), 
            .I3(\data_in_frame[8] [2]), .O(n12_adj_4985));   // verilog/coms.v(81[16:27])
    defparam i5_4_lut_adj_1438.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1439 (.I0(\data_in_frame[8] [1]), .I1(n12_adj_4985), 
            .I2(n57616), .I3(\data_in_frame[6][1] ), .O(n26482));   // verilog/coms.v(81[16:27])
    defparam i6_4_lut_adj_1439.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1440 (.I0(n52017), .I1(\data_in_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n57473));
    defparam i1_2_lut_adj_1440.LUT_INIT = 16'h6666;
    SB_DFFER setpoint_i0_i22 (.Q(setpoint[22]), .C(clk16MHz), .E(n27737), 
            .D(n4762[22]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i21 (.Q(setpoint[21]), .C(clk16MHz), .E(n27737), 
            .D(n4762[21]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i20 (.Q(setpoint[20]), .C(clk16MHz), .E(n27737), 
            .D(n4762[20]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i19 (.Q(setpoint[19]), .C(clk16MHz), .E(n27737), 
            .D(n4762[19]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i18 (.Q(setpoint[18]), .C(clk16MHz), .E(n27737), 
            .D(n4762[18]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i17 (.Q(setpoint[17]), .C(clk16MHz), .E(n27737), 
            .D(n4762[17]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i16 (.Q(setpoint[16]), .C(clk16MHz), .E(n27737), 
            .D(n4762[16]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i15 (.Q(setpoint[15]), .C(clk16MHz), .E(n27737), 
            .D(n4762[15]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_193_i2_4_lut (.I0(\data_out_frame[24] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4986));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_193_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFER setpoint_i0_i14 (.Q(setpoint[14]), .C(clk16MHz), .E(n27737), 
            .D(n4762[14]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i13 (.Q(setpoint[13]), .C(clk16MHz), .E(n27737), 
            .D(n4762[13]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i12 (.Q(setpoint[12]), .C(clk16MHz), .E(n27737), 
            .D(n4762[12]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i11 (.Q(setpoint[11]), .C(clk16MHz), .E(n27737), 
            .D(n4762[11]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i10 (.Q(setpoint[10]), .C(clk16MHz), .E(n27737), 
            .D(n4762[10]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i9 (.Q(setpoint[9]), .C(clk16MHz), .E(n27737), 
            .D(n4762[9]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i8 (.Q(setpoint[8]), .C(clk16MHz), .E(n27737), 
            .D(n4762[8]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i7 (.Q(setpoint[7]), .C(clk16MHz), .E(n27737), 
            .D(n4762[7]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1441 (.I0(n59574), .I1(n52017), .I2(\data_in_frame[16] [6]), 
            .I3(n52594), .O(n57226));
    defparam i1_2_lut_3_lut_4_lut_adj_1441.LUT_INIT = 16'h6996;
    SB_DFFER setpoint_i0_i6 (.Q(setpoint[6]), .C(clk16MHz), .E(n27737), 
            .D(n4762[6]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i5 (.Q(setpoint[5]), .C(clk16MHz), .E(n27737), 
            .D(n4762[5]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i4 (.Q(setpoint[4]), .C(clk16MHz), .E(n27737), 
            .D(n4762[4]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i3 (.Q(setpoint[3]), .C(clk16MHz), .E(n27737), 
            .D(n4762[3]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i2 (.Q(setpoint[2]), .C(clk16MHz), .E(n27737), 
            .D(n4762[2]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i1 (.Q(setpoint[1]), .C(clk16MHz), .E(n27737), 
            .D(n4762[1]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS \FRAME_MATCHER.state_FSM_i9  (.Q(\FRAME_MATCHER.i_31__N_2507 ), 
            .C(clk16MHz), .D(n69553), .S(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i8  (.Q(\FRAME_MATCHER.i_31__N_2508 ), 
            .C(clk16MHz), .D(n27011), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i7  (.Q(\FRAME_MATCHER.i_31__N_2509 ), 
            .C(clk16MHz), .D(n2048), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i6  (.Q(\FRAME_MATCHER.state[3] ), .C(clk16MHz), 
            .D(n2049), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i5  (.Q(\FRAME_MATCHER.i_31__N_2511 ), 
            .C(clk16MHz), .D(n20371), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i4  (.Q(\FRAME_MATCHER.i_31__N_2512 ), 
            .C(clk16MHz), .D(n55927), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i3  (.Q(\FRAME_MATCHER.i_31__N_2513 ), 
            .C(clk16MHz), .D(n2060), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i2  (.Q(\FRAME_MATCHER.i_31__N_2514 ), 
            .C(clk16MHz), .D(n27014), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 i1_2_lut_adj_1442 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n25899));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1442.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4987), .S(n56934));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1443 (.I0(\data_in_frame[20] [6]), .I1(n57441), 
            .I2(n51588), .I3(n57474), .O(n57463));
    defparam i3_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1444 (.I0(n52234), .I1(n26815), .I2(n25889), 
            .I3(GND_net), .O(n57467));
    defparam i2_3_lut_adj_1444.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_192_i2_4_lut (.I0(\data_out_frame[24] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4988));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_192_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1445 (.I0(\data_in_frame[9] [7]), .I1(n57467), 
            .I2(GND_net), .I3(GND_net), .O(n52607));
    defparam i1_2_lut_adj_1445.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1446 (.I0(n57576), .I1(n4_adj_4989), .I2(GND_net), 
            .I3(GND_net), .O(n57482));
    defparam i2_2_lut_adj_1446.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1447 (.I0(n25746), .I1(\data_in_frame[7] [6]), 
            .I2(\data_in_frame[8] [1]), .I3(\data_in_frame[10][2] ), .O(n62292));
    defparam i1_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4990), .S(n56933));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1448 (.I0(n57482), .I1(n57437), .I2(n25889), 
            .I3(n62292), .O(n51646));
    defparam i1_4_lut_adj_1448.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4991), .S(n56932));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1449 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n57259));
    defparam i1_2_lut_adj_1449.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4992), .S(n56931));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4993), .S(n56930));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1450 (.I0(\data_in_frame[14] [4]), .I1(n57259), 
            .I2(n25820), .I3(n51646), .O(n52017));
    defparam i3_4_lut_adj_1450.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1451 (.I0(n57662), .I1(\data_in_frame[10][1] ), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4994));
    defparam i2_2_lut_adj_1451.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1452 (.I0(\data_in_frame[14] [3]), .I1(\data_in_frame[12] [2]), 
            .I2(n6_adj_4994), .I3(n52607), .O(n57408));
    defparam i1_4_lut_adj_1452.LUT_INIT = 16'h9669;
    SB_LUT4 i52647_2_lut_3_lut_4_lut (.I0(n23938), .I1(\data_in_frame[7] [6]), 
            .I2(n57229), .I3(\data_in_frame[9] [7]), .O(n68333));   // verilog/coms.v(99[12:25])
    defparam i52647_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1453 (.I0(n51600), .I1(n57209), .I2(n25762), 
            .I3(\data_in_frame[11] [5]), .O(n12_adj_4995));
    defparam i5_4_lut_adj_1453.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1454 (.I0(\data_in_frame[14] [1]), .I1(n12_adj_4995), 
            .I2(n57602), .I3(n57576), .O(n57750));
    defparam i6_4_lut_adj_1454.LUT_INIT = 16'h9669;
    SB_LUT4 select_777_Select_191_i2_4_lut (.I0(\data_out_frame[23] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4996));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_191_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1455 (.I0(n57750), .I1(\data_in_frame[13] [7]), 
            .I2(n52655), .I3(GND_net), .O(n52651));
    defparam i2_3_lut_adj_1455.LUT_INIT = 16'h6969;
    SB_DFFESS data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4997), .S(n56929));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4998), .S(n56928));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4999), .S(n56927));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5000), .S(n56926));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5001), .S(n56925));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5002), .S(n56924));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_777_Select_190_i2_4_lut (.I0(\data_out_frame[23] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5003));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_190_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1456 (.I0(\data_in_frame[16] [3]), .I1(n52651), 
            .I2(GND_net), .I3(GND_net), .O(n57433));
    defparam i1_2_lut_adj_1456.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5004), .S(n56923));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5005), .S(n56922));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5006), .S(n56921));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1457 (.I0(n57226), .I1(\data_in_frame[18] [5]), 
            .I2(\data_in_frame[19][0] ), .I3(n57433), .O(n10_adj_4843));
    defparam i4_4_lut_adj_1457.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5007), .S(n56920));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5008), .S(n56919));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk16MHz), .D(n29480));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_4_lut_adj_1458 (.I0(n25169), .I1(n57463), .I2(n4_adj_4830), 
            .I3(\data_in_frame[21] [0]), .O(n57704));
    defparam i2_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1459 (.I0(\data_in_frame[16]_c [0]), .I1(\data_in_frame[13] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n57701));
    defparam i1_2_lut_adj_1459.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1460 (.I0(\data_in_frame[11] [6]), .I1(n23938), 
            .I2(GND_net), .I3(GND_net), .O(n57707));
    defparam i1_2_lut_adj_1460.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1271));   // verilog/coms.v(88[17:28])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1461 (.I0(\data_in_frame[9] [3]), .I1(n57209), 
            .I2(\data_in_frame[11] [4]), .I3(GND_net), .O(n25971));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_adj_1461.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1462 (.I0(\data_in_frame[14] [0]), .I1(n57707), 
            .I2(n25707), .I3(n26458), .O(n57125));
    defparam i3_4_lut_adj_1462.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1463 (.I0(n51613), .I1(n57367), .I2(n6_adj_4795), 
            .I3(\data_in_frame[9] [7]), .O(n57662));
    defparam i1_4_lut_adj_1463.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1464 (.I0(\data_in_frame[3][1] ), .I1(\data_in_frame[5] [3]), 
            .I2(\data_in_frame[7] [5]), .I3(n57726), .O(n10_adj_5009));   // verilog/coms.v(73[16:69])
    defparam i4_4_lut_adj_1464.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1465 (.I0(\data_in_frame[3][3] ), .I1(n10_adj_5009), 
            .I2(\data_in_frame[5] [4]), .I3(GND_net), .O(n52234));   // verilog/coms.v(73[16:69])
    defparam i5_3_lut_adj_1465.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1466 (.I0(n57331), .I1(\data_in_frame[11] [7]), 
            .I2(n52234), .I3(GND_net), .O(n57367));
    defparam i2_3_lut_adj_1466.LUT_INIT = 16'h9696;
    SB_LUT4 i4_2_lut_adj_1467 (.I0(\data_in_frame[6][3] ), .I1(\data_in_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_5010));
    defparam i4_2_lut_adj_1467.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1468 (.I0(n57573), .I1(\data_in_frame[8] [3]), 
            .I2(\data_in_frame[8] [2]), .I3(\data_in_frame[1] [6]), .O(n24_adj_5011));
    defparam i10_4_lut_adj_1468.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1469 (.I0(\data_in_frame[4] [2]), .I1(n57367), 
            .I2(\data_in_frame[12] [0]), .I3(n25868), .O(n22_adj_5012));
    defparam i8_4_lut_adj_1469.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1470 (.I0(\data_in_frame[8] [0]), .I1(n24_adj_5011), 
            .I2(n18_adj_5010), .I3(n57160), .O(n26_adj_5013));
    defparam i12_4_lut_adj_1470.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1471 (.I0(n68333), .I1(n26_adj_5013), .I2(n22_adj_5012), 
            .I3(\data_in_frame[1] [7]), .O(n57602));
    defparam i13_4_lut_adj_1471.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1472 (.I0(\data_in_frame[10]_c [0]), .I1(\data_in_frame[9] [6]), 
            .I2(n68333), .I3(GND_net), .O(n25820));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1472.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1473 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n57765));
    defparam i1_2_lut_adj_1473.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_1474 (.I0(n57522), .I1(n57108), .I2(n57262), 
            .I3(\data_in_frame[11] [6]), .O(n26_adj_5014));
    defparam i11_4_lut_adj_1474.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1475 (.I0(n57058), .I1(n25820), .I2(n57289), 
            .I3(n57602), .O(n24_adj_5015));
    defparam i9_4_lut_adj_1475.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1476 (.I0(n57163), .I1(n57765), .I2(\data_in_frame[7] [1]), 
            .I3(n57650), .O(n25_adj_5016));
    defparam i10_4_lut_adj_1476.LUT_INIT = 16'h6996;
    SB_LUT4 i8_3_lut_adj_1477 (.I0(\data_in_frame[5] [0]), .I1(\data_in_frame[14] [2]), 
            .I2(n57662), .I3(GND_net), .O(n23_adj_5017));
    defparam i8_3_lut_adj_1477.LUT_INIT = 16'h9696;
    SB_LUT4 i14_4_lut_adj_1478 (.I0(n23_adj_5017), .I1(n25_adj_5016), .I2(n24_adj_5015), 
            .I3(n26_adj_5014), .O(n52655));
    defparam i14_4_lut_adj_1478.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1479 (.I0(\data_in_frame[16][2] ), .I1(\data_in_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5018));
    defparam i1_2_lut_adj_1479.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1480 (.I0(n57125), .I1(n25971), .I2(Kp_23__N_1271), 
            .I3(n6_adj_5018), .O(n57143));
    defparam i4_4_lut_adj_1480.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1481 (.I0(n57143), .I1(n52655), .I2(GND_net), 
            .I3(GND_net), .O(n57441));
    defparam i1_2_lut_adj_1481.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1482 (.I0(n51745), .I1(n52327), .I2(\data_out_frame[20] [4]), 
            .I3(GND_net), .O(n51730));
    defparam i1_2_lut_3_lut_adj_1482.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_214_i3_3_lut_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(n25105), .I2(\FRAME_MATCHER.state[3] ), .I3(n57395), .O(n3_adj_5019));
    defparam select_777_Select_214_i3_3_lut_4_lut.LUT_INIT = 16'h6090;
    SB_LUT4 i1_4_lut_adj_1483 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[23] [5]), 
            .I2(neopxl_color[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5020));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1483.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_adj_1484 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26266));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1484.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1485 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n25707));
    defparam i1_2_lut_adj_1485.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1486 (.I0(\data_in_frame[9] [0]), .I1(Kp_23__N_974), 
            .I2(\data_in_frame[9] [1]), .I3(GND_net), .O(n25762));
    defparam i2_3_lut_adj_1486.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1487 (.I0(n26298), .I1(n25762), .I2(\data_in_frame[11] [2]), 
            .I3(GND_net), .O(n57680));
    defparam i2_3_lut_adj_1487.LUT_INIT = 16'h9696;
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk16MHz), .D(n29478));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1488 (.I0(n26193), .I1(n57097), .I2(n57333), 
            .I3(\data_in_frame[7] [4]), .O(n57650));
    defparam i1_4_lut_adj_1488.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1489 (.I0(\data_in_frame[4] [3]), .I1(n57157), 
            .I2(\data_in_frame[4] [4]), .I3(\data_in_frame[1] [7]), .O(Kp_23__N_878));   // verilog/coms.v(73[16:69])
    defparam i3_4_lut_adj_1489.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1490 (.I0(\data_in_frame[2] [7]), .I1(n35660), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n26193));
    defparam i1_3_lut_adj_1490.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1491 (.I0(n26652), .I1(n57726), .I2(n62190), 
            .I3(n57531), .O(n59504));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1491.LUT_INIT = 16'h6996;
    SB_LUT4 i52643_2_lut (.I0(n59504), .I1(\data_in_frame[7] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n68329));   // verilog/coms.v(99[12:25])
    defparam i52643_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1492 (.I0(\data_in_frame[6][3] ), .I1(\data_in_frame[6][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n25903));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1492.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1493 (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[0] [6]), 
            .I2(n35660), .I3(\data_in_frame[3][0] ), .O(n57097));
    defparam i1_4_lut_adj_1493.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1494 (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(reset), .I3(n3470), .O(n56625));
    defparam i1_2_lut_4_lut_adj_1494.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_adj_1495 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n57058));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1495.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1496 (.I0(\data_in_frame[6][0] ), .I1(n57599), 
            .I2(\data_in_frame[6][1] ), .I3(GND_net), .O(n57262));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_adj_1496.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1497 (.I0(n57115), .I1(\data_in_frame[2] [7]), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[2] [2]), .O(n62248));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1497.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1498 (.I0(\data_in_frame[3][3] ), .I1(\data_in_frame[5] [6]), 
            .I2(\data_in_frame[3][5] ), .I3(\data_in_frame[5] [7]), .O(n61990));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1498.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1499 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[4] [6]), 
            .I2(\data_in_frame[4] [0]), .I3(GND_net), .O(n61988));   // verilog/coms.v(81[16:27])
    defparam i1_3_lut_adj_1499.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1500 (.I0(n61988), .I1(n61990), .I2(\data_in_frame[4] [5]), 
            .I3(\data_in_frame[3] [7]), .O(n61994));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1500.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1501 (.I0(n62248), .I1(Kp_23__N_760), .I2(n57118), 
            .I3(n57557), .O(n62254));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1501.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1502 (.I0(n57567), .I1(n57531), .I2(n61994), 
            .I3(n57311), .O(n62000));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1502.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1503 (.I0(n57157), .I1(n62000), .I2(n62256), 
            .I3(n62254), .O(n62002));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1503.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5020), .S(n56832));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5003), .S(n56833));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1504 (.I0(n62002), .I1(n57097), .I2(n57229), 
            .I3(n26329), .O(n57163));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1504.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1505 (.I0(Kp_23__N_799), .I1(n57163), .I2(n57262), 
            .I3(n57619), .O(n57576));
    defparam i1_4_lut_adj_1505.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1506 (.I0(n26415), .I1(n57576), .I2(\data_in_frame[5] [6]), 
            .I3(GND_net), .O(n57437));
    defparam i1_3_lut_adj_1506.LUT_INIT = 16'h6969;
    SB_LUT4 i1_3_lut_adj_1507 (.I0(\data_in_frame[5] [4]), .I1(n57333), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n25746));
    defparam i1_3_lut_adj_1507.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1508 (.I0(\data_in_frame[7] [6]), .I1(n57229), 
            .I2(GND_net), .I3(GND_net), .O(n23942));
    defparam i1_2_lut_adj_1508.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1509 (.I0(n57150), .I1(n57160), .I2(\data_in_frame[1] [5]), 
            .I3(GND_net), .O(Kp_23__N_872));   // verilog/coms.v(73[16:69])
    defparam i2_3_lut_adj_1509.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1510 (.I0(\data_in_frame[6][4] ), .I1(\data_in_frame[8] [5]), 
            .I2(\data_in_frame[6][3] ), .I3(n6_adj_4808), .O(n25853));   // verilog/coms.v(78[16:43])
    defparam i4_4_lut_adj_1510.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4996), .S(n56834));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1511 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n25893));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_adj_1511.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1512 (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[5] [5]), 
            .I2(\data_in_frame[3][3] ), .I3(n4_adj_5021), .O(n4_adj_4989));
    defparam i1_4_lut_adj_1512.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1513 (.I0(\data_in_frame[1] [5]), .I1(n4_adj_4989), 
            .I2(GND_net), .I3(GND_net), .O(n25868));
    defparam i2_2_lut_adj_1513.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1514 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[3][5] ), 
            .I2(GND_net), .I3(GND_net), .O(n57206));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1514.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1515 (.I0(n25804), .I1(n26335), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_799));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1515.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1516 (.I0(\data_in_frame[4] [7]), .I1(n26329), 
            .I2(n26652), .I3(n6_adj_5022), .O(n57274));   // verilog/coms.v(73[16:27])
    defparam i4_4_lut_adj_1516.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1517 (.I0(\data_in_frame[4] [5]), .I1(n57274), 
            .I2(GND_net), .I3(GND_net), .O(n26286));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1517.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1518 (.I0(n25853), .I1(n25938), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1067));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1518.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1519 (.I0(\data_in_frame[8] [0]), .I1(n57593), 
            .I2(n57206), .I3(n26390), .O(n25889));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1519.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1520 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[3][4] ), .I3(GND_net), .O(n25906));   // verilog/coms.v(79[16:43])
    defparam i1_3_lut_adj_1520.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4988), .S(n56835));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1521 (.I0(\data_in_frame[5] [6]), .I1(n25906), 
            .I2(GND_net), .I3(GND_net), .O(n57616));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1521.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1522 (.I0(\data_in_frame[3][6] ), .I1(\data_in_frame[6][0] ), 
            .I2(GND_net), .I3(GND_net), .O(n26390));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1522.LUT_INIT = 16'h6666;
    SB_DFFESS data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4986), .S(n56836));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1523 (.I0(n26390), .I1(n57616), .I2(n57253), 
            .I3(\data_in_frame[1] [4]), .O(n26815));   // verilog/coms.v(79[16:43])
    defparam i3_4_lut_adj_1523.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4970), .S(n56837));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1524 (.I0(\data_in_frame[4] [6]), .I1(n26335), 
            .I2(\data_in_frame[7] [0]), .I3(\data_in_frame[6] [6]), .O(n57289));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1524.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1525 (.I0(\data_in_frame[4] [4]), .I1(n25804), 
            .I2(n26363), .I3(GND_net), .O(n26332));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1525.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1526 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[2] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n57557));
    defparam i1_2_lut_adj_1526.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_1527 (.I0(\data_in_frame[5] [1]), .I1(\data_in_frame[5] [0]), 
            .I2(\data_in_frame[2] [5]), .I3(GND_net), .O(n14_adj_5023));
    defparam i5_3_lut_adj_1527.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1528 (.I0(n57557), .I1(\data_in_frame[7] [2]), 
            .I2(\data_in_frame[3][0] ), .I3(n57122), .O(n15_adj_5024));
    defparam i6_4_lut_adj_1528.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1529 (.I0(n15_adj_5024), .I1(\data_in_frame[0] [2]), 
            .I2(n14_adj_5023), .I3(\data_in_frame[4] [6]), .O(n26458));
    defparam i8_4_lut_adj_1529.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n56736));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_DFFESS data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4969), .S(n56838));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1530 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n25915));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1530.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1531 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n57253));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1531.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1532 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[3][6] ), 
            .I2(\data_in_frame[1] [4]), .I3(GND_net), .O(n57311));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_adj_1532.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1533 (.I0(n57055), .I1(n57188), .I2(n26415), 
            .I3(GND_net), .O(n25924));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_adj_1533.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4956), .S(n56839));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4955), .S(n56840));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4954), .S(n56772));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1534 (.I0(\data_in_frame[1] [5]), .I1(n25915), 
            .I2(\data_in_frame[2] [0]), .I3(n6_adj_5025), .O(Kp_23__N_869));   // verilog/coms.v(81[16:27])
    defparam i4_4_lut_adj_1534.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4953), .S(n56782));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1535 (.I0(n25924), .I1(n26815), .I2(\data_in_frame[8] [2]), 
            .I3(GND_net), .O(n4_c));   // verilog/coms.v(79[16:43])
    defparam i2_3_lut_adj_1535.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1536 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[4] [1]), .I3(GND_net), .O(n25671));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1536.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4952), .S(n56841));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1537 (.I0(\data_in_frame[8] [3]), .I1(Kp_23__N_869), 
            .I2(\data_in_frame[6][2] ), .I3(n25924), .O(n26428));   // verilog/coms.v(78[16:43])
    defparam i3_4_lut_adj_1537.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1538 (.I0(\data_in_frame[8] [7]), .I1(\data_in_frame[8] [1]), 
            .I2(\data_in_frame[8] [6]), .I3(GND_net), .O(n57573));
    defparam i2_3_lut_adj_1538.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4950), .S(n56842));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1539 (.I0(n26298), .I1(n26458), .I2(GND_net), 
            .I3(GND_net), .O(n26724));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_adj_1539.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i176 (.Q(\data_in_frame[21] [7]), .C(clk16MHz), 
           .D(n29655));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4949), .S(n56843));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4948), .S(n56844));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4947), .S(n56918));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1540 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[7] [3]), .I3(GND_net), .O(n14_adj_4833));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1540.LUT_INIT = 16'h9696;
    SB_LUT4 i26904_3_lut (.I0(n40837), .I1(\data_in_frame[4] [6]), .I2(reset), 
            .I3(GND_net), .O(n29967));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i26904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1541 (.I0(n25889), .I1(n57738), .I2(Kp_23__N_974), 
            .I3(n62074), .O(n62080));
    defparam i1_4_lut_adj_1541.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1542 (.I0(n51600), .I1(n52662), .I2(n26470), 
            .I3(n62080), .O(n59043));
    defparam i1_4_lut_adj_1542.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1543 (.I0(\data_in_frame[9] [7]), .I1(n57522), 
            .I2(\data_in_frame[9] [6]), .I3(n25707), .O(Kp_23__N_1080));   // verilog/coms.v(88[17:63])
    defparam i3_4_lut_adj_1543.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1544 (.I0(n59043), .I1(n57331), .I2(\data_in_frame[10][7] ), 
            .I3(GND_net), .O(n57134));
    defparam i1_3_lut_adj_1544.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4928), .S(n56917));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4926), .S(n56916));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4925), .S(n56915));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4921), .S(n56845));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4920), .S(n56846));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4919), .S(n56847));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_4915), .S(n56848));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_adj_1545 (.I0(n7_adj_4826), .I1(n57134), .I2(Kp_23__N_1080), 
            .I3(GND_net), .O(n51720));
    defparam i1_3_lut_adj_1545.LUT_INIT = 16'h9696;
    SB_DFFESS data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4913), .S(n56754));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4798), .S(n56755));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i211 (.Q(\data_out_frame[26][2] ), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4770), .S(n56756));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4767), .S(n56752));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5026), .S(n56757));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5027), .S(n56750));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5019), .S(n56758));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4766), .S(n56759));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4757), .S(n56760));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4755), .S(n56761));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i219 (.Q(\data_out_frame[27][2] ), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4738), .S(n56762));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4737), .S(n56753));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_4731), .S(n56749));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5028), .S(n56751));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk16MHz), 
            .E(n2873), .D(n3), .S(n56763));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1546 (.I0(Kp_23__N_878), .I1(n57108), .I2(\data_in_frame[6][4] ), 
            .I3(GND_net), .O(Kp_23__N_974));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_adj_1546.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1547 (.I0(n25903), .I1(Kp_23__N_872), .I2(Kp_23__N_869), 
            .I3(\data_in_frame[8] [4]), .O(n25938));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1547.LUT_INIT = 16'h6996;
    SB_DFFESS tx_transmit_4011 (.Q(r_SM_Main_2__N_3545[0]), .C(clk16MHz), 
            .E(n2873), .D(n1), .S(n28912));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5029), .S(n56776));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS LED_4014 (.Q(LED_c), .C(clk16MHz), .E(n2873), .D(n5), 
            .S(n28911));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk16MHz), 
            .E(n2873), .D(n3_adj_5030), .S(n56764));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i1 (.Q(\byte_transmit_counter[1] ), 
            .C(clk16MHz), .E(n2873), .D(n1_adj_5031), .S(n56738));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i2 (.Q(\byte_transmit_counter[2] ), 
            .C(clk16MHz), .E(n2873), .D(n1_adj_5032), .S(n56739));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk16MHz), 
            .E(n2873), .D(n1_adj_5033), .S(n56740));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk16MHz), 
            .E(n2873), .D(n1_adj_5034), .S(n56741));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk16MHz), 
            .E(n2873), .D(n1_adj_5035), .S(n56742));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk16MHz), 
            .E(n2873), .D(n1_adj_5036), .S(n56743));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1548 (.I0(Kp_23__N_974), .I1(n57404), .I2(\data_in_frame[11] [0]), 
            .I3(\data_in_frame[10][7] ), .O(n57683));
    defparam i1_4_lut_adj_1548.LUT_INIT = 16'h6996;
    SB_DFFESS byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk16MHz), 
            .E(n2873), .D(n1_adj_5037), .S(n56737));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5038), .S(n56914));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS driver_enable_4015 (.Q(DE_c), .C(clk16MHz), .E(n2873), .D(n26912), 
            .S(n28901));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1549 (.I0(n57404), .I1(n57680), .I2(GND_net), 
            .I3(GND_net), .O(n52688));
    defparam i1_2_lut_adj_1549.LUT_INIT = 16'h6666;
    SB_DFFESS byte_transmit_counter_i0_i0 (.Q(\byte_transmit_counter[0] ), 
            .C(clk16MHz), .E(n2873), .D(n1_adj_5039), .S(n56744));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5040), .S(n56913));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5041), .S(n56912));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 data_in_frame_17__7__I_0_4040_2_lut (.I0(\data_in_frame[17] [7]), 
            .I1(\data_in_frame[17] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1389));   // verilog/coms.v(73[16:27])
    defparam data_in_frame_17__7__I_0_4040_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_53721 (.I0(byte_transmit_counter[3]), 
            .I1(n69207), .I2(n65479), .I3(byte_transmit_counter[4]), .O(n69336));
    defparam byte_transmit_counter_3__bdd_4_lut_53721.LUT_INIT = 16'he4aa;
    SB_DFFESS data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5042), .S(n56911));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1550 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[15][4] ), 
            .I2(\data_in_frame[13] [2]), .I3(\data_in_frame[13] [3]), .O(n62268));
    defparam i1_4_lut_adj_1550.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1551 (.I0(n52688), .I1(n57683), .I2(n25938), 
            .I3(n62268), .O(n60027));
    defparam i1_4_lut_adj_1551.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5043), .S(n56910));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1552 (.I0(n59636), .I1(n57635), .I2(GND_net), 
            .I3(GND_net), .O(n57490));
    defparam i1_2_lut_adj_1552.LUT_INIT = 16'h9999;
    SB_DFFE data_in_frame_0___i40 (.Q(\data_in_frame[4] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29969));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk16MHz), 
            .E(n2873), .D(n2_adj_5044), .S(n56909));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1553 (.I0(n57490), .I1(\data_in_frame[22] [4]), 
            .I2(\data_in_frame[20] [3]), .I3(n57710), .O(n10_adj_5045));
    defparam i4_4_lut_adj_1553.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1554 (.I0(\data_in_frame[20] [5]), .I1(n8_adj_4828), 
            .I2(\data_in_frame[18] [2]), .I3(\data_in_frame[18] [4]), .O(n59238));
    defparam i4_4_lut_adj_1554.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1555 (.I0(\data_in_frame[21] [1]), .I1(n57704), 
            .I2(n59162), .I3(\data_in_frame[23] [2]), .O(n58846));
    defparam i3_4_lut_adj_1555.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1556 (.I0(\data_in_frame[20] [2]), .I1(n10_adj_5045), 
            .I2(\data_in_frame[18] [2]), .I3(GND_net), .O(n58857));
    defparam i5_3_lut_adj_1556.LUT_INIT = 16'h9696;
    SB_LUT4 n69336_bdd_4_lut (.I0(n69336), .I1(n69267), .I2(n7_adj_5046), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n69336_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_777_Select_54_i2_4_lut (.I0(\data_out_frame[6] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5008));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_54_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1557 (.I0(n58857), .I1(n58846), .I2(n59238), 
            .I3(n59777), .O(n61950));
    defparam i1_4_lut_adj_1557.LUT_INIT = 16'h0008;
    SB_LUT4 i1_4_lut_adj_1558 (.I0(\data_in_frame[21] [2]), .I1(n61950), 
            .I2(n57494), .I3(\data_in_frame[23] [4]), .O(n61952));
    defparam i1_4_lut_adj_1558.LUT_INIT = 16'h8448;
    SB_LUT4 i1_4_lut_adj_1559 (.I0(n52747), .I1(n61952), .I2(n57500), 
            .I3(\data_in_frame[23] [3]), .O(n61954));
    defparam i1_4_lut_adj_1559.LUT_INIT = 16'h8448;
    SB_LUT4 i3_4_lut_adj_1560 (.I0(\data_in_frame[21] [7]), .I1(n57550), 
            .I2(n57101), .I3(\data_in_frame[22] [1]), .O(n59473));
    defparam i3_4_lut_adj_1560.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_53_i2_4_lut (.I0(\data_out_frame[6] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5007));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_53_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1561 (.I0(n59473), .I1(\data_in_frame[22] [5]), 
            .I2(n61954), .I3(n57389), .O(n61958));
    defparam i1_4_lut_adj_1561.LUT_INIT = 16'h4010;
    SB_LUT4 i1_3_lut_adj_1562 (.I0(\data_in_frame[21] [0]), .I1(\data_in_frame[20] [6]), 
            .I2(\data_in_frame[22] [7]), .I3(GND_net), .O(n62202));
    defparam i1_3_lut_adj_1562.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1563 (.I0(n62202), .I1(n57223), .I2(\data_in_frame[18] [5]), 
            .I3(\data_in_frame[18] [4]), .O(n62206));
    defparam i1_4_lut_adj_1563.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1564 (.I0(n52695), .I1(n52745), .I2(n52594), 
            .I3(n62206), .O(n62214));
    defparam i1_4_lut_adj_1564.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_52_i2_4_lut (.I0(\data_out_frame[6] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5006));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_52_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_51_i2_4_lut (.I0(\data_out_frame[6] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5005));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_51_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_50_i2_4_lut (.I0(\data_out_frame[6] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5004));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_50_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1565 (.I0(n57519), .I1(n51826), .I2(n57500), 
            .I3(n62214), .O(n62220));
    defparam i1_4_lut_adj_1565.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1566 (.I0(n59141), .I1(n61958), .I2(n57519), 
            .I3(\data_in_frame[22] [0]), .O(n61960));
    defparam i1_4_lut_adj_1566.LUT_INIT = 16'h8448;
    SB_LUT4 i3_4_lut_adj_1567 (.I0(\data_in_frame[23] [5]), .I1(n57223), 
            .I2(n52745), .I3(n23898), .O(n59377));
    defparam i3_4_lut_adj_1567.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1568 (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[20] [1]), 
            .I2(\data_in_frame[22] [2]), .I3(GND_net), .O(n62232));
    defparam i1_3_lut_adj_1568.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_49_i2_4_lut (.I0(\data_out_frame[6] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5002));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_49_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1569 (.I0(n57238), .I1(n57372), .I2(\data_in_frame[21] [6]), 
            .I3(\data_in_frame[23] [7]), .O(n59440));
    defparam i1_4_lut_adj_1569.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1570 (.I0(\data_in_frame[23] [6]), .I1(n59377), 
            .I2(n57168), .I3(n61960), .O(n61964));
    defparam i1_4_lut_adj_1570.LUT_INIT = 16'h8400;
    SB_LUT4 i1_4_lut_adj_1571 (.I0(n57238), .I1(n57783), .I2(n57550), 
            .I3(n62220), .O(n59860));
    defparam i1_4_lut_adj_1571.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_48_i2_4_lut (.I0(\data_out_frame[6] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5001));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_48_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1572 (.I0(n57101), .I1(n57476), .I2(n59212), 
            .I3(n62232), .O(n59259));
    defparam i1_4_lut_adj_1572.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1573 (.I0(\data_in_frame[20] [1]), .I1(\data_in_frame[22] [3]), 
            .I2(\data_in_frame[20] [2]), .I3(GND_net), .O(n62110));
    defparam i1_3_lut_adj_1573.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_47_i2_4_lut (.I0(\data_out_frame[5] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5000));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_47_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i11_3_lut_4_lut (.I0(rx_data[0]), .I1(\data_in_frame[16]_c [0]), 
            .I2(reset), .I3(n92), .O(n56177));   // verilog/coms.v(94[13:20])
    defparam i11_3_lut_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 select_777_Select_46_i2_4_lut (.I0(\data_out_frame[5] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4999));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_46_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1574 (.I0(n59259), .I1(n59860), .I2(n61964), 
            .I3(n59440), .O(n61970));
    defparam i1_4_lut_adj_1574.LUT_INIT = 16'h0010;
    SB_LUT4 i1_2_lut_adj_1575 (.I0(n57704), .I1(\data_in_frame[23] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n62170));
    defparam i1_2_lut_adj_1575.LUT_INIT = 16'h6666;
    SB_LUT4 select_777_Select_45_i2_4_lut (.I0(\data_out_frame[5] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4998));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_45_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_44_i2_4_lut (.I0(\data_out_frame[5] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4997));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_44_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_43_i2_4_lut (.I0(\data_out_frame[5] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4993));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_43_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_42_i2_4_lut (.I0(\data_out_frame[5] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4992));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_42_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1576 (.I0(n57302), .I1(n57710), .I2(n57635), 
            .I3(n62110), .O(n62116));
    defparam i1_4_lut_adj_1576.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1577 (.I0(\data_in_frame[23] [1]), .I1(n62170), 
            .I2(n61970), .I3(n57292), .O(n61974));
    defparam i1_4_lut_adj_1577.LUT_INIT = 16'h8010;
    SB_LUT4 select_777_Select_41_i2_4_lut (.I0(\data_out_frame[5] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4991));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_41_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1578 (.I0(n61974), .I1(n62116), .I2(\data_in_frame[19]_c [7]), 
            .I3(n57476), .O(n33761));
    defparam i1_4_lut_adj_1578.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_53617 (.I0(byte_transmit_counter[3]), 
            .I1(n69213), .I2(n65421), .I3(byte_transmit_counter[4]), .O(n69330));
    defparam byte_transmit_counter_3__bdd_4_lut_53617.LUT_INIT = 16'he4aa;
    SB_LUT4 select_777_Select_40_i2_4_lut (.I0(\data_out_frame[5] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4990));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_40_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1579 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[4] [7]), 
            .I2(ID[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_4987));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1579.LUT_INIT = 16'ha088;
    SB_LUT4 i51242_4_lut (.I0(n69201), .I1(n69219), .I2(byte_transmit_counter[3]), 
            .I3(\byte_transmit_counter[2] ), .O(n66928));
    defparam i51242_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i47012_3_lut (.I0(n69237), .I1(n66928), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(tx_data[4]));
    defparam i47012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46724_2_lut (.I0(n26298), .I1(n25938), .I2(GND_net), .I3(GND_net), 
            .O(n62400));
    defparam i46724_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6688_4_lut (.I0(\FRAME_MATCHER.i_31__N_2514 ), .I1(n1951), 
            .I2(n59002), .I3(n4452), .O(n20366));   // verilog/coms.v(148[4] 304[11])
    defparam i6688_4_lut.LUT_INIT = 16'ha0a2;
    SB_LUT4 i6_4_lut_adj_1580 (.I0(n57619), .I1(\data_in_frame[8] [1]), 
            .I2(n57055), .I3(n57599), .O(n15_adj_5047));
    defparam i6_4_lut_adj_1580.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1581 (.I0(n20366), .I1(n1951), .I2(n22702), .I3(n62408), 
            .O(n27014));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1581.LUT_INIT = 16'hbbba;
    SB_LUT4 i1_2_lut_adj_1582 (.I0(n52662), .I1(\data_in_frame[8] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n52467));
    defparam i1_2_lut_adj_1582.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1583 (.I0(n62400), .I1(n4_c), .I2(n26428), .I3(n57482), 
            .O(n16_adj_5048));
    defparam i7_4_lut_adj_1583.LUT_INIT = 16'h0100;
    SB_LUT4 i6_4_lut_adj_1584 (.I0(n26286), .I1(n52467), .I2(n59777), 
            .I3(n25853), .O(n15_adj_5049));
    defparam i6_4_lut_adj_1584.LUT_INIT = 16'h0004;
    SB_LUT4 i2_4_lut_adj_1585 (.I0(n62406), .I1(n52234), .I2(n23938), 
            .I3(n68329), .O(n8_adj_5050));
    defparam i2_4_lut_adj_1585.LUT_INIT = 16'h0010;
    SB_LUT4 i8_4_lut_adj_1586 (.I0(n15_adj_5047), .I1(n57163), .I2(n14_adj_5051), 
            .I3(n26335), .O(n59689));
    defparam i8_4_lut_adj_1586.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1587 (.I0(Kp_23__N_974), .I1(n15_adj_5049), .I2(\data_in_frame[8] [6]), 
            .I3(n16_adj_5048), .O(n7_adj_5052));
    defparam i1_4_lut_adj_1587.LUT_INIT = 16'h8400;
    SB_LUT4 i456_2_lut (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), .I2(GND_net), 
            .I3(GND_net), .O(n2060));   // verilog/coms.v(148[4] 304[11])
    defparam i456_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46652_4_lut (.I0(n1951), .I1(n1954), .I2(n3303), .I3(n1957), 
            .O(n62323));   // verilog/coms.v(139[4] 141[7])
    defparam i46652_4_lut.LUT_INIT = 16'h0a02;
    SB_LUT4 i1_4_lut_adj_1588 (.I0(\FRAME_MATCHER.i_31__N_2512 ), .I1(n1954), 
            .I2(n62323), .I3(n59835), .O(n55927));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1588.LUT_INIT = 16'hb3a0;
    SB_LUT4 i5_4_lut_adj_1589 (.I0(n23942), .I1(n7_adj_5052), .I2(n59689), 
            .I3(n8_adj_5050), .O(n33769));
    defparam i5_4_lut_adj_1589.LUT_INIT = 16'h0800;
    SB_LUT4 i6693_4_lut (.I0(n1955), .I1(\FRAME_MATCHER.state[3] ), .I2(n1957), 
            .I3(n25483), .O(n20371));   // verilog/coms.v(148[4] 304[11])
    defparam i6693_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i1_2_lut_adj_1590 (.I0(Kp_23__N_1748), .I1(n33761), .I2(GND_net), 
            .I3(GND_net), .O(n27696));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1590.LUT_INIT = 16'h8888;
    SB_LUT4 i445_2_lut (.I0(\FRAME_MATCHER.state_31__N_2612 [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(GND_net), .I3(GND_net), .O(n2049));   // verilog/coms.v(148[4] 304[11])
    defparam i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i444_2_lut (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), .I2(GND_net), 
            .I3(GND_net), .O(n2048));   // verilog/coms.v(148[4] 304[11])
    defparam i444_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_adj_1591 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5053));
    defparam i2_2_lut_adj_1591.LUT_INIT = 16'heeee;
    SB_LUT4 i28943_4_lut (.I0(n6_adj_5054), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n6_adj_5053), .I3(n25401), .O(n771));   // verilog/coms.v(160[9:60])
    defparam i28943_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i1_2_lut_adj_1592 (.I0(\FRAME_MATCHER.i [4]), .I1(n25580), .I2(GND_net), 
            .I3(GND_net), .O(n25401));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_adj_1592.LUT_INIT = 16'heeee;
    SB_LUT4 i28944_4_lut (.I0(n8_adj_12), .I1(\FRAME_MATCHER.i [31]), .I2(n25401), 
            .I3(\FRAME_MATCHER.i[3] ), .O(n3303));   // verilog/coms.v(230[9:54])
    defparam i28944_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i2_2_lut_adj_1593 (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(GND_net), .I3(GND_net), .O(n22702));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_adj_1593.LUT_INIT = 16'h4444;
    SB_LUT4 i3_2_lut_adj_1594 (.I0(n25483), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n27585));   // verilog/coms.v(148[4] 304[11])
    defparam i3_2_lut_adj_1594.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1595 (.I0(n4452), .I1(n27585), .I2(\FRAME_MATCHER.i_31__N_2514 ), 
            .I3(n22702), .O(n59226));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1595.LUT_INIT = 16'hffdc;
    SB_LUT4 i1_4_lut_adj_1596 (.I0(n25488), .I1(n1957), .I2(n1955), .I3(n59226), 
            .O(n27011));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1596.LUT_INIT = 16'hbaaa;
    SB_LUT4 i6_4_lut_adj_1597 (.I0(\data_in[0] [1]), .I1(\data_in[1] [2]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_5055));
    defparam i6_4_lut_adj_1597.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1598 (.I0(\data_in[1] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [3]), .O(n17_adj_5056));
    defparam i7_4_lut_adj_1598.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1599 (.I0(n17_adj_5056), .I1(\data_in[3] [7]), 
            .I2(n16_adj_5055), .I3(\data_in[2] [6]), .O(n25577));
    defparam i9_4_lut_adj_1599.LUT_INIT = 16'hfbff;
    SB_LUT4 i4_4_lut_adj_1600 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_5057));
    defparam i4_4_lut_adj_1600.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1601 (.I0(\data_in[2] [7]), .I1(n10_adj_5057), 
            .I2(\data_in[3] [4]), .I3(GND_net), .O(n25574));
    defparam i5_3_lut_adj_1601.LUT_INIT = 16'hdfdf;
    SB_LUT4 i5_3_lut_adj_1602 (.I0(\data_in[3] [0]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14_adj_5058));
    defparam i5_3_lut_adj_1602.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1603 (.I0(\data_in[0] [6]), .I1(n25574), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15_adj_5059));
    defparam i6_4_lut_adj_1603.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_1604 (.I0(n15_adj_5059), .I1(\data_in[2] [2]), 
            .I2(n14_adj_5058), .I3(\data_in[0] [3]), .O(n25427));
    defparam i8_4_lut_adj_1604.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_2_lut_adj_1605 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5060));
    defparam i2_2_lut_adj_1605.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1606 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_5061));
    defparam i6_4_lut_adj_1606.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_1607 (.I0(\data_in[3] [6]), .I1(n14_adj_5061), 
            .I2(n10_adj_5060), .I3(\data_in[2] [1]), .O(n25513));
    defparam i7_4_lut_adj_1607.LUT_INIT = 16'hfffd;
    SB_LUT4 i8_4_lut_adj_1608 (.I0(\data_in[2] [6]), .I1(\data_in[2] [0]), 
            .I2(n25513), .I3(\data_in[0] [1]), .O(n20_c));
    defparam i8_4_lut_adj_1608.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1609 (.I0(n25427), .I1(\data_in[3] [7]), .I2(\data_in[1] [6]), 
            .I3(\data_in[2] [5]), .O(n19_c));
    defparam i7_4_lut_adj_1609.LUT_INIT = 16'hfeff;
    SB_LUT4 i46829_4_lut (.I0(\data_in[1] [3]), .I1(\data_in[0] [5]), .I2(\data_in[3] [2]), 
            .I3(\data_in[1] [2]), .O(n62506));
    defparam i46829_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut (.I0(n62506), .I1(n19_c), .I2(n20_c), .I3(GND_net), 
            .O(n1951));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i7_4_lut_adj_1610 (.I0(\data_in[2] [4]), .I1(n25513), .I2(\data_in[1] [5]), 
            .I3(n25577), .O(n18_adj_5062));
    defparam i7_4_lut_adj_1610.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1611 (.I0(\data_in[0] [6]), .I1(n18_adj_5062), 
            .I2(\data_in[3] [0]), .I3(n25574), .O(n20_adj_5063));
    defparam i9_4_lut_adj_1611.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut_adj_1612 (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5064));
    defparam i4_2_lut_adj_1612.LUT_INIT = 16'heeee;
    SB_LUT4 i19768_4_lut (.I0(\FRAME_MATCHER.i_31__N_2513 ), .I1(Kp_23__N_1748), 
            .I2(n33769), .I3(n33761), .O(n27737));   // verilog/coms.v(18[27:29])
    defparam i19768_4_lut.LUT_INIT = 16'he420;
    SB_LUT4 i10_4_lut_adj_1613 (.I0(n15_adj_5064), .I1(n20_adj_5063), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n1954));
    defparam i10_4_lut_adj_1613.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut_adj_1614 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n25427), .O(n16_adj_5065));
    defparam i6_4_lut_adj_1614.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1615 (.I0(n25577), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [1]), .O(n17_adj_5066));
    defparam i7_4_lut_adj_1615.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1616 (.I0(n17_adj_5066), .I1(\data_in[3] [5]), 
            .I2(n16_adj_5065), .I3(\data_in[3] [3]), .O(n1957));
    defparam i9_4_lut_adj_1616.LUT_INIT = 16'hfbff;
    SB_LUT4 i362_2_lut (.I0(n1954), .I1(n1951), .I2(GND_net), .I3(GND_net), 
            .O(n1955));   // verilog/coms.v(142[4] 144[7])
    defparam i362_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1617 (.I0(Kp_23__N_1748), .I1(\FRAME_MATCHER.i_31__N_2513 ), 
            .I2(GND_net), .I3(GND_net), .O(n33763));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1617.LUT_INIT = 16'heeee;
    SB_LUT4 i5_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(GND_net), .I3(GND_net), .O(n28_adj_5067));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1618 (.I0(n43466), .I1(n59359), .I2(\FRAME_MATCHER.i_31__N_2511 ), 
            .I3(n42668), .O(n6_adj_5068));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1618.LUT_INIT = 16'hccec;
    SB_LUT4 i3_4_lut_adj_1619 (.I0(n33763), .I1(n6_adj_5068), .I2(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I3(\FRAME_MATCHER.i_31__N_2509 ), .O(n69553));   // verilog/coms.v(148[4] 304[11])
    defparam i3_4_lut_adj_1619.LUT_INIT = 16'hefee;
    SB_LUT4 i15_4_lut_adj_1620 (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [17]), .O(n38_adj_5069));
    defparam i15_4_lut_adj_1620.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1621 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [30]), 
            .I2(\FRAME_MATCHER.i [29]), .I3(\FRAME_MATCHER.i [24]), .O(n59867));
    defparam i3_4_lut_adj_1621.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1622 (.I0(\FRAME_MATCHER.i [15]), .I1(n59867), 
            .I2(\FRAME_MATCHER.i [28]), .I3(\FRAME_MATCHER.i [26]), .O(n36_adj_5070));
    defparam i13_4_lut_adj_1622.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.i [11]), .I1(n38_adj_5069), .I2(n28_adj_5067), 
            .I3(\FRAME_MATCHER.i [12]), .O(n42));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1623 (.I0(\FRAME_MATCHER.i [25]), .I1(\FRAME_MATCHER.i [7]), 
            .I2(\FRAME_MATCHER.i [19]), .I3(\FRAME_MATCHER.i [9]), .O(n40));
    defparam i17_4_lut_adj_1623.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [27]), .I1(n36_adj_5070), .I2(\FRAME_MATCHER.i [13]), 
            .I3(\FRAME_MATCHER.i [10]), .O(n41));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1624 (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i[5] ), 
            .I2(\FRAME_MATCHER.i [8]), .I3(\FRAME_MATCHER.i [23]), .O(n39));
    defparam i16_4_lut_adj_1624.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n39), .I1(n41), .I2(n40), .I3(n42), .O(n25580));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i28947_4_lut (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n25580), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(262[9:58])
    defparam i28947_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i464_2_lut (.I0(n4452), .I1(\FRAME_MATCHER.i_31__N_2514 ), .I2(GND_net), 
            .I3(GND_net), .O(n2068));   // verilog/coms.v(148[4] 304[11])
    defparam i464_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47160_3_lut (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[17] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62846));
    defparam i47160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47161_3_lut (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[19] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62847));
    defparam i47161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47158_3_lut (.I0(\data_out_frame[22] [0]), .I1(\data_out_frame[23] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62844));
    defparam i47158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47157_3_lut (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[21] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62843));
    defparam i47157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1625 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[4] [6]), 
            .I2(ID[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_4984));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1625.LUT_INIT = 16'ha088;
    SB_LUT4 select_777_Select_37_i2_4_lut (.I0(\data_out_frame[4] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_4983));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_37_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i47169_3_lut (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[17] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62855));
    defparam i47169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47170_3_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[19] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62856));
    defparam i47170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46939_3_lut (.I0(\data_out_frame[22] [7]), .I1(\data_out_frame[23] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62625));
    defparam i46939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_777_Select_36_i2_4_lut (.I0(\data_out_frame[4] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_4980));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_36_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i46938_3_lut (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[21] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62624));
    defparam i46938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_777_Select_35_i2_4_lut (.I0(\data_out_frame[4] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_4979));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_35_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i47145_3_lut (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[17] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62831));
    defparam i47145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_777_Select_34_i2_4_lut (.I0(\data_out_frame[4] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_4978));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_34_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i47146_3_lut (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[19] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62832));
    defparam i47146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47020_3_lut (.I0(\data_out_frame[22] [6]), .I1(\data_out_frame[23] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62706));
    defparam i47020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_777_Select_33_i2_4_lut (.I0(\data_out_frame[4] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_4977));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_33_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i47019_3_lut (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[21] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62705));
    defparam i47019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47133_3_lut (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[17] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62819));
    defparam i47133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_777_Select_32_i2_4_lut (.I0(\data_out_frame[4] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_4976));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_32_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i47134_3_lut (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[19] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62820));
    defparam i47134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47083_3_lut (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[23] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62769));
    defparam i47083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47082_3_lut (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[21] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62768));
    defparam i47082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47112_3_lut (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[17] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62798));
    defparam i47112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47113_3_lut (.I0(\data_out_frame[18] [2]), .I1(\data_out_frame[19] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62799));
    defparam i47113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47116_3_lut (.I0(\data_out_frame[22] [2]), .I1(\data_out_frame[23] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62802));
    defparam i47116_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47115_3_lut (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[21] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62801));
    defparam i47115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47034_3_lut (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[17] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62720));
    defparam i47034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47035_3_lut (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[19] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62721));
    defparam i47035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47038_3_lut (.I0(\data_out_frame[22] [1]), .I1(\data_out_frame[23] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62724));
    defparam i47038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47037_3_lut (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[21] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62723));
    defparam i47037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47043_4_lut (.I0(\data_out_frame[0][4] ), .I1(\data_out_frame[3][4] ), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n62729));
    defparam i47043_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i47181_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62867));
    defparam i47181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47182_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62868));
    defparam i47182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47023_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62709));
    defparam i47023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47022_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62708));
    defparam i47022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26873_4_lut (.I0(n28383), .I1(n106), .I2(rx_data[2]), .I3(\data_in_frame[20] [2]), 
            .O(n40807));   // verilog/coms.v(94[13:20])
    defparam i26873_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i47028_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62714));
    defparam i47028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47029_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62715));
    defparam i47029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26874_3_lut (.I0(n40807), .I1(\data_in_frame[20] [2]), .I2(reset), 
            .I3(GND_net), .O(n30195));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i26874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1626 (.I0(n40970), .I1(n145), .I2(GND_net), .I3(GND_net), 
            .O(n106));
    defparam i1_2_lut_adj_1626.LUT_INIT = 16'h8888;
    SB_LUT4 i26918_4_lut (.I0(n28383), .I1(n106), .I2(rx_data[1]), .I3(\data_in_frame[20] [1]), 
            .O(n40852));   // verilog/coms.v(94[13:20])
    defparam i26918_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i47041_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62727));
    defparam i47041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47040_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62726));
    defparam i47040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i26919_3_lut (.I0(n40852), .I1(\data_in_frame[20] [1]), .I2(reset), 
            .I3(GND_net), .O(n30199));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i26919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47100_3_lut (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[9] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62786));
    defparam i47100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47101_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62787));
    defparam i47101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47104_3_lut (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62790));
    defparam i47104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47103_3_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62789));
    defparam i47103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47121_3_lut (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[9] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62807));
    defparam i47121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1627 (.I0(\data_in_frame[19]_c [7]), .I1(n28379), 
            .I2(n28434), .I3(rx_data[7]), .O(n56067));
    defparam i12_4_lut_adj_1627.LUT_INIT = 16'h3a0a;
    SB_LUT4 i47122_3_lut (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[11] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62808));
    defparam i47122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47068_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62754));
    defparam i47068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47069_4_lut (.I0(n62754), .I1(n28175), .I2(\byte_transmit_counter[2] ), 
            .I3(\data_out_frame[1][0] ), .O(n62755));
    defparam i47069_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i47067_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62753));
    defparam i47067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47143_3_lut (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[15] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62829));
    defparam i47143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47142_3_lut (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[13] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62828));
    defparam i47142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50633_2_lut (.I0(n69303), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n65477));
    defparam i50633_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i47139_3_lut (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[9] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62825));
    defparam i47139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47140_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62826));
    defparam i47140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47032_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62718));
    defparam i47032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47031_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62717));
    defparam i47031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46935_3_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62621));
    defparam i46935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46936_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62622));
    defparam i46936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_779_Select_0_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n1_adj_5039));
    defparam select_779_Select_0_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_779_Select_7_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(byte_transmit_counter[7]), 
            .I3(GND_net), .O(n1_adj_5037));
    defparam select_779_Select_7_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i47191_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62877));
    defparam i47191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_779_Select_6_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(byte_transmit_counter[6]), 
            .I3(GND_net), .O(n1_adj_5036));
    defparam select_779_Select_6_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_779_Select_5_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(byte_transmit_counter[5]), 
            .I3(GND_net), .O(n1_adj_5035));
    defparam select_779_Select_5_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i47190_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62876));
    defparam i47190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_779_Select_4_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(n1_adj_5034));
    defparam select_779_Select_4_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_779_Select_3_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n1_adj_5033));
    defparam select_779_Select_3_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_779_Select_2_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n1_adj_5032));
    defparam select_779_Select_2_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1628 (.I0(\FRAME_MATCHER.i_31__N_2511 ), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n57007));
    defparam i1_2_lut_3_lut_adj_1628.LUT_INIT = 16'hfefe;
    SB_LUT4 select_779_Select_1_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2511 ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(\byte_transmit_counter[1] ), 
            .I3(GND_net), .O(n1_adj_5031));
    defparam select_779_Select_1_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i1_3_lut (.I0(\data_out_frame[0][3] ), 
            .I1(\data_out_frame[1][3] ), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n1_adj_5071));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50136_2_lut (.I0(\data_out_frame[3][3] ), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n65394));
    defparam i50136_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_5072));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i4_3_lut (.I0(\data_out_frame[4] [3]), 
            .I1(\data_out_frame[5] [3]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n4_adj_5073));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14118_3_lut (.I0(\data_out_frame[1][1] ), .I1(\data_out_frame[3][1] ), 
            .I2(\byte_transmit_counter[1] ), .I3(GND_net), .O(n28125));   // verilog/coms.v(109[34:55])
    defparam i14118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47092_3_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[7] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62778));
    defparam i47092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1629 (.I0(current_limit[14]), .I1(current_limit[15]), 
            .I2(n26), .I3(current_limit[13]), .O(n21));   // verilog/TinyFPGA_B.v(251[22:35])
    defparam i1_4_lut_adj_1629.LUT_INIT = 16'h3332;
    SB_LUT4 i47093_4_lut (.I0(n62778), .I1(n28125), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n62779));
    defparam i47093_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i47091_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62777));
    defparam i47091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50259_2_lut (.I0(n69531), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n65421));
    defparam i50259_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i52754_2_lut_3_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), 
            .I2(n43466), .I3(GND_net), .O(tx_transmit_N_3416));
    defparam i52754_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_2_lut_adj_1630 (.I0(n10_adj_11), .I1(\FRAME_MATCHER.i [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5076));
    defparam i1_2_lut_adj_1630.LUT_INIT = 16'heeee;
    SB_LUT4 i14440_4_lut (.I0(n5_adj_5076), .I1(reset), .I2(n57016), .I3(n43293), 
            .O(n57921));
    defparam i14440_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 n69330_bdd_4_lut (.I0(n69330), .I1(n69249), .I2(n7_adj_5077), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n69330_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i50152_3_lut (.I0(current_limit[14]), .I1(n26), .I2(current_limit[13]), 
            .I3(GND_net), .O(n65396));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i50152_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i21742_4_lut (.I0(n21), .I1(n65396), .I2(\current[15] ), .I3(current_limit[15]), 
            .O(n260));   // verilog/TinyFPGA_B.v(250[22:29])
    defparam i21742_4_lut.LUT_INIT = 16'hcafa;
    SB_LUT4 i50264_2_lut_3_lut (.I0(\FRAME_MATCHER.i[5] ), .I1(n8_adj_14), 
            .I2(n130), .I3(GND_net), .O(n65436));
    defparam i50264_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1631 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i[3] ), 
            .I2(\FRAME_MATCHER.i[5] ), .I3(GND_net), .O(n40970));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_3_lut_adj_1631.LUT_INIT = 16'h0202;
    SB_LUT4 i1_3_lut_4_lut_adj_1632 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(n57007), .I3(LED_c), .O(n27274));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1632.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_adj_1633 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n3470));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1633.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1634 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i[3] ), 
            .I2(n3470), .I3(n161), .O(n130));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_3_lut_4_lut_adj_1634.LUT_INIT = 16'h2000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.i[5] ), .I1(n8_adj_14), 
            .I2(n130), .I3(reset), .O(n28428));
    defparam i1_2_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i2_3_lut_4_lut_adj_1635 (.I0(\data_out_frame[11] [5]), .I1(n51541), 
            .I2(n26780), .I3(n26693), .O(n51832));
    defparam i2_3_lut_4_lut_adj_1635.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_31_i2_3_lut (.I0(\data_out_frame[3][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4972));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_31_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_3_lut_adj_1636 (.I0(\data_out_frame[11] [5]), .I1(n51541), 
            .I2(n26394), .I3(GND_net), .O(n52624));
    defparam i1_2_lut_3_lut_adj_1636.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1637 (.I0(byte_transmit_counter[6]), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5079));   // verilog/coms.v(216[6] 223[9])
    defparam i1_2_lut_adj_1637.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1638 (.I0(byte_transmit_counter[4]), .I1(\byte_transmit_counter[0] ), 
            .I2(\byte_transmit_counter[2] ), .I3(\byte_transmit_counter[1] ), 
            .O(n4_adj_5080));
    defparam i1_4_lut_adj_1638.LUT_INIT = 16'ha8a0;
    SB_LUT4 i29557_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[7]), 
            .I2(n4_adj_5080), .I3(n4_adj_5079), .O(n43466));
    defparam i29557_4_lut.LUT_INIT = 16'hffec;
    SB_LUT4 i1_4_lut_4_lut (.I0(reset), .I1(n28417), .I2(\data_in_frame[0] [4]), 
            .I3(rx_data[4]), .O(n56361));   // verilog/coms.v(94[13:20])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i28766_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3545[0]), .I2(GND_net), 
            .I3(GND_net), .O(n42668));
    defparam i28766_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_3_lut_4_lut_adj_1639 (.I0(\data_out_frame[4] [7]), .I1(n57792), 
            .I2(n26662), .I3(n10_adj_4821), .O(n51676));   // verilog/coms.v(88[17:70])
    defparam i5_3_lut_4_lut_adj_1639.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1640 (.I0(n10_adj_11), .I1(n57019), .I2(n40783), 
            .I3(\FRAME_MATCHER.i [0]), .O(n59230));
    defparam i3_4_lut_adj_1640.LUT_INIT = 16'hfeff;
    SB_LUT4 i5_3_lut_4_lut_adj_1641 (.I0(\data_out_frame[4] [7]), .I1(n57792), 
            .I2(\data_out_frame[11] [3]), .I3(n10_adj_4846), .O(n25095));   // verilog/coms.v(88[17:70])
    defparam i5_3_lut_4_lut_adj_1641.LUT_INIT = 16'h6996;
    SB_LUT4 i23230_3_lut_4_lut (.I0(deadband[1]), .I1(\data_in_frame[16][1] ), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29850));
    defparam i23230_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 select_777_Select_30_i2_3_lut (.I0(\data_out_frame[3][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4971));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_30_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i3_4_lut_adj_1642 (.I0(n56625), .I1(\FRAME_MATCHER.i [2]), .I2(n40970), 
            .I3(\FRAME_MATCHER.i [0]), .O(n57046));
    defparam i3_4_lut_adj_1642.LUT_INIT = 16'hbfff;
    SB_LUT4 i23224_3_lut_4_lut (.I0(deadband[0]), .I1(\data_in_frame[16]_c [0]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29505));
    defparam i23224_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i2_2_lut_3_lut_adj_1643 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[7] [4]), 
            .I2(\data_out_frame[9] [6]), .I3(GND_net), .O(n57622));   // verilog/coms.v(77[16:27])
    defparam i2_2_lut_3_lut_adj_1643.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1054_i24_3_lut_4_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[23]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i24_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1054_i23_3_lut_4_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[22]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i23_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1054_i22_3_lut_4_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[21]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i22_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1054_i21_3_lut_4_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[20]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i21_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i3_3_lut_4_lut_adj_1644 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[7] [4]), 
            .I2(\data_out_frame[5] [3]), .I3(n57185), .O(n26066));   // verilog/coms.v(77[16:27])
    defparam i3_3_lut_4_lut_adj_1644.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1054_i20_3_lut_4_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[19]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i20_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1054_i19_3_lut_4_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[18]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i19_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1054_i18_3_lut_4_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[17]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i18_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 select_777_Select_123_i2_4_lut (.I0(\data_out_frame[15] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4945));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_123_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 mux_1054_i17_3_lut_4_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[16]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i17_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1054_i16_3_lut_4_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[15]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i16_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1054_i15_3_lut_4_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[14]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i15_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1054_i14_3_lut_4_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[13]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i14_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1054_i13_3_lut_4_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[12]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i13_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1054_i12_3_lut_4_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[11]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i12_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_4_lut_adj_1645 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[8] [6]), 
            .I2(encoder0_position_scaled[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4823));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1645.LUT_INIT = 16'ha088;
    SB_LUT4 mux_1054_i11_3_lut_4_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[10]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i11_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1054_i10_3_lut_4_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[9]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i10_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 select_777_Select_28_i2_3_lut (.I0(\data_out_frame[3][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4968));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_28_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 mux_1054_i9_3_lut_4_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[8]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i9_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i21869_3_lut_4_lut (.I0(\data_in_frame[19]_c [7]), .I1(\data_in_frame[3] [7]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[7]));
    defparam i21869_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1054_i7_3_lut_4_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3][6] ), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[6]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i7_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1054_i6_3_lut_4_lut (.I0(\data_in_frame[19][5] ), .I1(\data_in_frame[3][5] ), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[5]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i6_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1054_i5_3_lut_4_lut (.I0(\data_in_frame[19][4] ), .I1(\data_in_frame[3][4] ), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[4]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i5_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1054_i4_3_lut_4_lut (.I0(\data_in_frame[19][3] ), .I1(\data_in_frame[3][3] ), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[3]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i4_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1054_i3_3_lut_4_lut (.I0(\data_in_frame[19][2] ), .I1(\data_in_frame[3][2] ), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[2]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i3_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 mux_1054_i2_3_lut_4_lut (.I0(\data_in_frame[19][1] ), .I1(\data_in_frame[3][1] ), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[1]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i2_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i2_3_lut_4_lut_adj_1646 (.I0(n1954), .I1(n1951), .I2(n1957), 
            .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n59359));   // verilog/coms.v(148[4] 304[11])
    defparam i2_3_lut_4_lut_adj_1646.LUT_INIT = 16'h8000;
    SB_LUT4 mux_1054_i1_3_lut_4_lut (.I0(\data_in_frame[19][0] ), .I1(\data_in_frame[3][0] ), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n4762[0]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1054_i1_3_lut_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i1_3_lut_4_lut_adj_1647 (.I0(\FRAME_MATCHER.i_31__N_2511 ), .I1(tx_active), 
            .I2(r_SM_Main_2__N_3545[0]), .I3(n43466), .O(n25483));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1647.LUT_INIT = 16'ha8aa;
    SB_LUT4 i5_3_lut_4_lut_adj_1648 (.I0(n25804), .I1(\data_in_frame[3][6] ), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[3][5] ), .O(n14_adj_5051));
    defparam i5_3_lut_4_lut_adj_1648.LUT_INIT = 16'h6996;
    SB_LUT4 i46730_2_lut_4_lut (.I0(n26458), .I1(\data_in_frame[4] [5]), 
            .I2(n57271), .I3(\data_in_frame[8] [7]), .O(n62406));
    defparam i46730_2_lut_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 select_777_Select_27_i2_3_lut (.I0(\data_out_frame[3][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4967));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_27_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i22862_3_lut_4_lut (.I0(deadband[13]), .I1(\data_in_frame[15] [5]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29838));
    defparam i22862_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 select_777_Select_122_i2_4_lut (.I0(\data_out_frame[15] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4944));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_122_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_69_i2_4_lut (.I0(\data_out_frame[8] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4815));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_69_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_68_i2_4_lut (.I0(\data_out_frame[8] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4814));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_68_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1649 (.I0(n60027), .I1(\data_in_frame[18] [0]), 
            .I2(\data_in_frame[17] [7]), .I3(\data_in_frame[17] [6]), .O(n57710));
    defparam i2_3_lut_4_lut_adj_1649.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1650 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[3][6] ), .I3(\data_in_frame[1] [4]), .O(n6_adj_5025));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_4_lut_adj_1650.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1651 (.I0(\data_in_frame[6][1] ), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[5] [7]), .I3(GND_net), .O(n57055));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1651.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1652 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[4] [0]), .I3(GND_net), .O(n57188));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1652.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1653 (.I0(n25853), .I1(n25938), .I2(\data_in_frame[4] [5]), 
            .I3(n57274), .O(n57738));
    defparam i1_2_lut_4_lut_adj_1653.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1654 (.I0(\data_in_frame[5] [0]), .I1(n25804), 
            .I2(n26335), .I3(GND_net), .O(n26329));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1654.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1655 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[1] [5]), 
            .I2(n4_adj_4989), .I3(GND_net), .O(n57593));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1655.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1656 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[4] [2]), .O(n57567));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_4_lut_adj_1656.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1657 (.I0(n25906), .I1(n26415), .I2(n57576), 
            .I3(\data_in_frame[5] [6]), .O(n52662));
    defparam i1_2_lut_4_lut_adj_1657.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1658 (.I0(reset), .I1(n3470), .I2(GND_net), .I3(GND_net), 
            .O(n57019));
    defparam i1_2_lut_adj_1658.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_1659 (.I0(n10), .I1(n56625), .I2(GND_net), .I3(GND_net), 
            .O(n57041));
    defparam i1_2_lut_adj_1659.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_1660 (.I0(n23938), .I1(\data_in_frame[7] [6]), 
            .I2(n57229), .I3(GND_net), .O(n26470));
    defparam i1_2_lut_3_lut_adj_1660.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1661 (.I0(Kp_23__N_760), .I1(\data_in_frame[2] [6]), 
            .I2(n57650), .I3(\data_in_frame[5] [2]), .O(n23938));
    defparam i1_3_lut_4_lut_adj_1661.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1662 (.I0(n25906), .I1(\data_in_frame[5] [4]), 
            .I2(n57333), .I3(\data_in_frame[5] [5]), .O(n57229));
    defparam i1_2_lut_4_lut_adj_1662.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1663 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[3][2] ), .O(n57333));   // verilog/coms.v(73[16:27])
    defparam i1_3_lut_4_lut_adj_1663.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1664 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[6][3] ), 
            .I2(\data_in_frame[6][2] ), .I3(GND_net), .O(n57599));
    defparam i1_2_lut_3_lut_adj_1664.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1665 (.I0(\data_in_frame[3][1] ), .I1(\data_in_frame[4] [7]), 
            .I2(\data_in_frame[5] [2]), .I3(\data_in_frame[5] [1]), .O(n57531));   // verilog/coms.v(88[17:70])
    defparam i1_3_lut_4_lut_adj_1665.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1666 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[9] [3]), .I3(GND_net), .O(n57522));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1666.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_121_i2_4_lut (.I0(\data_out_frame[15] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4943));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_121_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1667 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[12] [1]), .I3(GND_net), .O(n57352));
    defparam i1_2_lut_3_lut_adj_1667.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1668 (.I0(\data_in_frame[9] [3]), .I1(\data_in_frame[9] [4]), 
            .I2(n59504), .I3(\data_in_frame[7] [3]), .O(n51613));
    defparam i2_3_lut_4_lut_adj_1668.LUT_INIT = 16'h6996;
    SB_LUT4 i14168_2_lut (.I0(\byte_transmit_counter[1] ), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n28175));   // verilog/coms.v(109[34:55])
    defparam i14168_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i47077_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62763));
    defparam i47077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47078_4_lut (.I0(n62763), .I1(n28175), .I2(\byte_transmit_counter[2] ), 
            .I3(\data_out_frame[1][5] ), .O(n62764));
    defparam i47078_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i1_2_lut_3_lut_adj_1669 (.I0(\data_in_frame[9] [2]), .I1(n26298), 
            .I2(n26458), .I3(GND_net), .O(n57209));   // verilog/coms.v(76[16:42])
    defparam i1_2_lut_3_lut_adj_1669.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1670 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(n57474), .I3(n52594), .O(n25169));
    defparam i1_2_lut_4_lut_adj_1670.LUT_INIT = 16'h9669;
    SB_LUT4 select_777_Select_120_i2_4_lut (.I0(\data_out_frame[15] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4942));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_120_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1671 (.I0(n25899), .I1(n57226), .I2(\data_in_frame[19][0] ), 
            .I3(n59024), .O(n52747));
    defparam i1_2_lut_4_lut_adj_1671.LUT_INIT = 16'h9669;
    SB_LUT4 select_777_Select_119_i2_4_lut (.I0(\data_out_frame[14] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4941));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_119_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i47076_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62762));
    defparam i47076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1672 (.I0(n59162), .I1(\data_in_frame[21] [1]), 
            .I2(\data_in_frame[21] [2]), .I3(GND_net), .O(n57500));
    defparam i1_2_lut_3_lut_adj_1672.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1673 (.I0(\data_in_frame[20] [4]), .I1(\data_in_frame[18] [1]), 
            .I2(n25128), .I3(\data_in_frame[20] [3]), .O(n51826));
    defparam i2_3_lut_4_lut_adj_1673.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_118_i2_4_lut (.I0(\data_out_frame[14] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4940));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_118_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1674 (.I0(n60027), .I1(\data_in_frame[15] [5]), 
            .I2(n57401), .I3(GND_net), .O(n52637));
    defparam i1_2_lut_3_lut_adj_1674.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1675 (.I0(\data_out_frame[7] [7]), .I1(n57753), 
            .I2(n57235), .I3(\data_out_frame[17] [0]), .O(n26858));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_4_lut_adj_1675.LUT_INIT = 16'h6996;
    SB_LUT4 i29881125_i1_3_lut (.I0(n69507), .I1(n69231), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n14_adj_4786));
    defparam i29881125_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_777_Select_117_i2_4_lut (.I0(\data_out_frame[14] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4939));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_117_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i51825_3_lut (.I0(n69243), .I1(n69255), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n67511));
    defparam i51825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1676 (.I0(\data_in_frame[15][2] ), .I1(\data_in_frame[12] [6]), 
            .I2(n26031), .I3(\data_in_frame[12] [7]), .O(n57774));
    defparam i2_3_lut_4_lut_adj_1676.LUT_INIT = 16'h6996;
    SB_LUT4 i14110_3_lut (.I0(\data_out_frame[1][6] ), .I1(\data_out_frame[3][6] ), 
            .I2(\byte_transmit_counter[1] ), .I3(GND_net), .O(n28117));   // verilog/coms.v(109[34:55])
    defparam i14110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47071_3_lut (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[7] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62757));
    defparam i47071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47072_4_lut (.I0(n62757), .I1(n28117), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n62758));
    defparam i47072_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i47070_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62756));
    defparam i47070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1677 (.I0(Kp_23__N_1301), .I1(n57404), .I2(n57680), 
            .I3(GND_net), .O(n52705));
    defparam i1_2_lut_3_lut_adj_1677.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1678 (.I0(\data_in_frame[19][5] ), .I1(n59284), 
            .I2(n59141), .I3(n59212), .O(n57372));
    defparam i1_2_lut_4_lut_adj_1678.LUT_INIT = 16'h9669;
    SB_LUT4 i50315_2_lut (.I0(n69195), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n65442));
    defparam i50315_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1679 (.I0(\data_out_frame[7] [7]), .I1(n57753), 
            .I2(\data_out_frame[16] [3]), .I3(GND_net), .O(n57065));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1679.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1680 (.I0(\data_out_frame[7] [7]), .I1(n57753), 
            .I2(n57412), .I3(GND_net), .O(n57413));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1680.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1681 (.I0(\data_out_frame[7] [7]), .I1(n57753), 
            .I2(n26241), .I3(n51805), .O(n59466));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_4_lut_adj_1681.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_116_i2_4_lut (.I0(\data_out_frame[14] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4938));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_116_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_4_lut_adj_1682 (.I0(n59980), .I1(n57128), .I2(n57238), 
            .I3(\data_in_frame[21] [4]), .O(n57168));
    defparam i1_3_lut_4_lut_adj_1682.LUT_INIT = 16'h9669;
    SB_LUT4 select_777_Select_115_i2_4_lut (.I0(\data_out_frame[14] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4937));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_115_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_4_lut_adj_1683 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[18] [3]), 
            .I2(\data_in_frame[17] [7]), .I3(\data_in_frame[20] [0]), .O(n62160));
    defparam i1_3_lut_4_lut_adj_1683.LUT_INIT = 16'h6996;
    SB_LUT4 i14108_3_lut (.I0(\data_out_frame[1][7] ), .I1(\data_out_frame[3][7] ), 
            .I2(\byte_transmit_counter[1] ), .I3(GND_net), .O(n28115));   // verilog/coms.v(109[34:55])
    defparam i14108_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47062_3_lut (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[7] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62748));
    defparam i47062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47063_4_lut (.I0(n62748), .I1(n28115), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n62749));
    defparam i47063_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i47061_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62747));
    defparam i47061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50549_2_lut (.I0(n69225), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n65454));
    defparam i50549_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1684 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4946));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_adj_1684.LUT_INIT = 16'heeee;
    SB_LUT4 i29391_2_lut_3_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(\FRAME_MATCHER.i [2]), .I3(GND_net), .O(n43293));
    defparam i29391_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i50692_2_lut (.I0(\data_out_frame[0][2] ), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n65497));
    defparam i50692_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_777_Select_114_i2_4_lut (.I0(\data_out_frame[14] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4936));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_114_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_113_i2_4_lut (.I0(\data_out_frame[14] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4932));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_113_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i47086_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62772));
    defparam i47086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1685 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[14] [0]), 
            .I2(setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4931));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1685.LUT_INIT = 16'ha088;
    SB_LUT4 i47087_4_lut (.I0(n62772), .I1(n65497), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[1] ), .O(n62773));
    defparam i47087_4_lut.LUT_INIT = 16'ha0ac;
    SB_LUT4 select_777_Select_111_i2_4_lut (.I0(\data_out_frame[13] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4930));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_111_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i47085_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n62771));
    defparam i47085_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23229_3_lut (.I0(n375), .I1(n455), .I2(n11610), .I3(GND_net), 
            .O(n37189));
    defparam i23229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20_4_lut_adj_1686 (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15), .I3(n15_adj_15), .O(n19));
    defparam i20_4_lut_adj_1686.LUT_INIT = 16'h0aca;
    SB_LUT4 i2_2_lut_adj_1687 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5054));
    defparam i2_2_lut_adj_1687.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1688 (.I0(n40970), .I1(n3470), .I2(n161), 
            .I3(n8_adj_14), .O(n28375));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_4_lut_adj_1688.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1689 (.I0(n40970), .I1(n3470), .I2(n161), 
            .I3(n8_adj_12), .O(n56988));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_4_lut_adj_1689.LUT_INIT = 16'h0080;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53741 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[6] [4]), .I2(\data_out_frame[7] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n69318));
    defparam byte_transmit_counter_0__bdd_4_lut_53741.LUT_INIT = 16'he4aa;
    SB_LUT4 i21861_3_lut_4_lut (.I0(\Kp[7] ), .I1(\data_in_frame[3] [7]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29798));
    defparam i21861_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1690 (.I0(n40970), .I1(n3470), .I2(n161), 
            .I3(reset), .O(n40973));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_4_lut_adj_1690.LUT_INIT = 16'h0080;
    SB_LUT4 n69318_bdd_4_lut (.I0(n69318), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[4] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n62730));
    defparam n69318_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1691 (.I0(n26757), .I1(n57671), .I2(\data_out_frame[19] [4]), 
            .I3(n51682), .O(n59521));
    defparam i2_3_lut_4_lut_adj_1691.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1692 (.I0(n26757), .I1(n57671), .I2(n57317), 
            .I3(GND_net), .O(n57644));
    defparam i1_2_lut_3_lut_adj_1692.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1693 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n6_adj_5084));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1693.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1694 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[2] [4]), .I3(GND_net), .O(n25804));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1694.LUT_INIT = 16'h9696;
    SB_LUT4 i16304_3_lut_4_lut (.I0(n8_adj_14), .I1(n57037), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n30312));
    defparam i16304_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16464_3_lut_4_lut (.I0(n8_adj_14), .I1(n57037), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n30472));
    defparam i16464_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16468_3_lut_4_lut (.I0(n8_adj_14), .I1(n57037), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n30476));
    defparam i16468_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16474_3_lut_4_lut (.I0(n8_adj_14), .I1(n57037), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n30482));
    defparam i16474_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15442_3_lut_4_lut (.I0(n8_adj_14), .I1(n57037), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n29450));
    defparam i15442_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(\byte_transmit_counter[1] ), 
            .I1(n4_adj_5073), .I2(n5_adj_5072), .I3(\byte_transmit_counter[2] ), 
            .O(n69312));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i15439_3_lut_4_lut (.I0(n8_adj_14), .I1(n57037), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n29447));
    defparam i15439_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1695 (.I0(n40970), .I1(n3470), .I2(n161), 
            .I3(n8_adj_16), .O(n28381));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_4_lut_adj_1695.LUT_INIT = 16'hff7f;
    SB_LUT4 i15436_3_lut_4_lut (.I0(n8_adj_14), .I1(n57037), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n29444));
    defparam i15436_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15433_3_lut_4_lut (.I0(n8_adj_14), .I1(n57037), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n29441));
    defparam i15433_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1696 (.I0(n40970), .I1(n3470), .I2(n161), 
            .I3(n8), .O(n28379));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_4_lut_adj_1696.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_adj_1697 (.I0(n10_adj_11), .I1(n56625), .I2(GND_net), 
            .I3(GND_net), .O(n57037));
    defparam i1_2_lut_adj_1697.LUT_INIT = 16'heeee;
    SB_LUT4 n69312_bdd_4_lut (.I0(n69312), .I1(n65394), .I2(n1_adj_5071), 
            .I3(\byte_transmit_counter[2] ), .O(n69315));
    defparam n69312_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1698 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(rx_data_ready), .I3(\FRAME_MATCHER.rx_data_ready_prev ), 
            .O(n40783));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_4_lut_adj_1698.LUT_INIT = 16'hffbf;
    SB_LUT4 select_777_Select_213_i3_3_lut_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(n25105), .I2(\FRAME_MATCHER.state[3] ), .I3(n57487), .O(n3_adj_5027));
    defparam select_777_Select_213_i3_3_lut_4_lut.LUT_INIT = 16'h9060;
    SB_LUT4 i15466_3_lut_4_lut (.I0(n28391), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[15][7] ), .O(n29474));
    defparam i15466_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1699 (.I0(n59574), .I1(n52017), .I2(\data_in_frame[16] [6]), 
            .I3(GND_net), .O(n57474));
    defparam i1_2_lut_3_lut_adj_1699.LUT_INIT = 16'h6969;
    SB_LUT4 i15457_3_lut_4_lut (.I0(n28391), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[15][4] ), .O(n29465));
    defparam i15457_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n69528));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n69528_bdd_4_lut (.I0(n69528), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n69531));
    defparam n69528_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15454_3_lut_4_lut (.I0(n28391), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[15][3] ), .O(n29462));
    defparam i15454_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_777_Select_67_i2_4_lut (.I0(\data_out_frame[8] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4736));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_67_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i15451_3_lut_4_lut (.I0(n28391), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[15][2] ), .O(n29459));
    defparam i15451_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15448_3_lut_4_lut (.I0(n28391), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[15][1] ), .O(n29456));
    defparam i15448_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1700 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[2] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n57122));   // verilog/coms.v(80[16:27])
    defparam i1_2_lut_adj_1700.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1701 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[2] [3]), .I3(GND_net), .O(n26335));   // verilog/coms.v(78[16:43])
    defparam i1_3_lut_adj_1701.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1702 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n26363));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_adj_1702.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1703 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [4]), 
            .I2(ID[3]), .I3(ID[4]), .O(n12_adj_5086));   // verilog/coms.v(241[12:32])
    defparam i4_4_lut_adj_1703.LUT_INIT = 16'h7bde;
    SB_LUT4 i15445_3_lut_4_lut (.I0(n28391), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[15][0] ), .O(n29453));
    defparam i15445_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_4_lut_adj_1704 (.I0(\data_in_frame[0] [1]), .I1(ID[6]), .I2(ID[1]), 
            .I3(\data_in_frame[0] [6]), .O(n10_adj_5087));   // verilog/coms.v(241[12:32])
    defparam i2_4_lut_adj_1704.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_1705 (.I0(ID[7]), .I1(\data_in_frame[0] [2]), .I2(\data_in_frame[0] [7]), 
            .I3(ID[2]), .O(n11_adj_5088));   // verilog/coms.v(241[12:32])
    defparam i3_4_lut_adj_1705.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1706 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [5]), 
            .I2(ID[0]), .I3(ID[5]), .O(n9_adj_5089));   // verilog/coms.v(241[12:32])
    defparam i1_4_lut_adj_1706.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_2_lut_4_lut_adj_1707 (.I0(n3470), .I1(n6_adj_5054), .I2(n43293), 
            .I3(n10), .O(n28415));
    defparam i1_2_lut_4_lut_adj_1707.LUT_INIT = 16'hff7f;
    SB_LUT4 i7_4_lut_adj_1708 (.I0(n9_adj_5089), .I1(n11_adj_5088), .I2(n10_adj_5087), 
            .I3(n12_adj_5086), .O(n59777));   // verilog/coms.v(241[12:32])
    defparam i7_4_lut_adj_1708.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1709 (.I0(n3470), .I1(n6_adj_5054), .I2(n43293), 
            .I3(n10_adj_11), .O(n28391));
    defparam i1_2_lut_4_lut_adj_1709.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_adj_1710 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n57118));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_adj_1710.LUT_INIT = 16'h6666;
    SB_LUT4 i5_2_lut_adj_1711 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_760));   // verilog/coms.v(99[12:25])
    defparam i5_2_lut_adj_1711.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53776 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n69522));
    defparam byte_transmit_counter_0__bdd_4_lut_53776.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut_adj_1712 (.I0(Kp_23__N_760), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[0] [6]), .I3(n6_adj_5084), .O(Kp_23__N_748));   // verilog/coms.v(73[16:27])
    defparam i4_4_lut_adj_1712.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1713 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n57115));   // verilog/coms.v(169[9:87])
    defparam i1_2_lut_adj_1713.LUT_INIT = 16'h6666;
    SB_LUT4 i15912_3_lut_4_lut (.I0(n28409), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[3][0] ), .O(n29920));
    defparam i15912_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1714 (.I0(\data_in_frame[0] [0]), .I1(Kp_23__N_748), 
            .I2(GND_net), .I3(GND_net), .O(n57308));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1714.LUT_INIT = 16'h6666;
    SB_LUT4 i15915_3_lut_4_lut (.I0(n28409), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[3][1] ), .O(n29923));
    defparam i15915_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15918_3_lut_4_lut (.I0(n28409), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[3][2] ), .O(n29926));
    defparam i15918_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_1934_i10_2_lut (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5090));   // verilog/coms.v(169[9:87])
    defparam equal_1934_i10_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15921_3_lut_4_lut (.I0(n28409), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[3][3] ), .O(n29929));
    defparam i15921_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15925_3_lut_4_lut (.I0(n28409), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[3][4] ), .O(n29933));
    defparam i15925_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1715 (.I0(n25804), .I1(Kp_23__N_748), .I2(\data_in_frame[2] [1]), 
            .I3(GND_net), .O(n22_adj_5091));
    defparam i5_3_lut_adj_1715.LUT_INIT = 16'h1414;
    SB_LUT4 i10_4_lut_adj_1716 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[1] [6]), .O(n27_adj_5092));
    defparam i10_4_lut_adj_1716.LUT_INIT = 16'h8000;
    SB_LUT4 i15928_3_lut_4_lut (.I0(n28409), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[3][5] ), .O(n29936));
    defparam i15928_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_4_lut_adj_1717 (.I0(\data_in_frame[2] [0]), .I1(n10_adj_5090), 
            .I2(n57308), .I3(\data_in_frame[1] [5]), .O(n26_adj_5093));
    defparam i9_4_lut_adj_1717.LUT_INIT = 16'h2100;
    SB_LUT4 i15931_3_lut_4_lut (.I0(n28409), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[3][6] ), .O(n29939));
    defparam i15931_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_4_lut (.I0(n28409), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n56355));
    defparam i11_4_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12_4_lut_adj_1718 (.I0(n26652), .I1(n24_adj_4927), .I2(\data_in_frame[0] [7]), 
            .I3(n57118), .O(n29));
    defparam i12_4_lut_adj_1718.LUT_INIT = 16'h0440;
    SB_LUT4 i14_4_lut_adj_1719 (.I0(n27_adj_5092), .I1(n59777), .I2(n22_adj_5091), 
            .I3(n26363), .O(n31));
    defparam i14_4_lut_adj_1719.LUT_INIT = 16'h0020;
    SB_LUT4 i16_4_lut_adj_1720 (.I0(n31), .I1(n29), .I2(n62366), .I3(n26_adj_5093), 
            .O(\FRAME_MATCHER.state_31__N_2612 [3]));
    defparam i16_4_lut_adj_1720.LUT_INIT = 16'h0800;
    SB_LUT4 select_777_Select_66_i2_4_lut (.I0(\data_out_frame[8] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_4734));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_66_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i26888_4_lut (.I0(n172), .I1(n107), .I2(rx_data[5]), .I3(\data_in_frame[4] [5]), 
            .O(n40822));   // verilog/coms.v(94[13:20])
    defparam i26888_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53593 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(\byte_transmit_counter[1] ), .O(n69300));
    defparam byte_transmit_counter_0__bdd_4_lut_53593.LUT_INIT = 16'he4aa;
    SB_LUT4 i26889_3_lut (.I0(n40822), .I1(\data_in_frame[4] [5]), .I2(reset), 
            .I3(GND_net), .O(n29964));   // verilog/TinyFPGA_B.v(47[5:10])
    defparam i26889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n69522_bdd_4_lut (.I0(n69522), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n69525));
    defparam n69522_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n69300_bdd_4_lut (.I0(n69300), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(\byte_transmit_counter[1] ), 
            .O(n69303));
    defparam n69300_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 equal_298_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // verilog/coms.v(158[12:15])
    defparam equal_298_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 equal_307_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_16));   // verilog/coms.v(158[12:15])
    defparam equal_307_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i16495_3_lut_4_lut (.I0(n28417), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n30503));
    defparam i16495_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15754_3_lut_4_lut (.I0(n28417), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n29762));
    defparam i15754_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_777_Select_65_i2_4_lut (.I0(\data_out_frame[8] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5044));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_65_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53771 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(\byte_transmit_counter[1] ), .O(n69516));
    defparam byte_transmit_counter_0__bdd_4_lut_53771.LUT_INIT = 16'he4aa;
    SB_LUT4 i15705_3_lut_4_lut (.I0(n28417), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n29713));
    defparam i15705_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n69516_bdd_4_lut (.I0(n69516), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n62815));
    defparam n69516_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15670_3_lut_4_lut (.I0(n28417), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n29678));
    defparam i15670_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i23201_4_lut (.I0(PWMLimit[1]), .I1(n375), .I2(n376), .I3(PWMLimit[0]), 
            .O(n4));
    defparam i23201_4_lut.LUT_INIT = 16'h44d4;
    SB_LUT4 i15658_3_lut_4_lut (.I0(n28417), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n29666));
    defparam i15658_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53766 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(\byte_transmit_counter[1] ), .O(n69510));
    defparam byte_transmit_counter_0__bdd_4_lut_53766.LUT_INIT = 16'he4aa;
    SB_LUT4 i23223_3_lut_4_lut (.I0(n376), .I1(n456), .I2(n455), .I3(n375), 
            .O(n4_adj_17));
    defparam i23223_3_lut_4_lut.LUT_INIT = 16'h40f4;
    SB_LUT4 i24104_3_lut_4_lut (.I0(\Ki[14] ), .I1(\data_in_frame[4] [6]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29776));
    defparam i24104_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_3_lut_adj_1721 (.I0(n59380), .I1(\data_in_frame[13] [7]), 
            .I2(\data_in_frame[13] [6]), .I3(GND_net), .O(n52825));
    defparam i1_2_lut_3_lut_adj_1721.LUT_INIT = 16'h6969;
    SB_LUT4 select_777_Select_25_i2_3_lut (.I0(\data_out_frame[3][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4966));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_25_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_777_Select_15_i2_3_lut (.I0(\data_out_frame[1][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4965));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_15_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_777_Select_14_i2_3_lut (.I0(\data_out_frame[1][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4964));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_14_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n62755), .I3(n62753), 
            .O(n7_adj_5096));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1722 (.I0(\data_out_frame[20] [2]), .I1(n51652), 
            .I2(\data_out_frame[20] [3]), .I3(n23668), .O(n51837));
    defparam i1_2_lut_3_lut_4_lut_adj_1722.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53598 (.I0(\byte_transmit_counter[1] ), 
            .I1(n62876), .I2(n62877), .I3(\byte_transmit_counter[2] ), 
            .O(n69288));
    defparam byte_transmit_counter_1__bdd_4_lut_53598.LUT_INIT = 16'he4aa;
    SB_LUT4 n69510_bdd_4_lut (.I0(n69510), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n62818));
    defparam n69510_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n62779), .I3(n62777), 
            .O(n7_adj_5077));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n62773), .I3(n62771), 
            .O(n7_adj_5046));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n62764), .I3(n62762), 
            .O(n7_adj_4787));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i21021_3_lut (.I0(n30), .I1(PWMLimit[15]), .I2(n361), .I3(GND_net), 
            .O(n32));
    defparam i21021_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1723 (.I0(n40783), .I1(\FRAME_MATCHER.i [0]), 
            .I2(n3470), .I3(n10), .O(n172));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_4_lut_adj_1723.LUT_INIT = 16'hffef;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n62749), .I3(n62747), 
            .O(n7_adj_4784));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(\byte_transmit_counter[1] ), .I2(n62758), .I3(n62756), 
            .O(n7_adj_4785));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i2_3_lut_4_lut_adj_1724 (.I0(\data_out_frame[20] [2]), .I1(n51652), 
            .I2(n59153), .I3(\data_out_frame[22] [3]), .O(n25105));
    defparam i2_3_lut_4_lut_adj_1724.LUT_INIT = 16'h9669;
    SB_LUT4 n69288_bdd_4_lut (.I0(n69288), .I1(n62622), .I2(n62621), .I3(\byte_transmit_counter[2] ), 
            .O(n69291));
    defparam n69288_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_777_Select_13_i2_3_lut (.I0(\data_out_frame[1][5] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4963));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_13_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1725 (.I0(n40783), .I1(\FRAME_MATCHER.i [0]), 
            .I2(n3470), .I3(n40970), .O(n28383));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_3_lut_4_lut_adj_1725.LUT_INIT = 16'hefff;
    SB_LUT4 select_777_Select_64_i2_4_lut (.I0(\data_out_frame[8] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5043));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_64_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1726 (.I0(\data_out_frame[23] [4]), .I1(n59922), 
            .I2(n51617), .I3(GND_net), .O(n57359));
    defparam i1_2_lut_3_lut_adj_1726.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1727 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(Kp_23__N_1301), .I3(n52688), .O(n57401));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_4_lut_adj_1727.LUT_INIT = 16'h9669;
    SB_LUT4 select_777_Select_11_i2_3_lut (.I0(\data_out_frame[1][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4962));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_11_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_777_Select_63_i2_4_lut (.I0(\data_out_frame[7] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5042));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_63_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_777_Select_9_i2_3_lut (.I0(\data_out_frame[1][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4961));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_9_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i50159_2_lut (.I0(n69309), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n65479));
    defparam i50159_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5_3_lut_4_lut_adj_1728 (.I0(\data_out_frame[15] [4]), .I1(n1720), 
            .I2(n10_adj_4791), .I3(n57689), .O(n51652));
    defparam i5_3_lut_4_lut_adj_1728.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_4_lut (.I0(\data_out_frame[21] [7]), .I1(n10_adj_4788), 
            .I2(n51605), .I3(\data_out_frame[22] [6]), .O(n17));
    defparam i3_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53761 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n69504));
    defparam byte_transmit_counter_0__bdd_4_lut_53761.LUT_INIT = 16'he4aa;
    SB_LUT4 select_777_Select_8_i2_3_lut (.I0(\data_out_frame[1][0] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4960));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_8_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_3_lut_adj_1729 (.I0(\data_out_frame[21] [2]), .I1(\data_out_frame[16] [5]), 
            .I2(\data_out_frame[19] [0]), .I3(GND_net), .O(n9_adj_4908));
    defparam i1_2_lut_3_lut_adj_1729.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_4_i2_3_lut (.I0(\data_out_frame[0][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4959));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_4_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_4_lut_adj_1730 (.I0(\data_out_frame[21] [7]), .I1(n10_adj_4788), 
            .I2(n51605), .I3(n25), .O(n57633));
    defparam i1_2_lut_4_lut_adj_1730.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1731 (.I0(\FRAME_MATCHER.i[5] ), .I1(\FRAME_MATCHER.i [4]), 
            .I2(GND_net), .I3(GND_net), .O(n134));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_adj_1731.LUT_INIT = 16'hbbbb;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(156[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 n69504_bdd_4_lut (.I0(n69504), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n69507));
    defparam n69504_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1732 (.I0(n52737), .I1(n68335), .I2(n57674), 
            .I3(n26100), .O(n57606));
    defparam i2_3_lut_4_lut_adj_1732.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1733 (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[12] [3]), 
            .I2(\data_out_frame[5] [7]), .I3(GND_net), .O(n6_adj_4882));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1733.LUT_INIT = 16'h9696;
    SB_LUT4 i49879_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65257));   // verilog/coms.v(158[12:15])
    defparam i49879_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49815_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65258));   // verilog/coms.v(158[12:15])
    defparam i49815_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49816_2_lut (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65259));   // verilog/coms.v(158[12:15])
    defparam i49816_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53579 (.I0(\byte_transmit_counter[1] ), 
            .I1(n62717), .I2(n62718), .I3(\byte_transmit_counter[2] ), 
            .O(n69282));
    defparam byte_transmit_counter_1__bdd_4_lut_53579.LUT_INIT = 16'he4aa;
    SB_LUT4 i15885_3_lut_4_lut (.I0(n8_adj_16), .I1(n57041), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n29893));
    defparam i15885_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_777_Select_62_i2_4_lut (.I0(\data_out_frame[7] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5041));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_62_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1734 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[10] [2]), .I3(n57653), .O(n6_adj_4881));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_4_lut_adj_1734.LUT_INIT = 16'h6996;
    SB_LUT4 i15888_3_lut_4_lut (.I0(n8_adj_16), .I1(n57041), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n29896));
    defparam i15888_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n69282_bdd_4_lut (.I0(n69282), .I1(n62826), .I2(n62825), .I3(\byte_transmit_counter[2] ), 
            .O(n69285));
    defparam n69282_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15891_3_lut_4_lut (.I0(n8_adj_16), .I1(n57041), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n29899));
    defparam i15891_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15895_3_lut_4_lut (.I0(n8_adj_16), .I1(n57041), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n29903));
    defparam i15895_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_777_Select_3_i2_3_lut (.I0(\data_out_frame[0][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4958));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_3_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_3_lut_adj_1735 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[10] [2]), .I3(GND_net), .O(n25731));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_3_lut_adj_1735.LUT_INIT = 16'h9696;
    SB_LUT4 i15898_3_lut_4_lut (.I0(n8_adj_16), .I1(n57041), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n29906));
    defparam i15898_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i49817_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65260));   // verilog/coms.v(158[12:15])
    defparam i49817_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1736 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[6] [2]), .I3(GND_net), .O(n25667));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1736.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1737 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[9] [7]), .O(n57154));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1737.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_61_i2_4_lut (.I0(\data_out_frame[7] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5040));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_61_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i49818_2_lut (.I0(\FRAME_MATCHER.i[5] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65261));   // verilog/coms.v(158[12:15])
    defparam i49818_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15902_3_lut_4_lut (.I0(n8_adj_16), .I1(n57041), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n29910));
    defparam i15902_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i49819_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65262));   // verilog/coms.v(158[12:15])
    defparam i49819_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49820_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65263));   // verilog/coms.v(158[12:15])
    defparam i49820_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15905_3_lut_4_lut (.I0(n8_adj_16), .I1(n57041), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n29913));
    defparam i15905_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_3_lut_4_lut_adj_1738 (.I0(n25918), .I1(n68337), .I2(\data_out_frame[19] [0]), 
            .I3(n51811), .O(n20));
    defparam i7_3_lut_4_lut_adj_1738.LUT_INIT = 16'h9669;
    SB_LUT4 i15909_3_lut_4_lut (.I0(n8_adj_16), .I1(n57041), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n29917));
    defparam i15909_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1739 (.I0(n25918), .I1(n68337), .I2(n59466), 
            .I3(n57171), .O(n59591));
    defparam i2_3_lut_4_lut_adj_1739.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n69171), .I2(n65477), .I3(byte_transmit_counter[4]), .O(n69498));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1740 (.I0(n51656), .I1(n26607), .I2(\data_out_frame[13] [1]), 
            .I3(GND_net), .O(n22_adj_4855));
    defparam i1_2_lut_3_lut_adj_1740.LUT_INIT = 16'h9696;
    SB_LUT4 i49821_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65264));   // verilog/coms.v(158[12:15])
    defparam i49821_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3_2_lut_4_lut_adj_1741 (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[14] [7]), 
            .I2(n57191), .I3(\data_out_frame[12] [5]), .O(n24_adj_4852));
    defparam i3_2_lut_4_lut_adj_1741.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1742 (.I0(\data_out_frame[9] [5]), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[9] [4]), .I3(GND_net), .O(n18_adj_4839));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_3_lut_adj_1742.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1743 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_14));
    defparam i2_3_lut_adj_1743.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_adj_1744 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[5] [6]), .I3(GND_net), .O(n57564));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1744.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1745 (.I0(n59636), .I1(n57143), .I2(n52655), 
            .I3(n57062), .O(n62014));
    defparam i1_2_lut_3_lut_4_lut_adj_1745.LUT_INIT = 16'h6996;
    SB_LUT4 i49822_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65265));   // verilog/coms.v(158[12:15])
    defparam i49822_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49823_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65266));   // verilog/coms.v(158[12:15])
    defparam i49823_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15760_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57046), 
            .I2(rx_data[7]), .I3(\data_in_frame[23] [7]), .O(n29768));
    defparam i15760_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15757_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57046), 
            .I2(rx_data[6]), .I3(\data_in_frame[23] [6]), .O(n29765));
    defparam i15757_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15751_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57046), 
            .I2(rx_data[5]), .I3(\data_in_frame[23] [5]), .O(n29759));
    defparam i15751_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15748_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57046), 
            .I2(rx_data[4]), .I3(\data_in_frame[23] [4]), .O(n29756));
    defparam i15748_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53574 (.I0(\byte_transmit_counter[1] ), 
            .I1(n62828), .I2(n62829), .I3(\byte_transmit_counter[2] ), 
            .O(n69276));
    defparam byte_transmit_counter_1__bdd_4_lut_53574.LUT_INIT = 16'he4aa;
    SB_LUT4 i15732_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57046), 
            .I2(rx_data[3]), .I3(\data_in_frame[23] [3]), .O(n29740));
    defparam i15732_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i49824_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65267));   // verilog/coms.v(158[12:15])
    defparam i49824_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15729_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57046), 
            .I2(rx_data[2]), .I3(\data_in_frame[23] [2]), .O(n29737));
    defparam i15729_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n69498_bdd_4_lut (.I0(n69498), .I1(n69261), .I2(n7_adj_5096), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n69498_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1746 (.I0(\data_in_frame[4] [5]), .I1(n57271), 
            .I2(n59504), .I3(\data_in_frame[7] [3]), .O(n51600));
    defparam i1_2_lut_3_lut_4_lut_adj_1746.LUT_INIT = 16'h6996;
    SB_LUT4 i49825_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65268));   // verilog/coms.v(158[12:15])
    defparam i49825_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15720_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57046), 
            .I2(rx_data[1]), .I3(\data_in_frame[23] [1]), .O(n29728));
    defparam i15720_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i49885_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65275));   // verilog/coms.v(158[12:15])
    defparam i49885_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15691_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57046), 
            .I2(rx_data[0]), .I3(\data_in_frame[23] [0]), .O(n29699));
    defparam i15691_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i49854_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65276));   // verilog/coms.v(158[12:15])
    defparam i49854_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49855_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65277));   // verilog/coms.v(158[12:15])
    defparam i49855_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16011_3_lut_4_lut (.I0(n8_adj_14), .I1(n57041), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n30019));
    defparam i16011_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16008_3_lut_4_lut (.I0(n8_adj_14), .I1(n57041), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n30016));
    defparam i16008_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16005_3_lut_4_lut (.I0(n8_adj_14), .I1(n57041), .I2(rx_data[5]), 
            .I3(\data_in_frame[6][5] ), .O(n30013));
    defparam i16005_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1747 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[9] [6]), .I3(GND_net), .O(n57587));
    defparam i1_2_lut_3_lut_adj_1747.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1748 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[11] [4]), 
            .I2(n10_adj_4824), .I3(n1130), .O(n26394));
    defparam i5_3_lut_4_lut_adj_1748.LUT_INIT = 16'h6996;
    SB_LUT4 i50130_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65279));   // verilog/coms.v(158[12:15])
    defparam i50130_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50018_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65282));   // verilog/coms.v(158[12:15])
    defparam i50018_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16002_3_lut_4_lut (.I0(n8_adj_14), .I1(n57041), .I2(rx_data[4]), 
            .I3(\data_in_frame[6][4] ), .O(n30010));
    defparam i16002_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15999_3_lut_4_lut (.I0(n8_adj_14), .I1(n57041), .I2(rx_data[3]), 
            .I3(\data_in_frame[6][3] ), .O(n30007));
    defparam i15999_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i50120_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65284));   // verilog/coms.v(158[12:15])
    defparam i50120_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15996_3_lut_4_lut (.I0(n8_adj_14), .I1(n57041), .I2(rx_data[2]), 
            .I3(\data_in_frame[6][2] ), .O(n30004));
    defparam i15996_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15993_3_lut_4_lut (.I0(n8_adj_14), .I1(n57041), .I2(rx_data[1]), 
            .I3(\data_in_frame[6][1] ), .O(n30001));
    defparam i15993_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i23217_3_lut (.I0(n43_adj_18), .I1(n375), .I2(n401), .I3(GND_net), 
            .O(n4_adj_19));
    defparam i23217_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i15990_3_lut_4_lut (.I0(n8_adj_14), .I1(n57041), .I2(rx_data[0]), 
            .I3(\data_in_frame[6][0] ), .O(n29998));
    defparam i15990_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n69276_bdd_4_lut (.I0(n69276), .I1(n62808), .I2(n62807), .I3(\byte_transmit_counter[2] ), 
            .O(n69279));
    defparam n69276_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i49921_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65286));   // verilog/coms.v(158[12:15])
    defparam i49921_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50128_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65290));   // verilog/coms.v(158[12:15])
    defparam i50128_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16029_3_lut_4_lut (.I0(n28415), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n30037));
    defparam i16029_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16026_3_lut_4_lut (.I0(n28415), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n30034));
    defparam i16026_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16023_3_lut_4_lut (.I0(n28415), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n30031));
    defparam i16023_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1749 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [6]), 
            .I2(\data_out_frame[7] [2]), .I3(\data_out_frame[5] [1]), .O(n26083));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_4_lut_adj_1749.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1750 (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[7] [0]), 
            .I2(\data_out_frame[4] [6]), .I3(GND_net), .O(n57744));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_4_lut_adj_1750.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_2_i2_3_lut (.I0(\data_out_frame[0][2] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_4957));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_2_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i50663_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65297));   // verilog/coms.v(158[12:15])
    defparam i50663_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16020_3_lut_4_lut (.I0(n28415), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n30028));
    defparam i16020_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16017_3_lut_4_lut (.I0(n28415), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n30025));
    defparam i16017_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16113_3_lut_4_lut (.I0(n8_adj_16), .I1(n57037), .I2(rx_data[7]), 
            .I3(\data_in_frame[10][7] ), .O(n30121));
    defparam i16113_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i49964_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65307));   // verilog/coms.v(158[12:15])
    defparam i49964_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16110_3_lut_4_lut (.I0(n8_adj_16), .I1(n57037), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n30118));
    defparam i16110_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16106_3_lut_4_lut (.I0(n8_adj_16), .I1(n57037), .I2(rx_data[5]), 
            .I3(\data_in_frame[10][5] ), .O(n30114));
    defparam i16106_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i49987_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65311));   // verilog/coms.v(158[12:15])
    defparam i49987_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49992_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65312));   // verilog/coms.v(158[12:15])
    defparam i49992_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16103_3_lut_4_lut (.I0(n8_adj_16), .I1(n57037), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n30111));
    defparam i16103_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16100_3_lut_4_lut (.I0(n8_adj_16), .I1(n57037), .I2(rx_data[3]), 
            .I3(\data_in_frame[10][3] ), .O(n30108));
    defparam i16100_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53569 (.I0(\byte_transmit_counter[1] ), 
            .I1(n62789), .I2(n62790), .I3(\byte_transmit_counter[2] ), 
            .O(n69264));
    defparam byte_transmit_counter_1__bdd_4_lut_53569.LUT_INIT = 16'he4aa;
    SB_LUT4 n69264_bdd_4_lut (.I0(n69264), .I1(n62787), .I2(n62786), .I3(\byte_transmit_counter[2] ), 
            .O(n69267));
    defparam n69264_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_3_lut_4_lut_adj_1751 (.I0(\data_out_frame[4] [0]), .I1(n57090), 
            .I2(\data_out_frame[6] [6]), .I3(n1130), .O(n14_adj_4820));   // verilog/coms.v(100[12:26])
    defparam i5_3_lut_4_lut_adj_1751.LUT_INIT = 16'h6996;
    SB_LUT4 i16097_3_lut_4_lut (.I0(n8_adj_16), .I1(n57037), .I2(rx_data[2]), 
            .I3(\data_in_frame[10][2] ), .O(n30105));
    defparam i16097_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i49998_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65313));   // verilog/coms.v(158[12:15])
    defparam i49998_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16094_3_lut_4_lut (.I0(n8_adj_16), .I1(n57037), .I2(rx_data[1]), 
            .I3(\data_in_frame[10][1] ), .O(n30102));
    defparam i16094_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53560 (.I0(\byte_transmit_counter[1] ), 
            .I1(n62726), .I2(n62727), .I3(\byte_transmit_counter[2] ), 
            .O(n69258));
    defparam byte_transmit_counter_1__bdd_4_lut_53560.LUT_INIT = 16'he4aa;
    SB_LUT4 n69258_bdd_4_lut (.I0(n69258), .I1(n62715), .I2(n62714), .I3(\byte_transmit_counter[2] ), 
            .O(n69261));
    defparam n69258_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53555 (.I0(\byte_transmit_counter[1] ), 
            .I1(\data_out_frame[21] [5]), .I2(\data_out_frame[23] [5]), 
            .I3(\byte_transmit_counter[0] ), .O(n69252));
    defparam byte_transmit_counter_1__bdd_4_lut_53555.LUT_INIT = 16'he4aa;
    SB_LUT4 i16090_3_lut_4_lut (.I0(n8_adj_16), .I1(n57037), .I2(rx_data[0]), 
            .I3(\data_in_frame[10]_c [0]), .O(n30098));
    defparam i16090_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n69252_bdd_4_lut (.I0(n69252), .I1(\data_out_frame[22] [5]), 
            .I2(\data_out_frame[20] [5]), .I3(\byte_transmit_counter[0] ), 
            .O(n69255));
    defparam n69252_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i50655_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65355));   // verilog/coms.v(158[12:15])
    defparam i50655_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_2_lut_3_lut_adj_1752 (.I0(\data_out_frame[9] [1]), .I1(n26423), 
            .I2(\data_out_frame[11] [2]), .I3(GND_net), .O(n10_adj_4818));   // verilog/coms.v(88[17:28])
    defparam i2_2_lut_3_lut_adj_1752.LUT_INIT = 16'h9696;
    SB_LUT4 i50089_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65359));   // verilog/coms.v(158[12:15])
    defparam i50089_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16138_3_lut_4_lut (.I0(n28399), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n30146));
    defparam i16138_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i50092_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65360));   // verilog/coms.v(158[12:15])
    defparam i50092_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16134_3_lut_4_lut (.I0(n28399), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n30142));
    defparam i16134_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i50093_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65361));   // verilog/coms.v(158[12:15])
    defparam i50093_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50094_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65362));   // verilog/coms.v(158[12:15])
    defparam i50094_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i50116_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n65365));   // verilog/coms.v(158[12:15])
    defparam i50116_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16131_3_lut_4_lut (.I0(n28399), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n30139));
    defparam i16131_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53550 (.I0(\byte_transmit_counter[1] ), 
            .I1(n62708), .I2(n62709), .I3(\byte_transmit_counter[2] ), 
            .O(n69246));
    defparam byte_transmit_counter_1__bdd_4_lut_53550.LUT_INIT = 16'he4aa;
    SB_LUT4 n69246_bdd_4_lut (.I0(n69246), .I1(n62868), .I2(n62867), .I3(\byte_transmit_counter[2] ), 
            .O(n69249));
    defparam n69246_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16128_3_lut_4_lut (.I0(n28399), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n30136));
    defparam i16128_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53588 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n69240));
    defparam byte_transmit_counter_0__bdd_4_lut_53588.LUT_INIT = 16'he4aa;
    SB_LUT4 n69240_bdd_4_lut (.I0(n69240), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n69243));
    defparam n69240_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1753 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[8] [5]), 
            .I2(\data_out_frame[8] [4]), .I3(GND_net), .O(n57052));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1753.LUT_INIT = 16'h9696;
    SB_LUT4 i14367_1_lut (.I0(n3470), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n28374));   // verilog/coms.v(148[4] 304[11])
    defparam i14367_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52638_3_lut_4_lut (.I0(n28399), .I1(reset), .I2(\data_in_frame[11] [3]), 
            .I3(rx_data[3]), .O(n56283));
    defparam i52638_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i52637_3_lut_4_lut (.I0(n28399), .I1(reset), .I2(\data_in_frame[11] [2]), 
            .I3(rx_data[2]), .O(n56273));
    defparam i52637_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(n62818), .I2(n62815), .I3(byte_transmit_counter[3]), .O(n69234));
    defparam byte_transmit_counter_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i52636_3_lut_4_lut (.I0(n28399), .I1(reset), .I2(\data_in_frame[11] [1]), 
            .I3(rx_data[1]), .O(n56257));
    defparam i52636_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 n69234_bdd_4_lut (.I0(n69234), .I1(n62730), .I2(n62729), .I3(byte_transmit_counter[3]), 
            .O(n69237));
    defparam n69234_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i50280_2_lut_3_lut (.I0(\FRAME_MATCHER.i[5] ), .I1(n8), .I2(n130), 
            .I3(GND_net), .O(n65432));
    defparam i50280_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i2_3_lut_4_lut_adj_1754 (.I0(\data_out_frame[7] [3]), .I1(n57516), 
            .I2(\data_out_frame[9] [4]), .I3(n26083), .O(n57265));
    defparam i2_3_lut_4_lut_adj_1754.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53540 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n69228));
    defparam byte_transmit_counter_0__bdd_4_lut_53540.LUT_INIT = 16'he4aa;
    SB_LUT4 n69228_bdd_4_lut (.I0(n69228), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n69231));
    defparam n69228_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1755 (.I0(\data_out_frame[9] [5]), .I1(\data_out_frame[7] [3]), 
            .I2(n57516), .I3(GND_net), .O(n57185));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1755.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53531 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(\byte_transmit_counter[1] ), .O(n69222));
    defparam byte_transmit_counter_0__bdd_4_lut_53531.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1756 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[4] [0]), 
            .I2(\data_out_frame[8] [4]), .I3(\data_out_frame[5] [7]), .O(n57596));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_4_lut_adj_1756.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1757 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[1] [1]), .I3(n25906), .O(n4_adj_5021));
    defparam i1_2_lut_3_lut_4_lut_adj_1757.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1758 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[1] [1]), .I3(n25797), .O(n62190));
    defparam i1_2_lut_3_lut_4_lut_adj_1758.LUT_INIT = 16'h6996;
    SB_LUT4 n69222_bdd_4_lut (.I0(n69222), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(\byte_transmit_counter[1] ), 
            .O(n69225));
    defparam n69222_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1759 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[1] [1]), .I3(n57732), .O(n62256));
    defparam i1_2_lut_3_lut_4_lut_adj_1759.LUT_INIT = 16'h6996;
    SB_LUT4 i15647_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57046), 
            .I2(rx_data[7]), .I3(\data_in_frame[21] [7]), .O(n29655));
    defparam i15647_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15643_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57046), 
            .I2(rx_data[6]), .I3(\data_in_frame[21] [6]), .O(n29651));
    defparam i15643_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15624_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57046), 
            .I2(rx_data[5]), .I3(\data_in_frame[21] [5]), .O(n29632));
    defparam i15624_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1760 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[0] [4]), 
            .I2(n57115), .I3(\data_in_frame[7] [1]), .O(n6_adj_5022));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1760.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53526 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(\byte_transmit_counter[1] ), .O(n69216));
    defparam byte_transmit_counter_0__bdd_4_lut_53526.LUT_INIT = 16'he4aa;
    SB_LUT4 n69216_bdd_4_lut (.I0(n69216), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n69219));
    defparam n69216_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53545 (.I0(\byte_transmit_counter[1] ), 
            .I1(n62723), .I2(n62724), .I3(\byte_transmit_counter[2] ), 
            .O(n69210));
    defparam byte_transmit_counter_1__bdd_4_lut_53545.LUT_INIT = 16'he4aa;
    SB_LUT4 n69210_bdd_4_lut (.I0(n69210), .I1(n62721), .I2(n62720), .I3(\byte_transmit_counter[2] ), 
            .O(n69213));
    defparam n69210_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53516 (.I0(\byte_transmit_counter[1] ), 
            .I1(n62801), .I2(n62802), .I3(\byte_transmit_counter[2] ), 
            .O(n69204));
    defparam byte_transmit_counter_1__bdd_4_lut_53516.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1761 (.I0(\data_out_frame[13] [5]), .I1(n25095), 
            .I2(\data_out_frame[15] [6]), .I3(GND_net), .O(n57560));
    defparam i1_2_lut_3_lut_adj_1761.LUT_INIT = 16'h9696;
    SB_LUT4 n69204_bdd_4_lut (.I0(n69204), .I1(n62799), .I2(n62798), .I3(\byte_transmit_counter[2] ), 
            .O(n69207));
    defparam n69204_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53511 (.I0(\byte_transmit_counter[1] ), 
            .I1(n62768), .I2(n62769), .I3(\byte_transmit_counter[2] ), 
            .O(n69198));
    defparam byte_transmit_counter_1__bdd_4_lut_53511.LUT_INIT = 16'he4aa;
    SB_LUT4 i15621_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57046), 
            .I2(rx_data[4]), .I3(\data_in_frame[21] [4]), .O(n29629));
    defparam i15621_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n69198_bdd_4_lut (.I0(n69198), .I1(n62820), .I2(n62819), .I3(\byte_transmit_counter[2] ), 
            .O(n69201));
    defparam n69198_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i52651_2_lut_3_lut (.I0(n51753), .I1(\data_out_frame[18] [7]), 
            .I2(\data_out_frame[18] [6]), .I3(GND_net), .O(n68337));
    defparam i52651_2_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53521 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n69192));
    defparam byte_transmit_counter_0__bdd_4_lut_53521.LUT_INIT = 16'he4aa;
    SB_LUT4 n69192_bdd_4_lut (.I0(n69192), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n69195));
    defparam n69192_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15613_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57046), 
            .I2(rx_data[3]), .I3(\data_in_frame[21] [3]), .O(n29621));
    defparam i15613_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53506 (.I0(\byte_transmit_counter[1] ), 
            .I1(n62705), .I2(n62706), .I3(\byte_transmit_counter[2] ), 
            .O(n69186));
    defparam byte_transmit_counter_1__bdd_4_lut_53506.LUT_INIT = 16'he4aa;
    SB_LUT4 n69186_bdd_4_lut (.I0(n69186), .I1(n62832), .I2(n62831), .I3(\byte_transmit_counter[2] ), 
            .O(n69189));
    defparam n69186_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15610_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57046), 
            .I2(rx_data[2]), .I3(\data_in_frame[21] [2]), .O(n29618));
    defparam i15610_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1762 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[15] [5]), 
            .I2(n26257), .I3(n51676), .O(n52737));
    defparam i1_2_lut_4_lut_adj_1762.LUT_INIT = 16'h6996;
    SB_LUT4 i15606_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57046), 
            .I2(rx_data[1]), .I3(\data_in_frame[21] [1]), .O(n29614));
    defparam i15606_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53497 (.I0(\byte_transmit_counter[1] ), 
            .I1(n62624), .I2(n62625), .I3(\byte_transmit_counter[2] ), 
            .O(n69180));
    defparam byte_transmit_counter_1__bdd_4_lut_53497.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_53756 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n69486));
    defparam byte_transmit_counter_0__bdd_4_lut_53756.LUT_INIT = 16'he4aa;
    SB_LUT4 n69486_bdd_4_lut (.I0(n69486), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n69489));
    defparam n69486_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1763 (.I0(\data_out_frame[17] [2]), .I1(\data_out_frame[15] [1]), 
            .I2(\data_out_frame[15] [0]), .I3(n51656), .O(n57671));
    defparam i2_3_lut_4_lut_adj_1763.LUT_INIT = 16'h6996;
    SB_LUT4 n69180_bdd_4_lut (.I0(n69180), .I1(n62856), .I2(n62855), .I3(\byte_transmit_counter[2] ), 
            .O(n69183));
    defparam n69180_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1764 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[16] [7]), 
            .I2(\data_out_frame[19] [2]), .I3(GND_net), .O(n26626));
    defparam i1_2_lut_3_lut_adj_1764.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53492 (.I0(\byte_transmit_counter[1] ), 
            .I1(n62711), .I2(n62712), .I3(\byte_transmit_counter[2] ), 
            .O(n69174));
    defparam byte_transmit_counter_1__bdd_4_lut_53492.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1765 (.I0(\data_out_frame[22] [4]), .I1(n51837), 
            .I2(n23709), .I3(GND_net), .O(n8_adj_4797));
    defparam i1_2_lut_3_lut_adj_1765.LUT_INIT = 16'h9696;
    SB_LUT4 n69174_bdd_4_lut (.I0(n69174), .I1(n62859), .I2(n62858), .I3(\byte_transmit_counter[2] ), 
            .O(n69177));
    defparam n69174_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1766 (.I0(n23668), .I1(\data_out_frame[20] [1]), 
            .I2(\data_out_frame[20] [3]), .I3(n59054), .O(n52618));
    defparam i2_3_lut_4_lut_adj_1766.LUT_INIT = 16'h9669;
    SB_LUT4 i15601_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n57046), 
            .I2(rx_data[0]), .I3(\data_in_frame[21] [0]), .O(n29609));
    defparam i15601_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1767 (.I0(\data_out_frame[17] [4]), .I1(\data_out_frame[15] [3]), 
            .I2(\data_out_frame[15] [2]), .I3(n51656), .O(n57590));
    defparam i2_3_lut_4_lut_adj_1767.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1768 (.I0(DE_c), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(n6_adj_4858), .I3(\FRAME_MATCHER.i_31__N_2512 ), .O(n26912));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1768.LUT_INIT = 16'haaa8;
    SB_LUT4 i1_2_lut_4_lut_adj_1769 (.I0(\data_out_frame[13] [6]), .I1(\data_out_frame[11] [5]), 
            .I2(n51541), .I3(n26394), .O(n57422));
    defparam i1_2_lut_4_lut_adj_1769.LUT_INIT = 16'h6996;
    SB_LUT4 select_777_Select_60_i2_4_lut (.I0(\data_out_frame[7] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder0_position_scaled[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5038));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_60_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1770 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n25483), .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n62408));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_4_lut_adj_1770.LUT_INIT = 16'hfff4;
    SB_LUT4 i2_3_lut_4_lut_adj_1771 (.I0(n59193), .I1(n51364), .I2(\data_out_frame[18] [4]), 
            .I3(\data_out_frame[18] [3]), .O(n52767));
    defparam i2_3_lut_4_lut_adj_1771.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1772 (.I0(\data_out_frame[20] [0]), .I1(n59193), 
            .I2(\data_out_frame[18] [4]), .I3(GND_net), .O(n6_c));
    defparam i1_2_lut_3_lut_adj_1772.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_53487 (.I0(\byte_transmit_counter[1] ), 
            .I1(n62843), .I2(n62844), .I3(\byte_transmit_counter[2] ), 
            .O(n69168));
    defparam byte_transmit_counter_1__bdd_4_lut_53487.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1773 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[20] [7]), .I3(GND_net), .O(n57232));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_3_lut_adj_1773.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1774 (.I0(n52677), .I1(n57450), .I2(\data_out_frame[16] [1]), 
            .I3(\data_out_frame[16] [2]), .O(n51364));
    defparam i2_3_lut_4_lut_adj_1774.LUT_INIT = 16'h6996;
    SB_LUT4 n69168_bdd_4_lut (.I0(n69168), .I1(n62847), .I2(n62846), .I3(\byte_transmit_counter[2] ), 
            .O(n69171));
    defparam n69168_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1775 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(n51832), .I3(GND_net), .O(n52677));
    defparam i1_2_lut_3_lut_adj_1775.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1776 (.I0(\data_out_frame[18] [3]), .I1(n52677), 
            .I2(n57450), .I3(n26100), .O(n51745));
    defparam i1_2_lut_4_lut_adj_1776.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1777 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[18] [2]), 
            .I2(n10_adj_4773), .I3(\data_out_frame[16] [1]), .O(n52327));
    defparam i5_3_lut_4_lut_adj_1777.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1778 (.I0(n59521), .I1(n51640), .I2(\data_out_frame[21] [6]), 
            .I3(GND_net), .O(n57322));
    defparam i1_2_lut_3_lut_adj_1778.LUT_INIT = 16'h6969;
    SB_LUT4 i23231_3_lut_4_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10]_c [0]), 
            .I2(Kp_23__N_1748), .I3(n33761), .O(n29640));
    defparam i23231_3_lut_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i1_2_lut_3_lut_adj_1779 (.I0(\data_out_frame[21] [4]), .I1(n26626), 
            .I2(n57317), .I3(GND_net), .O(n8_adj_4769));
    defparam i1_2_lut_3_lut_adj_1779.LUT_INIT = 16'h9696;
    SB_LUT4 select_777_Select_212_i3_3_lut_4_lut (.I0(\data_out_frame[24] [2]), 
            .I1(n25158), .I2(\FRAME_MATCHER.state[3] ), .I3(n57487), .O(n3_adj_5026));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_212_i3_3_lut_4_lut.LUT_INIT = 16'h9060;
    SB_LUT4 i1_2_lut_4_lut_adj_1780 (.I0(\data_out_frame[24] [5]), .I1(n23668), 
            .I2(n57460), .I3(n59054), .O(n57395));
    defparam i1_2_lut_4_lut_adj_1780.LUT_INIT = 16'h9669;
    SB_LUT4 select_777_Select_223_i3_4_lut (.I0(n26374), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n57328), .I3(\data_out_frame[25] [6]), .O(n3_adj_5030));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_223_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i2_3_lut_4_lut_adj_1781 (.I0(n51654), .I1(n59466), .I2(\data_out_frame[21] [1]), 
            .I3(n25716), .O(n57626));
    defparam i2_3_lut_4_lut_adj_1781.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1782 (.I0(LED_c), .I1(n33769), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5103));   // verilog/TinyFPGA_B.v(4[10:13])
    defparam i1_2_lut_adj_1782.LUT_INIT = 16'heeee;
    SB_LUT4 i14903_4_lut (.I0(n2873), .I1(n23_adj_5103), .I2(n27274), 
            .I3(\FRAME_MATCHER.i_31__N_2513 ), .O(n28911));   // verilog/coms.v(130[12] 305[6])
    defparam i14903_4_lut.LUT_INIT = 16'ha8a0;
    SB_LUT4 i2_3_lut_4_lut_adj_1783 (.I0(n57350), .I1(\data_out_frame[23] [2]), 
            .I2(\data_out_frame[23] [3]), .I3(n59922), .O(n25071));
    defparam i2_3_lut_4_lut_adj_1783.LUT_INIT = 16'h9669;
    SB_LUT4 i19758_4_lut (.I0(Kp_23__N_1748), .I1(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(LED_c), .O(n33766));   // verilog/coms.v(118[11:12])
    defparam i19758_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i1_2_lut_4_lut_adj_1784 (.I0(\data_out_frame[20] [5]), .I1(n57065), 
            .I2(n57412), .I3(n51784), .O(n9));
    defparam i1_2_lut_4_lut_adj_1784.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1785 (.I0(n33766), .I1(n27696), .I2(GND_net), 
            .I3(GND_net), .O(n5));
    defparam i1_2_lut_adj_1785.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_1786 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[16] [4]), 
            .I2(\data_out_frame[22] [7]), .I3(GND_net), .O(n57377));
    defparam i1_2_lut_3_lut_adj_1786.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1787 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[7] [3]), 
            .I2(encoder0_position_scaled[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5029));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1787.LUT_INIT = 16'ha088;
    SB_LUT4 select_777_Select_221_i3_3_lut_4_lut (.I0(\data_out_frame[25] [3]), 
            .I1(n51598), .I2(\FRAME_MATCHER.state[3] ), .I3(n57484), .O(n3_adj_5028));   // verilog/coms.v(148[4] 304[11])
    defparam select_777_Select_221_i3_3_lut_4_lut.LUT_INIT = 16'h9060;
    SB_LUT4 i1_2_lut_4_lut_adj_1788 (.I0(\data_out_frame[25] [4]), .I1(n57350), 
            .I2(n57659), .I3(n59922), .O(n57484));
    defparam i1_2_lut_4_lut_adj_1788.LUT_INIT = 16'h9669;
    SB_LUT4 select_1650_Select_0_i1_2_lut (.I0(tx_transmit_N_3416), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n1));   // verilog/coms.v(148[4] 304[11])
    defparam select_1650_Select_0_i1_2_lut.LUT_INIT = 16'h8888;
    uart_tx tx (.\r_SM_Main_2__N_3536[1] (r_SM_Main_2__N_3536[1]), .r_SM_Main({r_SM_Main}), 
            .GND_net(GND_net), .n57935(n57935), .n58550(n58550), .\r_SM_Main_2__N_3545[0] (r_SM_Main_2__N_3545[0]), 
            .n6(n6), .tx_o(tx_o), .clk16MHz(clk16MHz), .tx_data({tx_data}), 
            .n29661(n29661), .tx_active(tx_active), .r_Clock_Count({r_Clock_Count}), 
            .VCC_net(VCC_net), .n4940(n4940), .n29(n29_adj_5105), .n23(n23_adj_5106), 
            .\o_Rx_DV_N_3488[12] (o_Rx_DV_N_3488[12]), .\o_Rx_DV_N_3488[24] (o_Rx_DV_N_3488[24]), 
            .n27(n27), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(110[25:94])
    uart_rx rx (.\r_Bit_Index[0] (\r_Bit_Index[0] ), .GND_net(GND_net), 
            .\o_Rx_DV_N_3488[12] (o_Rx_DV_N_3488[12]), .n4937(n4937), .\o_Rx_DV_N_3488[8] (\o_Rx_DV_N_3488[8] ), 
            .\o_Rx_DV_N_3488[24] (o_Rx_DV_N_3488[24]), .n29(n29_adj_5105), 
            .n23(n23_adj_5106), .n60724(n60724), .baudrate({baudrate}), 
            .n4940(n4940), .\r_SM_Main[0] (r_SM_Main[0]), .n27(n27), .n58550(n58550), 
            .VCC_net(VCC_net), .clk16MHz(clk16MHz), .\r_SM_Main[2] (\r_SM_Main[2]_adj_20 ), 
            .n25530(n25530), .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), .\r_SM_Main[1] (\r_SM_Main[1]_adj_21 ), 
            .n27966(n27966), .n56959(n56959), .n60740(n60740), .n29884(n29884), 
            .rx_data({rx_data}), .n60788(n60788), .n60756(n60756), .n29866(n29866), 
            .\o_Rx_DV_N_3488[7] (\o_Rx_DV_N_3488[7] ), .\o_Rx_DV_N_3488[6] (\o_Rx_DV_N_3488[6] ), 
            .\o_Rx_DV_N_3488[5] (\o_Rx_DV_N_3488[5] ), .\o_Rx_DV_N_3488[4] (\o_Rx_DV_N_3488[4] ), 
            .\o_Rx_DV_N_3488[3] (\o_Rx_DV_N_3488[3] ), .\o_Rx_DV_N_3488[2] (\o_Rx_DV_N_3488[2] ), 
            .\o_Rx_DV_N_3488[1] (\o_Rx_DV_N_3488[1] ), .\o_Rx_DV_N_3488[0] (\o_Rx_DV_N_3488[0] ), 
            .n29774(n29774), .n29773(n29773), .n29772(n29772), .r_Clock_Count({r_Clock_Count_adj_30}), 
            .n58000(n58000), .n30502(n30502), .n52851(n52851), .rx_data_ready(rx_data_ready), 
            .n30498(n30498), .n30201(n30201), .n30200(n30200), .\r_SM_Main_2__N_3536[1] (r_SM_Main_2__N_3536[1]), 
            .n60708(n60708), .n60692(n60692), .n60804(n60804), .n27724(n27724), 
            .n60772(n60772)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(96[25:68])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (\r_SM_Main_2__N_3536[1] , r_SM_Main, GND_net, n57935, 
            n58550, \r_SM_Main_2__N_3545[0] , n6, tx_o, clk16MHz, 
            tx_data, n29661, tx_active, r_Clock_Count, VCC_net, n4940, 
            n29, n23, \o_Rx_DV_N_3488[12] , \o_Rx_DV_N_3488[24] , n27, 
            tx_enable) /* synthesis syn_module_defined=1 */ ;
    input \r_SM_Main_2__N_3536[1] ;
    output [2:0]r_SM_Main;
    input GND_net;
    input n57935;
    input n58550;
    input \r_SM_Main_2__N_3545[0] ;
    output n6;
    output tx_o;
    input clk16MHz;
    input [7:0]tx_data;
    input n29661;
    output tx_active;
    output [8:0]r_Clock_Count;
    input VCC_net;
    input n4940;
    input n29;
    input n23;
    input \o_Rx_DV_N_3488[12] ;
    input \o_Rx_DV_N_3488[24] ;
    input n27;
    output tx_enable;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n58521, n56768, n29192;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(34[16:27])
    wire [2:0]n460;
    
    wire n3, n40591, n25035;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(35[16:25])
    
    wire n52883, n65301;
    wire [8:0]n41;
    
    wire n50554, n50553, n50552, n50551, n50550, n50549, n50548, 
        n50547, n58022, n40563, n52881, n69552, n3_adj_4725, n60522, 
        n60528, n65295, n65292, n9, n69297, n14, n15, n62837, 
        n62838, n62871, n62870, n69294;
    
    SB_LUT4 i42167_rep_29_2_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(GND_net), .I3(GND_net), .O(n58521));
    defparam i42167_rep_29_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(n57935), .I1(n58521), .I2(r_SM_Main[1]), .I3(n56768), 
            .O(n29192));
    defparam i1_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i16_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n460[1]));   // verilog/uart_tx.v(34[16:27])
    defparam i16_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i17_4_lut (.I0(r_SM_Main[0]), .I1(n58550), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n6));
    defparam i17_4_lut.LUT_INIT = 16'h3530;
    SB_DFFE o_Tx_Serial_51 (.Q(tx_o), .C(clk16MHz), .E(n40591), .D(n3));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk16MHz), .E(n25035), 
            .D(tx_data[0]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n52883), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i50684_2_lut_3_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n65301));   // verilog/uart_tx.v(32[16:25])
    defparam i50684_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_DFF r_Tx_Active_53 (.Q(tx_active), .C(clk16MHz), .D(n29661));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 r_Clock_Count_1953_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n50554), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1953_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1953_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n50553), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1953_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1953_add_4_9 (.CI(n50553), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n50554));
    SB_LUT4 r_Clock_Count_1953_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n50552), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1953_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1953_add_4_8 (.CI(n50552), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n50553));
    SB_LUT4 r_Clock_Count_1953_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n50551), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1953_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1953_add_4_7 (.CI(n50551), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n50552));
    SB_LUT4 r_Clock_Count_1953_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n50550), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1953_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1953_add_4_6 (.CI(n50550), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n50551));
    SB_LUT4 r_Clock_Count_1953_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n50549), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1953_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1953_add_4_5 (.CI(n50549), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n50550));
    SB_LUT4 r_Clock_Count_1953_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n50548), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1953_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1953_add_4_4 (.CI(n50548), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n50549));
    SB_LUT4 r_Clock_Count_1953_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n50547), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1953_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1953_add_4_3 (.CI(n50547), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n50548));
    SB_LUT4 r_Clock_Count_1953_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1953_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1953_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n50547));
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n58022), 
            .D(n460[1]), .R(n29192));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n58022), 
            .D(n460[2]), .R(n29192));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Clock_Count_1953__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n40591), .D(n41[1]), .R(n40563));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1953__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n40591), .D(n41[2]), .R(n40563));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1953__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n40591), .D(n41[3]), .R(n40563));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1953__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n40591), .D(n41[4]), .R(n40563));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1953__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n40591), .D(n41[5]), .R(n40563));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1953__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n40591), .D(n41[6]), .R(n40563));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1953__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n40591), .D(n41[7]), .R(n40563));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1953__i8 (.Q(r_Clock_Count[8]), .C(clk16MHz), 
            .E(n40591), .D(n41[8]), .R(n40563));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_1953__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n40591), .D(n41[0]), .R(n40563));   // verilog/uart_tx.v(119[34:51])
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk16MHz), .E(VCC_net), 
            .D(n52881));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n69552));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3_adj_4725), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk16MHz), .E(n25035), 
            .D(tx_data[7]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk16MHz), .E(n25035), 
            .D(tx_data[6]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk16MHz), .E(n25035), 
            .D(tx_data[5]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk16MHz), .E(n25035), 
            .D(tx_data[4]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk16MHz), .E(n25035), 
            .D(tx_data[3]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk16MHz), .E(n25035), 
            .D(tx_data[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk16MHz), .E(n25035), 
            .D(tx_data[1]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i1_2_lut (.I0(n4940), .I1(r_SM_Main[0]), .I2(GND_net), .I3(GND_net), 
            .O(n60522));
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_adj_1089 (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3488[12] ), 
            .I3(n60522), .O(n60528));
    defparam i1_4_lut_adj_1089.LUT_INIT = 16'h0100;
    SB_LUT4 i10_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(r_SM_Main[1]), .I2(n27), 
            .I3(n60528), .O(n3_adj_4725));   // verilog/uart_tx.v(32[16:25])
    defparam i10_4_lut.LUT_INIT = 16'hc9cc;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(n56768));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i50659_3_lut (.I0(n56768), .I1(\o_Rx_DV_N_3488[12] ), .I2(n4940), 
            .I3(GND_net), .O(n65295));   // verilog/uart_tx.v(32[16:25])
    defparam i50659_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i50656_4_lut (.I0(n65295), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n65292));   // verilog/uart_tx.v(32[16:25])
    defparam i50656_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i23_4_lut (.I0(\r_SM_Main_2__N_3545[0] ), .I1(n65292), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n9));   // verilog/uart_tx.v(32[16:25])
    defparam i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_3_lut (.I0(n9), .I1(\r_SM_Main_2__N_3536[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n52883));   // verilog/uart_tx.v(32[16:25])
    defparam i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40591));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_SM_Main_2__I_0_62_i3_3_lut (.I0(r_SM_Main[0]), .I1(n69297), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(44[7] 143[14])
    defparam r_SM_Main_2__I_0_62_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[24] ), .I2(n27), 
            .I3(GND_net), .O(n14));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3488[12] ), .I2(n23), .I3(n4940), 
            .O(n15));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(n40591), .I2(n14), .I3(r_SM_Main[1]), 
            .O(n69552));
    defparam i8_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i47151_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n62837));
    defparam i47151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47152_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n62838));
    defparam i47152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47185_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n62871));
    defparam i47185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47184_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n62870));
    defparam i47184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n25035));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i12_4_lut (.I0(n65301), .I1(n58022), .I2(r_Bit_Index[0]), 
            .I3(n58521), .O(n52881));   // verilog/uart_tx.v(32[16:25])
    defparam i12_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 r_Bit_Index_2__bdd_4_lut (.I0(r_Bit_Index[2]), .I1(n62870), 
            .I2(n62871), .I3(r_Bit_Index[1]), .O(n69294));
    defparam r_Bit_Index_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n69294_bdd_4_lut (.I0(n69294), .I1(n62838), .I2(n62837), .I3(r_Bit_Index[1]), 
            .O(n69297));
    defparam n69294_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i53398_4_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n40563));
    defparam i53398_4_lut.LUT_INIT = 16'h1113;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(39[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53460_2_lut_4_lut (.I0(\r_SM_Main_2__N_3536[1] ), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[0]), .O(n58022));
    defparam i53460_2_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i26646_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n460[2]));   // verilog/uart_tx.v(34[16:27])
    defparam i26646_3_lut.LUT_INIT = 16'h6a6a;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (\r_Bit_Index[0] , GND_net, \o_Rx_DV_N_3488[12] , n4937, 
            \o_Rx_DV_N_3488[8] , \o_Rx_DV_N_3488[24] , n29, n23, n60724, 
            baudrate, n4940, \r_SM_Main[0] , n27, n58550, VCC_net, 
            clk16MHz, \r_SM_Main[2] , n25530, r_Rx_Data, RX_N_2, \r_SM_Main[1] , 
            n27966, n56959, n60740, n29884, rx_data, n60788, n60756, 
            n29866, \o_Rx_DV_N_3488[7] , \o_Rx_DV_N_3488[6] , \o_Rx_DV_N_3488[5] , 
            \o_Rx_DV_N_3488[4] , \o_Rx_DV_N_3488[3] , \o_Rx_DV_N_3488[2] , 
            \o_Rx_DV_N_3488[1] , \o_Rx_DV_N_3488[0] , n29774, n29773, 
            n29772, r_Clock_Count, n58000, n30502, n52851, rx_data_ready, 
            n30498, n30201, n30200, \r_SM_Main_2__N_3536[1] , n60708, 
            n60692, n60804, n27724, n60772) /* synthesis syn_module_defined=1 */ ;
    output \r_Bit_Index[0] ;
    input GND_net;
    output \o_Rx_DV_N_3488[12] ;
    input n4937;
    output \o_Rx_DV_N_3488[8] ;
    output \o_Rx_DV_N_3488[24] ;
    output n29;
    output n23;
    output n60724;
    input [31:0]baudrate;
    input n4940;
    input \r_SM_Main[0] ;
    output n27;
    output n58550;
    input VCC_net;
    input clk16MHz;
    output \r_SM_Main[2] ;
    output n25530;
    output r_Rx_Data;
    input RX_N_2;
    output \r_SM_Main[1] ;
    output n27966;
    input n56959;
    output n60740;
    input n29884;
    output [7:0]rx_data;
    output n60788;
    output n60756;
    input n29866;
    output \o_Rx_DV_N_3488[7] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[0] ;
    input n29774;
    input n29773;
    input n29772;
    output [7:0]r_Clock_Count;
    output n58000;
    input n30502;
    input n52851;
    output rx_data_ready;
    input n30498;
    input n30201;
    input n30200;
    output \r_SM_Main_2__N_3536[1] ;
    output n60708;
    output n60692;
    output n60804;
    output n27724;
    output n60772;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    wire [2:0]n479;
    
    wire n60712, n60718, n67986, n2713, n60328, n2845, n25622;
    wire [23:0]n294;
    
    wire n60382, n68298, n2827, n25644, n60330, n2957, n68310, 
        n2938, n60332, n3066, n1261;
    wire [23:0]n8035;
    
    wire n1408, n1266, n1413, n1262, n1409, n45, n49310, n1265, 
        n1412, n62574, n3;
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n39, n1264, n1411, n41, n49309, n60276, r_Rx_Data_R, 
        n1263, n1410, n43, n1267, n1414, n1415, n34, n67604, 
        n67605, n66138, n67021, n36, n38, n62610, n49308, n60376, 
        n66774, n67696, n1111;
    wire [23:0]n8009;
    
    wire n1115, n1112, n1113, n1114, n41_adj_4454, n49307;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n49306, n60374, n1116, n36_adj_4455, n38_adj_4456, n40, 
        n66151, n68083, n68084, n67909, n959, n58551, n44, n46, 
        n57842, n49305, n60372;
    wire [2:0]r_SM_Main_2__N_3446;
    
    wire n960, n11428, n20929, n20931, n49304, n961, n40_adj_4457, 
        n25545, n48, n962, n42, n43_adj_4458, n67391, n3046, n60334, 
        n3172, n49303, n60370, n38_adj_4459, n40_adj_4460, n42_adj_4461, 
        n66159, n68059, n68060, n49302, n60368, n25629, n49301, 
        n60274, n805, n42_adj_4462, n14, n15, n69533, n60728, 
        n60734, n60776, n60782, n803, n58597, n44_adj_4463, n46_adj_4464, 
        n57840, n61900, n804, n60744, n60750, n42863, n20919, 
        n20921, n61902, n61798, n61794, n61796, n61792, n61778, 
        n61676, n61790, n61666, n61658, n61656, n58123, n49300, 
        n60366, n42_adj_4465, n67626, n67627, n57838, n49299, n49298, 
        n49297, n49296, n62568, n62570, n25589, n65720, n48_adj_4466, 
        n68343, n44_adj_4467, n25632, n48_adj_4468, n42_adj_4469, 
        n67628, n67629, n48_adj_4470, n49295, n49294, n49293, n49292, 
        n49291, n49290, n49289, n49288, n49287, n59155, n25619, 
        n62318, n60908, n58609, n59474, n65325, n57899, n60962, 
        n65326, n61898, n60642, n62534, n60670, n62532, n62472, 
        n62450, n62602, n62592, n65714, n60990, n61804, n61748, 
        n61744, n61650, n61648, n61646, n60974, n60966, n61806, 
        n65404, n46_adj_4471, n60292, n61644, n62486, n42865, n60294, 
        n62504, n60252, n62556, n62540, n60586, n60604, n62604, 
        n3155;
    wire [23:0]n8425;
    
    wire n39_adj_4472, n3154, n41_adj_4473, n3158, n33, n3157, n35, 
        n3156, n37, n3163, n23_adj_4474, n3162, n25, n3160, n29_adj_4475, 
        n3159, n31, n3171, n7, n3152, n45_adj_4476, n3153, n43_adj_4477, 
        n3170, n9, n3166, n17, n3165, n19, n3164, n21, n3169, 
        n11, n3168, n13, n4, n3167, n15_adj_4478, n3161, n27_adj_4479, 
        n65618, n65625, n16, n65596, n8, n24, n3274, n65636, 
        n66526, n66522, n67882, n67255, n68113, n12, n60336, n48_adj_4480, 
        n4_adj_4481, n67813, n67814, n65610, n10, n30, n65612, 
        n68169, n67754, n68295, n68296, n6, n67815, n67816, n65601, 
        n67397, n67752, n68234, n65603, n68001, n40_adj_4482, n60264, 
        n3151, n3253, n68003, n61746, n60272, n62448, n60826, 
        n60822, n60824, n60820, n62514, n62512, n62600;
    wire [23:0]n8399;
    
    wire n3047, n3048, n3049, n3063, n60830, n62572, n3050, n3053, 
        n33_adj_4483, n3054, n31_adj_4484, n3051, n37_adj_4485, n3052, 
        n35_adj_4486, n3058, n3059, n21_adj_4487, n23_adj_4488, n3057, 
        n3056, n25_adj_4489, n27_adj_4490, n3065, n9_adj_4491, n3055, 
        n3062, n3061, n13_adj_4492, n15_adj_4493, n17_adj_4494, n29_adj_4495, 
        n3060, n3064, n11_adj_4496, n19_adj_4497, n62546;
    wire [23:0]n8087;
    
    wire n48_adj_4498, n1702, n61904, n25552, n65669, n66629, n67303, 
        n67301, n65682, n6_adj_4499, n67821, n14_adj_4500, n32, 
        n67822, n65662, n12_adj_4501, n65660, n68167, n67744, n62350;
    wire [23:0]n8165;
    
    wire n48_adj_4502, n2110, n8_adj_4503, n67995, n67996;
    wire [7:0]n1;
    
    wire n50546, n50545, n50544, n65696, n66615, n10_adj_4507, n67393, 
        n67742, n67600, n68293, n67817, n68315, n68316, n50543, 
        n68306, n68107, n50542, n68108, n50541, n50540, n27767, 
        n29148;
    wire [23:0]n8373;
    
    wire n2946, n2939, n2940, n2941, n2944, n35_adj_4513, n2942, 
        n39_adj_4514, n2945, n33_adj_4515, n2943, n37_adj_4516, n2947, 
        n2948, n27_adj_4517, n29_adj_4518, n2949, n2950, n23_adj_4519, 
        n25_adj_4520, n2956, n3186, n50386, n3082, n50385, n3188, 
        n50384, n3084, n50383, n2977, n50382, n2867, n50381, n2754, 
        n50380, n2638, n50379, n2519, n50378, n2397, n50377, n11_adj_4521, 
        n2272, n50376, n2144, n50375, n2013, n50374, n1879, n50373, 
        n1742, n50372, n1602, n50371, n1459, n50370, n1460, n50369, 
        n1011, n50368, n856, n50367, n698, n50366, n858, n50365, 
        n538, n50364, n58062, n50363, n50362, n2955, n50361, n50360, 
        n50359, n50358, n50357, n50356, n50355, n50354, n50353, 
        n50352, n50351, n50350, n50349, n50348, n50347, n50346, 
        n50345, n50344, n50343, n58066, n50342, n50341, n50340, 
        n2951, n50339, n50338, n50337, n50336, n50335, n50334, 
        n50333, n50332, n50331, n50330, n50329, n2952, n50328, 
        n2953, n50327, n13_adj_4522, n2954, n50326, n50325, n50324, 
        n50323, n58070;
    wire [23:0]n8347;
    
    wire n50322, n21_adj_4523, n2828, n50321, n2829, n50320, n2830, 
        n50319, n2831, n50318, n2832, n50317, n15_adj_4524, n2833, 
        n50316, n17_adj_4525, n2834, n50315, n2835, n50314, n2836, 
        n50313, n19_adj_4526, n31_adj_4527, n2837, n50312, n2838, 
        n50311, n2839, n50310, n2840, n50309, n65742, n2841, n50308, 
        n2842, n50307, n2843, n50306, n2844, n50305, n50304, n58074;
    wire [23:0]n8321;
    
    wire n50303, n66669, n2714, n50302, n2715, n50301, n67323, 
        n67321, n65744, n2716, n50300, n2717, n50299, n2718, n50298, 
        n8_adj_4528, n2719, n50297, n67825, n67826, n2720, n50296, 
        n2721, n50295, n2722, n50294, n2723, n50293, n2724, n50292, 
        n2725, n50291, n2726, n50290, n2727, n50289, n2728, n50288, 
        n2729, n50287, n2730, n50286, n16_adj_4529, n34_adj_4530, 
        n58078;
    wire [23:0]n8295;
    
    wire n2596, n50285, n2597, n50284, n2598, n50283, n2599, n50282, 
        n2600, n50281, n2601, n50280, n2602, n50279, n2603, n50278, 
        n65734, n2604, n50277, n2605, n50276, n14_adj_4531, n65728, 
        n68165, n67738, n2606, n50275, n10_adj_4532, n67827, n67828, 
        n2607, n50274, n65757, n66657, n2608, n50273, n12_adj_4533, 
        n20, n2609, n50272, n2610, n50271, n2611, n50270, n26, 
        n2612, n50269, n67634, n68291, n60326, n58082;
    wire [23:0]n8269;
    
    wire n2476, n50268, n2477, n50267, n67389, n2478, n50266, 
        n2479, n50265, n2480, n50264, n2481, n50263, n2482, n50262, 
        n68317, n2483, n50261, n2484, n50260, n2485, n50259, n2486, 
        n50258, n2487, n50257, n2488, n50256, n2489, n50255, n2490, 
        n50254, n2491, n50253, n60324, n58086;
    wire [23:0]n8243;
    
    wire n2353, n50252, n2354, n50251, n2355, n50250, n2356, n50249, 
        n2357, n50248, n2358, n50247, n2359, n50246, n2360, n50245, 
        n2361, n50244, n2362, n50243, n2363, n50242, n2364, n50241, 
        n2365, n50240, n2366, n50239, n68318, n68304, n2367, n50238, 
        n60322, n58090;
    wire [23:0]n8217;
    
    wire n2227, n50237, n2228, n50236, n2229, n50235, n2230, n50234, 
        n2231, n50233, n37_adj_4534, n2232, n50232, n2233, n50231, 
        n2234, n50230, n2235, n50229, n41_adj_4535, n2236, n50228, 
        n2237, n50227, n2238, n50226, n2239, n50225, n2240, n50224, 
        n60320, n58094;
    wire [23:0]n8191;
    
    wire n2098, n50223, n2099, n50222, n2100, n50221, n2101, n50220, 
        n2102, n50219, n2103, n50218, n35_adj_4536, n2104, n50217, 
        n39_adj_4537, n29_adj_4538, n2105, n50216, n2106, n50215, 
        n2107, n50214, n2108, n50213, n60760, n31_adj_4539, n2109, 
        n50212, n1966, n50211, n1967, n50210, n1968, n50209, n1969, 
        n50208, n1970, n50207, n23_adj_4540, n1971, n50206, n1972, 
        n50205, n3_adj_4541, n1973, n50204, n25_adj_4542, n27_adj_4543, 
        n1974, n50203, n1975, n50202, n1976, n50201, n17_adj_4544, 
        n1977, n50200, n19_adj_4545;
    wire [23:0]n8139;
    
    wire n1831, n50199, n1832, n50198, n67903, n1693, n25639, 
        n1833, n50197, n1834, n50196, n1835, n50195, n1836, n50194, 
        n21_adj_4546, n1837, n50193, n33_adj_4547, n13_adj_4548, n1838, 
        n50192, n1839, n50191, n1840, n50190, n1841, n50189, n60318, 
        n58103;
    wire [23:0]n8113;
    
    wire n50188, n1694, n50187, n1695, n50186, n1696, n50185, 
        n1697, n50184, n1698, n50183, n1699, n50182, n15_adj_4549, 
        n65792, n1700, n50181, n1701, n50180, n1552, n50179, n66703, 
        n67337, n1553, n50178, n1554, n50177, n1555, n50176, n1556, 
        n50175, n1557, n50174, n1558, n50173, n1559, n50172, n1560, 
        n50171;
    wire [23:0]n8061;
    
    wire n50170, n50169, n50168, n50167, n50166, n50165, n50164, 
        n50163, n67335, n60316, n58112, n50162, n50161, n50160, 
        n50159, n50158, n65794, n50157, n50156, n60314, n58116, 
        n50155, n50154, n50153, n50152, n10_adj_4550, n50151, n67831, 
        n67832, n50150, n18, n36_adj_4551, n60312, n58120, n65788, 
        n16_adj_4552, n65786, n68163, n67732, n14_adj_4553, n22, 
        n61766, n12_adj_4554, n65800, n68161, n68162, n68046, n67646, 
        n68289, n67990, n68313, n68314, n30_adj_4555, n66094, n43_adj_4556, 
        n32_adj_4557, n37_adj_4558, n39_adj_4559, n41_adj_4560, n31_adj_4561, 
        n33_adj_4562, n25_adj_4563, n27_adj_4564, n29_adj_4565, n15_adj_4566, 
        n17_adj_4567, n19_adj_4568, n21_adj_4569, n23_adj_4570, n35_adj_4571, 
        n65849, n66763, n67361, n67357, n65853, n12_adj_4572, n67837, 
        n20_adj_4573, n38_adj_4574, n67838, n65841, n18_adj_4575, 
        n65834, n67835, n67724, n16_adj_4576, n24_adj_4577, n14_adj_4578, 
        n65861, n68159, n68160, n68048, n67674, n68150, n67988, 
        n68297, n65381, n56722, n65387, n65378, n65384, n45_adj_4579, 
        n39_adj_4580, n41_adj_4581, n33_adj_4582, n35_adj_4583, n27_adj_4584, 
        n29_adj_4585, n31_adj_4586, n43_adj_4587, n17_adj_4588, n19_adj_4589, 
        n21_adj_4590, n23_adj_4591, n25_adj_4592, n28, n66080, n37_adj_4593, 
        n65889, n66849, n67395, n67381, n65893, n14_adj_4594, n67843, 
        n67844, n22_adj_4595, n40_adj_4596, n65882, n20_adj_4597, 
        n65880, n67385, n67720, n18_adj_4598, n26_adj_4599, n16_adj_4600, 
        n65902, n68157, n68158, n68050, n67700, n67984, n30_adj_4601, 
        n67983, n37_adj_4602, n43_adj_4603, n39_adj_4604, n41_adj_4605, 
        n31_adj_4606, n33_adj_4607, n35_adj_4608, n27_adj_4609, n29_adj_4610, 
        n19_adj_4611, n21_adj_4612, n23_adj_4613, n25_adj_4614, n17_adj_4615, 
        n65947, n65941, n67767, n16_adj_4616, n67560, n67561, n65943, 
        n66859, n22_adj_4617, n67715, n66836, n60348, n20_adj_4618, 
        n28_adj_4619, n18_adj_4620, n65939, n68095, n68096, n67879, 
        n66861, n67874, n66834, n68185, n68186, n68188, n25607, 
        n28_adj_4621, n66064, n30_adj_4622, n60696, n60702, n60680, 
        n60686, n39_adj_4623, n45_adj_4624, n43_adj_4625, n48_adj_4626, 
        n33_adj_4627, n35_adj_4628, n37_adj_4629, n41_adj_4630, n29_adj_4631, 
        n31_adj_4632, n21_adj_4633, n23_adj_4634, n25_adj_4635, n27_adj_4636, 
        n19_adj_4637, n66005, n65999, n67773, n18_adj_4638, n67572, 
        n67573, n66003, n66879, n24_adj_4639, n26_adj_4640, n66830, 
        n22_adj_4641, n30_adj_4642, n20_adj_4643, n65992, n68093, 
        n68094, n67885, n66883, n67712, n66828, n67714, n41_adj_4644, 
        n39_adj_4645, n37_adj_4646, n35_adj_4647, n29_adj_4648, n31_adj_4649, 
        n33_adj_4650, n24_adj_4651, n23_adj_4652, n25_adj_4653, n27_adj_4654, 
        n21_adj_4655, n66044, n66030, n66026, n26_adj_4656, n20_adj_4657, 
        n26_adj_4658, n28_adj_4659, n24_adj_4660, n32_adj_4661, n22_adj_4662, 
        n66024, n68091, n68092, n67887, n67775, n66028, n68155, 
        n66824, n68241, n68242, n66052, n28_adj_4663, n68218, n43_adj_4664, 
        n41_adj_4665, n39_adj_4666, n37_adj_4667, n48_adj_4668, n31_adj_4669, 
        n33_adj_4670, n35_adj_4671, n25_adj_4672, n27_adj_4673, n29_adj_4674, 
        n23_adj_4675, n66054, n66046, n22_adj_4676, n30_adj_4677, 
        n34_adj_4678, n68089, n68090, n67891, n67779, n67972, n66818, 
        n68055, n68056, n60792, n60798, n35_adj_4679, n37_adj_4680, 
        n41_adj_4681, n39_adj_4682, n29_adj_4683, n31_adj_4684, n33_adj_4685, 
        n61800, n61750, n60848, n61808, n27_adj_4686, n60306, n66072, 
        n61386, n3_adj_4687, n38_adj_4688, n58097, n61390, n5, n26_adj_4689, 
        n67588, n61394, n8_adj_4690, n67589, n66066, n68087, n66804, 
        n68253, n68254, n58912, n37_adj_4691, n35_adj_4692, n41_adj_4693, 
        n29_adj_4694, n33_adj_4695, n31_adj_4696, n39_adj_4697, n27_adj_4698, 
        n66086, n38_adj_4699, n26_adj_4700, n67592, n67593, n66082, 
        n68085, n66792, n68251, n68252, n68194, n60440, n60446, 
        n62500, n62596, n2, n11645, n37_adj_4701, n39_adj_4702, 
        n43_adj_4703, n48_adj_4704, n41_adj_4705, n31_adj_4706, n33_adj_4707, 
        n35_adj_4708, n29_adj_4709, n66102, n40_adj_4710, n28_adj_4711, 
        n67594, n67595, n66098, n68057, n66790, n68281, n68282, 
        n43_adj_4712, n37_adj_4713, n41_adj_4714, n39_adj_4715, n61776, 
        n58106, n32_adj_4716, n67598, n67599, n66116, n67005, n34_adj_4717, 
        n67702, n66785, n67902, n37_adj_4718, n39_adj_4719, n43_adj_4720, 
        n41_adj_4721, n32_adj_4722, n67602, n67603, n66128, n67013, 
        n34_adj_4723, n67698, n66780, n67904, n67905, n6_adj_4724, 
        n65352, n65349, n60766, n60828, n60868, n60842, n60844, 
        n65372, n65369, n65366, n60400, n60406;
    
    SB_LUT4 i2162_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n479[2]));   // verilog/uart_rx.v(103[36:51])
    defparam i2162_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i2155_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n479[1]));   // verilog/uart_rx.v(103[36:51])
    defparam i2155_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4937), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n60712), .O(n60718));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_970 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n60718), .O(n60724));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_970.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut (.I0(n67986), .I1(baudrate[18]), .I2(n2713), 
            .I3(n60328), .O(n2845));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h7100;
    SB_LUT4 i53441_2_lut_4_lut (.I0(n67986), .I1(baudrate[18]), .I2(n2713), 
            .I3(n25622), .O(n294[5]));   // verilog/uart_rx.v(119[33:55])
    defparam i53441_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_4_lut_adj_971 (.I0(n23), .I1(\o_Rx_DV_N_3488[12] ), .I2(n4940), 
            .I3(\r_SM_Main[0] ), .O(n60382));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_971.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_972 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n27), .I2(n29), 
            .I3(n60382), .O(n58550));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_972.LUT_INIT = 16'hfffe;
    SB_LUT4 i53448_2_lut_4_lut (.I0(n68298), .I1(baudrate[19]), .I2(n2827), 
            .I3(n25644), .O(n294[4]));   // verilog/uart_rx.v(119[33:55])
    defparam i53448_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_973 (.I0(n68298), .I1(baudrate[19]), .I2(n2827), 
            .I3(n60330), .O(n2957));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_973.LUT_INIT = 16'h7100;
    SB_LUT4 i1_2_lut_4_lut_adj_974 (.I0(n68310), .I1(baudrate[20]), .I2(n2938), 
            .I3(n60332), .O(n3066));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_974.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_i942_3_lut (.I0(n1261), .I1(n8035[23]), .I2(n294[16]), 
            .I3(GND_net), .O(n1408));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i947_3_lut (.I0(n1266), .I1(n8035[18]), .I2(n294[16]), 
            .I3(GND_net), .O(n1413));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i943_3_lut (.I0(n1262), .I1(n8035[22]), .I2(n294[16]), 
            .I3(GND_net), .O(n1409));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i45_2_lut (.I0(n1409), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_38_add_2_26_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n49310), .O(\o_Rx_DV_N_3488[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i946_3_lut (.I0(n1265), .I1(n8035[19]), .I2(n294[16]), 
            .I3(GND_net), .O(n1412));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53451_2_lut_4_lut (.I0(n68310), .I1(baudrate[20]), .I2(n2938), 
            .I3(n62574), .O(n294[3]));   // verilog/uart_rx.v(119[33:55])
    defparam i53451_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n3), .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_965_i39_2_lut (.I0(n1412), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i945_3_lut (.I0(n1264), .I1(n8035[20]), .I2(n294[16]), 
            .I3(GND_net), .O(n1411));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i41_2_lut (.I0(n1411), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_38_add_2_25_lut (.I0(n60276), .I1(n25530), .I2(VCC_net), 
            .I3(n49309), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_DFF r_Rx_Data_56 (.Q(r_Rx_Data), .C(clk16MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(42[10] 46[8])
    SB_DFF r_Rx_Data_R_55 (.Q(r_Rx_Data_R), .C(clk16MHz), .D(RX_N_2));   // verilog/uart_rx.v(42[10] 46[8])
    SB_LUT4 div_37_i944_3_lut (.I0(n1263), .I1(n8035[21]), .I2(n294[16]), 
            .I3(GND_net), .O(n1410));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_965_i43_2_lut (.I0(n1410), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i948_3_lut (.I0(n1267), .I1(n8035[17]), .I2(n294[16]), 
            .I3(GND_net), .O(n1414));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_25 (.CI(n49309), .I0(n25530), .I1(VCC_net), 
            .CO(n49310));
    SB_LUT4 div_37_LessThan_965_i34_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1415), .I3(GND_net), .O(n34));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i34_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51918_3_lut (.I0(n34), .I1(baudrate[5]), .I2(n41), .I3(GND_net), 
            .O(n67604));   // verilog/uart_rx.v(119[33:55])
    defparam i51918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51919_3_lut (.I0(n67604), .I1(baudrate[6]), .I2(n43), .I3(GND_net), 
            .O(n67605));   // verilog/uart_rx.v(119[33:55])
    defparam i51919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51335_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n66138), 
            .O(n67021));
    defparam i51335_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_965_i38_3_lut (.I0(n36), .I1(baudrate[4]), .I2(n39), 
            .I3(GND_net), .O(n38));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_38_add_2_24_lut (.I0(n60376), .I1(n62610), .I2(VCC_net), 
            .I3(n49308), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i51088_3_lut (.I0(n67605), .I1(baudrate[7]), .I2(n45), .I3(GND_net), 
            .O(n66774));   // verilog/uart_rx.v(119[33:55])
    defparam i51088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52010_4_lut (.I0(n66774), .I1(n38), .I2(n45), .I3(n67021), 
            .O(n67696));   // verilog/uart_rx.v(119[33:55])
    defparam i52010_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY sub_38_add_2_24 (.CI(n49308), .I0(n62610), .I1(VCC_net), 
            .CO(n49309));
    SB_LUT4 div_37_i843_3_lut (.I0(n1111), .I1(n8009[23]), .I2(n294[17]), 
            .I3(GND_net), .O(n1261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i847_3_lut (.I0(n1115), .I1(n8009[19]), .I2(n294[17]), 
            .I3(GND_net), .O(n1265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i844_3_lut (.I0(n1112), .I1(n8009[22]), .I2(n294[17]), 
            .I3(GND_net), .O(n1262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i845_3_lut (.I0(n1113), .I1(n8009[21]), .I2(n294[17]), 
            .I3(GND_net), .O(n1263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i846_3_lut (.I0(n1114), .I1(n8009[20]), .I2(n294[17]), 
            .I3(GND_net), .O(n1264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i41_2_lut (.I0(n1264), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4454));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_38_add_2_23_lut (.I0(o_Rx_DV_N_3488[18]), .I1(n294[21]), 
            .I2(VCC_net), .I3(n49307), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_23 (.CI(n49307), .I0(n294[21]), .I1(VCC_net), 
            .CO(n49308));
    SB_LUT4 sub_38_add_2_22_lut (.I0(n60374), .I1(n294[20]), .I2(VCC_net), 
            .I3(n49306), .O(n60376)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_i848_3_lut (.I0(n1116), .I1(n8009[18]), .I2(n294[17]), 
            .I3(GND_net), .O(n1266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i36_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1267), .I3(GND_net), .O(n36_adj_4455));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i36_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_866_i40_3_lut (.I0(n38_adj_4456), .I1(baudrate[4]), 
            .I2(n41_adj_4454), .I3(GND_net), .O(n40));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52397_4_lut (.I0(n40), .I1(n36_adj_4455), .I2(n41_adj_4454), 
            .I3(n66151), .O(n68083));   // verilog/uart_rx.v(119[33:55])
    defparam i52397_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52398_3_lut (.I0(n68083), .I1(baudrate[5]), .I2(n1263), .I3(GND_net), 
            .O(n68084));   // verilog/uart_rx.v(119[33:55])
    defparam i52398_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52223_3_lut (.I0(n68084), .I1(baudrate[6]), .I2(n1262), .I3(GND_net), 
            .O(n67909));   // verilog/uart_rx.v(119[33:55])
    defparam i52223_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i5763_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n58551), .I3(n44), 
            .O(n46));   // verilog/uart_rx.v(119[33:55])
    defparam i5763_4_lut.LUT_INIT = 16'hb3a0;
    SB_CARRY sub_38_add_2_22 (.CI(n49306), .I0(n294[20]), .I1(VCC_net), 
            .CO(n49307));
    SB_LUT4 div_37_i742_4_lut (.I0(n57842), .I1(n294[18]), .I2(n46), .I3(baudrate[5]), 
            .O(n1111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i742_4_lut.LUT_INIT = 16'h9559;
    SB_LUT4 sub_38_add_2_21_lut (.I0(n60372), .I1(n294[19]), .I2(VCC_net), 
            .I3(n49305), .O(n60374)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_21 (.CI(n49305), .I0(n294[19]), .I1(VCC_net), 
            .CO(n49306));
    SB_LUT4 i52673_2_lut_3_lut_4_lut (.I0(r_SM_Main_2__N_3446[1]), .I1(\r_SM_Main[1] ), 
            .I2(r_SM_Main[0]), .I3(\r_SM_Main[2] ), .O(n27966));
    defparam i52673_2_lut_3_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i7244_4_lut (.I0(n960), .I1(n11428), .I2(n20929), .I3(baudrate[3]), 
            .O(n20931));   // verilog/uart_rx.v(119[33:55])
    defparam i7244_4_lut.LUT_INIT = 16'ha8aa;
    SB_LUT4 sub_38_add_2_20_lut (.I0(GND_net), .I1(n294[18]), .I2(VCC_net), 
            .I3(n49304), .O(o_Rx_DV_N_3488[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i743_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n294[18]), 
            .I3(n44), .O(n1112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i743_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i745_4_lut (.I0(n961), .I1(n40_adj_4457), .I2(n294[18]), 
            .I3(baudrate[2]), .O(n1114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i745_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i1_3_lut (.I0(n25545), .I1(n48), .I2(baudrate[0]), .I3(GND_net), 
            .O(n1116));
    defparam i1_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i5741_2_lut (.I0(n962), .I1(baudrate[1]), .I2(GND_net), .I3(GND_net), 
            .O(n40_adj_4457));   // verilog/uart_rx.v(119[33:55])
    defparam i5741_2_lut.LUT_INIT = 16'hbbbb;
    SB_CARRY sub_38_add_2_20 (.CI(n49304), .I0(n294[18]), .I1(VCC_net), 
            .CO(n49305));
    SB_LUT4 i7243_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), .I3(baudrate[1]), 
            .O(n20929));   // verilog/uart_rx.v(119[33:55])
    defparam i7243_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 div_37_i744_4_lut (.I0(n960), .I1(baudrate[3]), .I2(n294[18]), 
            .I3(n42), .O(n1113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i744_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_LessThan_765_i43_2_lut (.I0(n1113), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4458));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_975 (.I0(n67391), .I1(baudrate[21]), .I2(n3046), 
            .I3(n60334), .O(n3172));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_975.LUT_INIT = 16'h7100;
    SB_LUT4 sub_38_add_2_19_lut (.I0(n60370), .I1(n294[17]), .I2(VCC_net), 
            .I3(n49303), .O(n60372)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_19 (.CI(n49303), .I0(n294[17]), .I1(VCC_net), 
            .CO(n49304));
    SB_LUT4 div_37_LessThan_765_i38_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1116), .I3(GND_net), .O(n38_adj_4459));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i38_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_765_i42_3_lut (.I0(n40_adj_4460), .I1(baudrate[4]), 
            .I2(n43_adj_4458), .I3(GND_net), .O(n42_adj_4461));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i42_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52373_4_lut (.I0(n42_adj_4461), .I1(n38_adj_4459), .I2(n43_adj_4458), 
            .I3(n66159), .O(n68059));   // verilog/uart_rx.v(119[33:55])
    defparam i52373_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52374_3_lut (.I0(n68059), .I1(baudrate[5]), .I2(n1112), .I3(GND_net), 
            .O(n68060));   // verilog/uart_rx.v(119[33:55])
    defparam i52374_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 sub_38_add_2_18_lut (.I0(n60368), .I1(n294[16]), .I2(VCC_net), 
            .I3(n49302), .O(n60370)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i53456_2_lut_4_lut (.I0(n67391), .I1(baudrate[21]), .I2(n3046), 
            .I3(n25629), .O(n294[2]));   // verilog/uart_rx.v(119[33:55])
    defparam i53456_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_CARRY sub_38_add_2_18 (.CI(n49302), .I0(n294[16]), .I1(VCC_net), 
            .CO(n49303));
    SB_LUT4 sub_38_add_2_17_lut (.I0(n60274), .I1(n294[15]), .I2(VCC_net), 
            .I3(n49301), .O(n60276)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i5578_2_lut_4_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n42_adj_4462));   // verilog/uart_rx.v(119[33:55])
    defparam i5578_2_lut_4_lut_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[24] ), .I2(n27), 
            .I3(GND_net), .O(n14));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3488[12] ), .I2(n23), .I3(n4937), 
            .O(n15));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(\o_Rx_DV_N_3488[8] ), .I2(n14), .I3(n56959), 
            .O(n69533));
    defparam i8_4_lut.LUT_INIT = 16'h2000;
    SB_CARRY sub_38_add_2_17 (.CI(n49301), .I0(n294[15]), .I1(VCC_net), 
            .CO(n49302));
    SB_LUT4 i1_4_lut_adj_976 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4937), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n60728), .O(n60734));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_976.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_977 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n60734), .O(n60740));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_977.LUT_INIT = 16'hfffe;
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk16MHz), .D(n29884));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i1_4_lut_adj_978 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4937), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n60776), .O(n60782));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_978.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_979 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n60782), .O(n60788));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_979.LUT_INIT = 16'hfffe;
    SB_LUT4 i5592_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n58597), .I3(n44_adj_4463), 
            .O(n46_adj_4464));   // verilog/uart_rx.v(119[33:55])
    defparam i5592_4_lut.LUT_INIT = 16'hb3a0;
    SB_LUT4 div_37_i639_4_lut (.I0(n57840), .I1(n294[19]), .I2(n46_adj_4464), 
            .I3(baudrate[4]), .O(n57842));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i639_4_lut.LUT_INIT = 16'h6aa6;
    SB_LUT4 i1_2_lut (.I0(baudrate[25]), .I1(baudrate[29]), .I2(GND_net), 
            .I3(GND_net), .O(n61900));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i641_4_lut (.I0(n804), .I1(n42_adj_4462), .I2(n294[19]), 
            .I3(baudrate[2]), .O(n960));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i641_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i1_4_lut_adj_980 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4937), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n60744), .O(n60750));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_980.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_981 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n60750), .O(n60756));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_981.LUT_INIT = 16'hfffe;
    SB_LUT4 i7237_4_lut (.I0(n804), .I1(n42863), .I2(n20919), .I3(baudrate[2]), 
            .O(n20921));   // verilog/uart_rx.v(119[33:55])
    defparam i7237_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 div_37_i640_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n294[19]), 
            .I3(n44_adj_4463), .O(n959));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i640_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i642_4_lut (.I0(n805), .I1(baudrate[1]), .I2(n294[19]), 
            .I3(baudrate[0]), .O(n961));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i642_4_lut.LUT_INIT = 16'h9a6a;
    SB_LUT4 i1_2_lut_adj_982 (.I0(baudrate[24]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n61902));
    defparam i1_2_lut_adj_982.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_983 (.I0(n61798), .I1(n61794), .I2(n61796), .I3(n61792), 
            .O(n61778));
    defparam i1_4_lut_adj_983.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_984 (.I0(n61900), .I1(n61676), .I2(n61790), .I3(n61666), 
            .O(n25629));
    defparam i1_4_lut_adj_984.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_985 (.I0(n61658), .I1(n25629), .I2(n61778), .I3(n61656), 
            .O(n25545));
    defparam i1_4_lut_adj_985.LUT_INIT = 16'hfffe;
    SB_LUT4 i28970_rep_6_2_lut (.I0(baudrate[0]), .I1(n294[19]), .I2(GND_net), 
            .I3(GND_net), .O(n58123));   // verilog/uart_rx.v(119[33:55])
    defparam i28970_rep_6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_38_add_2_16_lut (.I0(n60366), .I1(n294[14]), .I2(VCC_net), 
            .I3(n49300), .O(n60368)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 div_37_LessThan_662_i42_4_lut (.I0(n58123), .I1(baudrate[2]), 
            .I2(n961), .I3(baudrate[1]), .O(n42_adj_4465));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i42_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i51940_3_lut (.I0(n42_adj_4465), .I1(baudrate[3]), .I2(n960), 
            .I3(GND_net), .O(n67626));   // verilog/uart_rx.v(119[33:55])
    defparam i51940_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51941_3_lut (.I0(n67626), .I1(baudrate[4]), .I2(n959), .I3(GND_net), 
            .O(n67627));   // verilog/uart_rx.v(119[33:55])
    defparam i51941_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_662_i48_3_lut (.I0(n67627), .I1(baudrate[5]), 
            .I2(n57842), .I3(GND_net), .O(n48));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i52835_2_lut (.I0(n48), .I1(n25545), .I2(GND_net), .I3(GND_net), 
            .O(n294[18]));   // verilog/uart_rx.v(119[33:55])
    defparam i52835_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_37_i534_3_lut (.I0(n57838), .I1(n294[20]), .I2(baudrate[3]), 
            .I3(GND_net), .O(n57840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i534_3_lut.LUT_INIT = 16'h6a6a;
    SB_CARRY sub_38_add_2_16 (.CI(n49300), .I0(n294[14]), .I1(VCC_net), 
            .CO(n49301));
    SB_LUT4 sub_38_add_2_15_lut (.I0(o_Rx_DV_N_3488[10]), .I1(n294[13]), 
            .I2(VCC_net), .I3(n49299), .O(n60366)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_15 (.CI(n49299), .I0(n294[13]), .I1(VCC_net), 
            .CO(n49300));
    SB_LUT4 sub_38_add_2_14_lut (.I0(GND_net), .I1(n294[12]), .I2(VCC_net), 
            .I3(n49298), .O(\o_Rx_DV_N_3488[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_14 (.CI(n49298), .I0(n294[12]), .I1(VCC_net), 
            .CO(n49299));
    SB_LUT4 sub_38_add_2_13_lut (.I0(o_Rx_DV_N_3488[9]), .I1(n294[11]), 
            .I2(VCC_net), .I3(n49297), .O(n60274)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_13_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_13 (.CI(n49297), .I0(n294[11]), .I1(VCC_net), 
            .CO(n49298));
    SB_LUT4 sub_38_add_2_12_lut (.I0(GND_net), .I1(n294[10]), .I2(VCC_net), 
            .I3(n49296), .O(o_Rx_DV_N_3488[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_12 (.CI(n49296), .I0(n294[10]), .I1(VCC_net), 
            .CO(n49297));
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk16MHz), .D(n29866));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i46893_2_lut (.I0(baudrate[8]), .I1(n62568), .I2(GND_net), 
            .I3(GND_net), .O(n62570));
    defparam i46893_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i50609_4_lut (.I0(n25589), .I1(n65720), .I2(n48_adj_4466), 
            .I3(baudrate[0]), .O(n804));
    defparam i50609_4_lut.LUT_INIT = 16'h3633;
    SB_LUT4 div_37_i535_4_lut (.I0(n68343), .I1(n44_adj_4467), .I2(n294[20]), 
            .I3(baudrate[2]), .O(n803));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i535_4_lut.LUT_INIT = 16'h9565;
    SB_LUT4 i1_3_lut_adj_986 (.I0(n25632), .I1(n48_adj_4468), .I2(baudrate[0]), 
            .I3(GND_net), .O(n805));
    defparam i1_3_lut_adj_986.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_LessThan_557_i42_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n805), .I3(GND_net), .O(n42_adj_4469));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i42_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51942_3_lut (.I0(n42_adj_4469), .I1(baudrate[2]), .I2(n804), 
            .I3(GND_net), .O(n67628));   // verilog/uart_rx.v(119[33:55])
    defparam i51942_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51943_3_lut (.I0(n67628), .I1(baudrate[3]), .I2(n803), .I3(GND_net), 
            .O(n67629));   // verilog/uart_rx.v(119[33:55])
    defparam i51943_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_557_i48_3_lut (.I0(n67629), .I1(baudrate[4]), 
            .I2(n57840), .I3(GND_net), .O(n48_adj_4470));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 sub_38_add_2_11_lut (.I0(GND_net), .I1(n294[9]), .I2(VCC_net), 
            .I3(n49295), .O(o_Rx_DV_N_3488[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_11 (.CI(n49295), .I0(n294[9]), .I1(VCC_net), 
            .CO(n49296));
    SB_LUT4 sub_38_add_2_10_lut (.I0(GND_net), .I1(n294[8]), .I2(VCC_net), 
            .I3(n49294), .O(\o_Rx_DV_N_3488[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_10 (.CI(n49294), .I0(n294[8]), .I1(VCC_net), 
            .CO(n49295));
    SB_LUT4 sub_38_add_2_9_lut (.I0(GND_net), .I1(n294[7]), .I2(VCC_net), 
            .I3(n49293), .O(\o_Rx_DV_N_3488[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_9 (.CI(n49293), .I0(n294[7]), .I1(VCC_net), 
            .CO(n49294));
    SB_LUT4 sub_38_add_2_8_lut (.I0(GND_net), .I1(n294[6]), .I2(VCC_net), 
            .I3(n49292), .O(\o_Rx_DV_N_3488[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_8 (.CI(n49292), .I0(n294[6]), .I1(VCC_net), 
            .CO(n49293));
    SB_LUT4 sub_38_add_2_7_lut (.I0(GND_net), .I1(n294[5]), .I2(VCC_net), 
            .I3(n49291), .O(\o_Rx_DV_N_3488[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_7 (.CI(n49291), .I0(n294[5]), .I1(VCC_net), 
            .CO(n49292));
    SB_LUT4 sub_38_add_2_6_lut (.I0(GND_net), .I1(n294[4]), .I2(VCC_net), 
            .I3(n49290), .O(\o_Rx_DV_N_3488[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_6 (.CI(n49290), .I0(n294[4]), .I1(VCC_net), 
            .CO(n49291));
    SB_LUT4 sub_38_add_2_5_lut (.I0(GND_net), .I1(n294[3]), .I2(VCC_net), 
            .I3(n49289), .O(\o_Rx_DV_N_3488[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_5 (.CI(n49289), .I0(n294[3]), .I1(VCC_net), 
            .CO(n49290));
    SB_LUT4 sub_38_add_2_4_lut (.I0(GND_net), .I1(n294[2]), .I2(VCC_net), 
            .I3(n49288), .O(\o_Rx_DV_N_3488[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_4 (.CI(n49288), .I0(n294[2]), .I1(VCC_net), 
            .CO(n49289));
    SB_LUT4 sub_38_add_2_3_lut (.I0(GND_net), .I1(n294[1]), .I2(VCC_net), 
            .I3(n49287), .O(\o_Rx_DV_N_3488[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_3 (.CI(n49287), .I0(n294[1]), .I1(VCC_net), 
            .CO(n49288));
    SB_LUT4 sub_38_add_2_2_lut (.I0(GND_net), .I1(n59155), .I2(GND_net), 
            .I3(VCC_net), .O(\o_Rx_DV_N_3488[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_2 (.CI(VCC_net), .I0(n59155), .I1(GND_net), 
            .CO(n49287));
    SB_LUT4 i46648_2_lut (.I0(baudrate[17]), .I1(n25619), .I2(GND_net), 
            .I3(GND_net), .O(n62318));
    defparam i46648_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_987 (.I0(n61656), .I1(n61798), .I2(baudrate[16]), 
            .I3(n42863), .O(n60908));
    defparam i1_4_lut_adj_987.LUT_INIT = 16'h0100;
    SB_LUT4 i50740_3_lut (.I0(n58609), .I1(n59474), .I2(baudrate[2]), 
            .I3(GND_net), .O(n65325));   // verilog/uart_rx.v(119[33:55])
    defparam i50740_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i50590_4_lut (.I0(n57899), .I1(n60908), .I2(n61658), .I3(n60962), 
            .O(n65326));   // verilog/uart_rx.v(119[33:55])
    defparam i50590_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 div_37_i427_4_lut (.I0(n65326), .I1(n65325), .I2(n294[21]), 
            .I3(n62318), .O(n57838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i427_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i1_2_lut_adj_988 (.I0(baudrate[26]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n61898));
    defparam i1_2_lut_adj_988.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_989 (.I0(baudrate[23]), .I1(baudrate[28]), .I2(baudrate[27]), 
            .I3(baudrate[0]), .O(n60642));
    defparam i1_4_lut_adj_989.LUT_INIT = 16'h0100;
    SB_LUT4 i46857_4_lut (.I0(baudrate[25]), .I1(baudrate[31]), .I2(baudrate[24]), 
            .I3(baudrate[29]), .O(n62534));
    defparam i46857_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_990 (.I0(n57899), .I1(n60642), .I2(n61898), .I3(baudrate[16]), 
            .O(n60670));
    defparam i1_4_lut_adj_990.LUT_INIT = 16'h0004;
    SB_LUT4 i46925_4_lut (.I0(n62534), .I1(n62532), .I2(n62472), .I3(n62450), 
            .O(n62602));
    defparam i46925_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52657_4_lut (.I0(n62592), .I1(n65714), .I2(n62602), .I3(n60670), 
            .O(n68343));
    defparam i52657_4_lut.LUT_INIT = 16'hc9cc;
    SB_LUT4 i1_2_lut_adj_991 (.I0(baudrate[16]), .I1(baudrate[17]), .I2(GND_net), 
            .I3(GND_net), .O(n61796));
    defparam i1_2_lut_adj_991.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_992 (.I0(baudrate[28]), .I1(baudrate[27]), .I2(baudrate[31]), 
            .I3(baudrate[26]), .O(n60990));
    defparam i1_4_lut_adj_992.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_993 (.I0(n60990), .I1(n61804), .I2(n61748), .I3(n61744), 
            .O(n25644));
    defparam i1_4_lut_adj_993.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_994 (.I0(baudrate[6]), .I1(baudrate[7]), .I2(GND_net), 
            .I3(GND_net), .O(n61650));
    defparam i1_2_lut_adj_994.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_995 (.I0(baudrate[8]), .I1(baudrate[9]), .I2(GND_net), 
            .I3(GND_net), .O(n61648));
    defparam i1_2_lut_adj_995.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_996 (.I0(baudrate[4]), .I1(baudrate[5]), .I2(GND_net), 
            .I3(GND_net), .O(n60962));
    defparam i1_2_lut_adj_996.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_997 (.I0(n60962), .I1(n61648), .I2(n61650), .I3(n61646), 
            .O(n60974));
    defparam i1_4_lut_adj_997.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_998 (.I0(n60974), .I1(n25644), .I2(n60966), .I3(n61806), 
            .O(n25632));
    defparam i1_4_lut_adj_998.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_450_i46_4_lut (.I0(n65404), .I1(baudrate[2]), 
            .I2(n68343), .I3(n48_adj_4466), .O(n46_adj_4471));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i46_4_lut.LUT_INIT = 16'hc0e8;
    SB_LUT4 div_37_LessThan_450_i48_3_lut (.I0(n46_adj_4471), .I1(baudrate[3]), 
            .I2(n57838), .I3(GND_net), .O(n48_adj_4468));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i52832_2_lut (.I0(n48_adj_4468), .I1(n25632), .I2(GND_net), 
            .I3(GND_net), .O(n294[20]));   // verilog/uart_rx.v(119[33:55])
    defparam i52832_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_3_lut_4_lut (.I0(baudrate[30]), .I1(baudrate[31]), .I2(baudrate[27]), 
            .I3(baudrate[24]), .O(n60292));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_999 (.I0(baudrate[14]), .I1(baudrate[15]), .I2(GND_net), 
            .I3(GND_net), .O(n61798));
    defparam i1_2_lut_adj_999.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1000 (.I0(baudrate[12]), .I1(baudrate[13]), .I2(GND_net), 
            .I3(GND_net), .O(n61644));
    defparam i1_2_lut_adj_1000.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1001 (.I0(baudrate[10]), .I1(baudrate[11]), .I2(GND_net), 
            .I3(GND_net), .O(n61646));
    defparam i1_2_lut_adj_1001.LUT_INIT = 16'heeee;
    SB_LUT4 i46809_2_lut (.I0(baudrate[21]), .I1(baudrate[22]), .I2(GND_net), 
            .I3(GND_net), .O(n62486));
    defparam i46809_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i46915_4_lut (.I0(n62486), .I1(n60966), .I2(n61646), .I3(baudrate[9]), 
            .O(n62592));
    defparam i46915_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i28963_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n42865));
    defparam i28963_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1002 (.I0(baudrate[18]), .I1(baudrate[19]), .I2(GND_net), 
            .I3(GND_net), .O(n61794));
    defparam i1_2_lut_adj_1002.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1003 (.I0(n61804), .I1(n60294), .I2(n60292), 
            .I3(n61794), .O(n25619));
    defparam i1_4_lut_adj_1003.LUT_INIT = 16'hfffe;
    SB_LUT4 i28961_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n42863));
    defparam i28961_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1004 (.I0(baudrate[17]), .I1(n62504), .I2(baudrate[2]), 
            .I3(n42863), .O(n60252));
    defparam i1_4_lut_adj_1004.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1005 (.I0(n62556), .I1(n60252), .I2(n25619), 
            .I3(n62532), .O(n59474));
    defparam i1_4_lut_adj_1005.LUT_INIT = 16'h0004;
    SB_LUT4 i46863_3_lut_4_lut (.I0(baudrate[30]), .I1(baudrate[31]), .I2(baudrate[26]), 
            .I3(baudrate[24]), .O(n62540));
    defparam i46863_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1006 (.I0(baudrate[23]), .I1(baudrate[27]), .I2(baudrate[25]), 
            .I3(n42865), .O(n60586));
    defparam i1_4_lut_adj_1006.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1007 (.I0(n60586), .I1(baudrate[29]), .I2(baudrate[16]), 
            .I3(baudrate[28]), .O(n60604));
    defparam i1_4_lut_adj_1007.LUT_INIT = 16'h0002;
    SB_LUT4 i46927_4_lut (.I0(n62540), .I1(n62532), .I2(n62472), .I3(n62450), 
            .O(n62604));
    defparam i46927_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1008 (.I0(n62592), .I1(n62604), .I2(n57899), 
            .I3(n60604), .O(n58609));
    defparam i1_4_lut_adj_1008.LUT_INIT = 16'h0100;
    SB_LUT4 div_37_LessThan_341_i48_3_lut (.I0(n58609), .I1(baudrate[2]), 
            .I2(n59474), .I3(GND_net), .O(n48_adj_4466));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_341_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i53463_2_lut (.I0(n48_adj_4466), .I1(n25589), .I2(GND_net), 
            .I3(GND_net), .O(n294[21]));
    defparam i53463_2_lut.LUT_INIT = 16'h1111;
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk16MHz), .D(n29774));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk16MHz), .D(n29773));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk16MHz), .D(n29772));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(clk16MHz), .D(n69533));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_2210_i39_4_lut (.I0(n3155), .I1(baudrate[19]), 
            .I2(n8425[19]), .I3(n294[1]), .O(n39_adj_4472));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i39_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i41_4_lut (.I0(n3154), .I1(baudrate[20]), 
            .I2(n8425[20]), .I3(n294[1]), .O(n41_adj_4473));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i41_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i33_4_lut (.I0(n3158), .I1(baudrate[16]), 
            .I2(n8425[16]), .I3(n294[1]), .O(n33));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i33_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i35_4_lut (.I0(n3157), .I1(baudrate[17]), 
            .I2(n8425[17]), .I3(n294[1]), .O(n35));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i35_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i37_4_lut (.I0(n3156), .I1(baudrate[18]), 
            .I2(n8425[18]), .I3(n294[1]), .O(n37));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i37_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i23_4_lut (.I0(n3163), .I1(baudrate[11]), 
            .I2(n8425[11]), .I3(n294[1]), .O(n23_adj_4474));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i23_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i25_4_lut (.I0(n3162), .I1(baudrate[12]), 
            .I2(n8425[12]), .I3(n294[1]), .O(n25));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i25_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i29_4_lut (.I0(n3160), .I1(baudrate[14]), 
            .I2(n8425[14]), .I3(n294[1]), .O(n29_adj_4475));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i29_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i31_4_lut (.I0(n3159), .I1(baudrate[15]), 
            .I2(n8425[15]), .I3(n294[1]), .O(n31));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i31_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i7_4_lut (.I0(n3171), .I1(baudrate[3]), 
            .I2(n8425[3]), .I3(n294[1]), .O(n7));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i7_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i45_4_lut (.I0(n3152), .I1(baudrate[22]), 
            .I2(n8425[22]), .I3(n294[1]), .O(n45_adj_4476));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i45_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i43_4_lut (.I0(n3153), .I1(baudrate[21]), 
            .I2(n8425[21]), .I3(n294[1]), .O(n43_adj_4477));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i43_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i9_4_lut (.I0(n3170), .I1(baudrate[4]), 
            .I2(n8425[4]), .I3(n294[1]), .O(n9));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i9_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i17_4_lut (.I0(n3166), .I1(baudrate[8]), 
            .I2(n8425[8]), .I3(n294[1]), .O(n17));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i17_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i19_4_lut (.I0(n3165), .I1(baudrate[9]), 
            .I2(n8425[9]), .I3(n294[1]), .O(n19));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i19_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i21_4_lut (.I0(n3164), .I1(baudrate[10]), 
            .I2(n8425[10]), .I3(n294[1]), .O(n21));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i21_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i11_4_lut (.I0(n3169), .I1(baudrate[5]), 
            .I2(n8425[5]), .I3(n294[1]), .O(n11));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i11_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i13_4_lut (.I0(n3168), .I1(baudrate[6]), 
            .I2(n8425[6]), .I3(n294[1]), .O(n13));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i13_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i1_2_lut_3_lut (.I0(\r_SM_Main[1] ), .I1(r_SM_Main[0]), .I2(\r_SM_Main[2] ), 
            .I3(GND_net), .O(n4));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 div_37_LessThan_2210_i15_4_lut (.I0(n3167), .I1(baudrate[7]), 
            .I2(n8425[7]), .I3(n294[1]), .O(n15_adj_4478));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i15_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i27_4_lut (.I0(n3161), .I1(baudrate[13]), 
            .I2(n8425[13]), .I3(n294[1]), .O(n27_adj_4479));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i27_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i49932_4_lut (.I0(n27_adj_4479), .I1(n15_adj_4478), .I2(n13), 
            .I3(n11), .O(n65618));
    defparam i49932_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i49939_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n65625));
    defparam i49939_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2210_i16_3_lut (.I0(baudrate[9]), .I1(baudrate[21]), 
            .I2(n43_adj_4477), .I3(GND_net), .O(n16));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49910_2_lut (.I0(n43_adj_4477), .I1(n19), .I2(GND_net), .I3(GND_net), 
            .O(n65596));
    defparam i49910_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2210_i8_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n17), .I3(GND_net), .O(n8));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i24_3_lut (.I0(n16), .I1(baudrate[22]), 
            .I2(n45_adj_4476), .I3(GND_net), .O(n24));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2208_3_lut (.I0(n3172), .I1(n8425[2]), .I2(n294[1]), 
            .I3(GND_net), .O(n3274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49950_3_lut (.I0(n7), .I1(n3274), .I2(baudrate[2]), .I3(GND_net), 
            .O(n65636));
    defparam i49950_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 i50840_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n65636), 
            .O(n66526));
    defparam i50840_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i50836_4_lut (.I0(n19), .I1(n17), .I2(n15_adj_4478), .I3(n66526), 
            .O(n66522));
    defparam i50836_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52196_4_lut (.I0(n25), .I1(n23_adj_4474), .I2(n21), .I3(n66522), 
            .O(n67882));
    defparam i52196_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51569_4_lut (.I0(n31), .I1(n29_adj_4475), .I2(n27_adj_4479), 
            .I3(n67882), .O(n67255));
    defparam i51569_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52427_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n67255), 
            .O(n68113));
    defparam i52427_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2210_i12_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n33), .I3(GND_net), .O(n12));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i4_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n60336), .I3(n48_adj_4480), .O(n4_adj_4481));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i4_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i52127_3_lut (.I0(n4_adj_4481), .I1(baudrate[13]), .I2(n27_adj_4479), 
            .I3(GND_net), .O(n67813));   // verilog/uart_rx.v(119[33:55])
    defparam i52127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52128_3_lut (.I0(n67813), .I1(baudrate[14]), .I2(n29_adj_4475), 
            .I3(GND_net), .O(n67814));   // verilog/uart_rx.v(119[33:55])
    defparam i52128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49924_2_lut (.I0(n33), .I1(n15_adj_4478), .I2(GND_net), .I3(GND_net), 
            .O(n65610));
    defparam i49924_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2210_i10_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n13), .I3(GND_net), .O(n10));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i30_3_lut (.I0(n12), .I1(baudrate[17]), 
            .I2(n35), .I3(GND_net), .O(n30));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49926_4_lut (.I0(n33), .I1(n31), .I2(n29_adj_4475), .I3(n65618), 
            .O(n65612));
    defparam i49926_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52483_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n65610), 
            .O(n68169));   // verilog/uart_rx.v(119[33:55])
    defparam i52483_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52068_3_lut (.I0(n67814), .I1(baudrate[15]), .I2(n31), .I3(GND_net), 
            .O(n67754));   // verilog/uart_rx.v(119[33:55])
    defparam i52068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52609_4_lut (.I0(n67754), .I1(n68169), .I2(n35), .I3(n65612), 
            .O(n68295));   // verilog/uart_rx.v(119[33:55])
    defparam i52609_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52610_3_lut (.I0(n68295), .I1(baudrate[18]), .I2(n37), .I3(GND_net), 
            .O(n68296));   // verilog/uart_rx.v(119[33:55])
    defparam i52610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i6_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n7), .I3(GND_net), .O(n6));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52129_3_lut (.I0(n6), .I1(baudrate[10]), .I2(n21), .I3(GND_net), 
            .O(n67815));   // verilog/uart_rx.v(119[33:55])
    defparam i52129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52130_3_lut (.I0(n67815), .I1(baudrate[11]), .I2(n23_adj_4474), 
            .I3(GND_net), .O(n67816));   // verilog/uart_rx.v(119[33:55])
    defparam i52130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49915_4_lut (.I0(n43_adj_4477), .I1(n25), .I2(n23_adj_4474), 
            .I3(n65625), .O(n65601));
    defparam i49915_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51711_4_lut (.I0(n24), .I1(n8), .I2(n45_adj_4476), .I3(n65596), 
            .O(n67397));   // verilog/uart_rx.v(119[33:55])
    defparam i51711_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52066_3_lut (.I0(n67816), .I1(baudrate[12]), .I2(n25), .I3(GND_net), 
            .O(n67752));   // verilog/uart_rx.v(119[33:55])
    defparam i52066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52548_3_lut (.I0(n68296), .I1(baudrate[19]), .I2(n39_adj_4472), 
            .I3(GND_net), .O(n68234));   // verilog/uart_rx.v(119[33:55])
    defparam i52548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49917_4_lut (.I0(n43_adj_4477), .I1(n41_adj_4473), .I2(n39_adj_4472), 
            .I3(n68113), .O(n65603));
    defparam i49917_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52315_4_lut (.I0(n67752), .I1(n67397), .I2(n45_adj_4476), 
            .I3(n65601), .O(n68001));   // verilog/uart_rx.v(119[33:55])
    defparam i52315_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52541_3_lut (.I0(n68234), .I1(baudrate[20]), .I2(n41_adj_4473), 
            .I3(GND_net), .O(n40_adj_4482));   // verilog/uart_rx.v(119[33:55])
    defparam i52541_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1009 (.I0(baudrate[25]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n60264));
    defparam i1_2_lut_adj_1009.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i2187_3_lut (.I0(n3151), .I1(n8425[23]), .I2(n294[1]), 
            .I3(GND_net), .O(n3253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52317_4_lut (.I0(n40_adj_4482), .I1(n68001), .I2(n45_adj_4476), 
            .I3(n65603), .O(n68003));   // verilog/uart_rx.v(119[33:55])
    defparam i52317_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_adj_1010 (.I0(baudrate[30]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n61744));
    defparam i1_2_lut_adj_1010.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1011 (.I0(n61898), .I1(n61748), .I2(n60264), 
            .I3(n61746), .O(n60272));
    defparam i1_4_lut_adj_1011.LUT_INIT = 16'hfffe;
    SB_LUT4 i53023_4_lut (.I0(n60272), .I1(n68003), .I2(baudrate[23]), 
            .I3(n3253), .O(n59155));   // verilog/uart_rx.v(119[33:55])
    defparam i53023_4_lut.LUT_INIT = 16'h1501;
    SB_LUT4 i46771_2_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62448));
    defparam i46771_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i46879_4_lut (.I0(n60826), .I1(n60822), .I2(n60824), .I3(n60820), 
            .O(n62556));
    defparam i46879_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i42262_2_lut (.I0(baudrate[2]), .I1(baudrate[3]), .I2(GND_net), 
            .I3(GND_net), .O(n57899));
    defparam i42262_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i46837_3_lut (.I0(baudrate[31]), .I1(baudrate[21]), .I2(baudrate[27]), 
            .I3(GND_net), .O(n62514));
    defparam i46837_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i46897_4_lut (.I0(n62514), .I1(n61790), .I2(n62512), .I3(n61744), 
            .O(n62574));
    defparam i46897_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i46923_4_lut (.I0(n62574), .I1(n62532), .I2(n57899), .I3(baudrate[4]), 
            .O(n62600));
    defparam i46923_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53445_4_lut (.I0(n62556), .I1(n62450), .I2(n62600), .I3(n62448), 
            .O(n62610));
    defparam i53445_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_i2118_3_lut (.I0(n3046), .I1(n8399[23]), .I2(n294[2]), 
            .I3(GND_net), .O(n3151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2119_3_lut (.I0(n3047), .I1(n8399[22]), .I2(n294[2]), 
            .I3(GND_net), .O(n3152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2120_3_lut (.I0(n3048), .I1(n8399[21]), .I2(n294[2]), 
            .I3(GND_net), .O(n3153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2121_3_lut (.I0(n3049), .I1(n8399[20]), .I2(n294[2]), 
            .I3(GND_net), .O(n3154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2135_3_lut (.I0(n3063), .I1(n8399[6]), .I2(n294[2]), 
            .I3(GND_net), .O(n3168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1012 (.I0(n60830), .I1(n62572), .I2(baudrate[0]), 
            .I3(n48_adj_4470), .O(n962));
    defparam i1_3_lut_4_lut_adj_1012.LUT_INIT = 16'h0010;
    SB_LUT4 div_37_i2122_3_lut (.I0(n3050), .I1(n8399[19]), .I2(n294[2]), 
            .I3(GND_net), .O(n3155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2125_3_lut (.I0(n3053), .I1(n8399[16]), .I2(n294[2]), 
            .I3(GND_net), .O(n3158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i33_2_lut (.I0(n3158), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4483));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2126_3_lut (.I0(n3054), .I1(n8399[15]), .I2(n294[2]), 
            .I3(GND_net), .O(n3159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i31_2_lut (.I0(n3159), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4484));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2123_3_lut (.I0(n3051), .I1(n8399[18]), .I2(n294[2]), 
            .I3(GND_net), .O(n3156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i37_2_lut (.I0(n3156), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4485));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2124_3_lut (.I0(n3052), .I1(n8399[17]), .I2(n294[2]), 
            .I3(GND_net), .O(n3157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i35_2_lut (.I0(n3157), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4486));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2130_3_lut (.I0(n3058), .I1(n8399[11]), .I2(n294[2]), 
            .I3(GND_net), .O(n3163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2131_3_lut (.I0(n3059), .I1(n8399[10]), .I2(n294[2]), 
            .I3(GND_net), .O(n3164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i21_2_lut (.I0(n3164), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4487));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i23_2_lut (.I0(n3163), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4488));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2129_3_lut (.I0(n3057), .I1(n8399[12]), .I2(n294[2]), 
            .I3(GND_net), .O(n3162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2128_3_lut (.I0(n3056), .I1(n8399[13]), .I2(n294[2]), 
            .I3(GND_net), .O(n3161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i25_2_lut (.I0(n3162), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4489));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i27_2_lut (.I0(n3161), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4490));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2137_3_lut (.I0(n3065), .I1(n8399[4]), .I2(n294[2]), 
            .I3(GND_net), .O(n3170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2138_3_lut (.I0(n3066), .I1(n8399[3]), .I2(n294[2]), 
            .I3(GND_net), .O(n3171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i9_2_lut (.I0(n3170), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4491));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2127_3_lut (.I0(n3055), .I1(n8399[14]), .I2(n294[2]), 
            .I3(GND_net), .O(n3160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2134_3_lut (.I0(n3062), .I1(n8399[7]), .I2(n294[2]), 
            .I3(GND_net), .O(n3167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2133_3_lut (.I0(n3061), .I1(n8399[8]), .I2(n294[2]), 
            .I3(GND_net), .O(n3166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i13_2_lut (.I0(n3168), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4492));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i15_2_lut (.I0(n3167), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4493));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i17_2_lut (.I0(n3166), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4494));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i29_2_lut (.I0(n3160), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4495));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2132_3_lut (.I0(n3060), .I1(n8399[9]), .I2(n294[2]), 
            .I3(GND_net), .O(n3165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2136_3_lut (.I0(n3064), .I1(n8399[5]), .I2(n294[2]), 
            .I3(GND_net), .O(n3169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i11_2_lut (.I0(n3169), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4496));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i19_2_lut (.I0(n3165), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4497));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1013 (.I0(n61646), .I1(n62546), .I2(n8087[14]), 
            .I3(n48_adj_4498), .O(n1702));
    defparam i1_3_lut_4_lut_adj_1013.LUT_INIT = 16'h0010;
    SB_LUT4 i1_4_lut_adj_1014 (.I0(n61902), .I1(n61904), .I2(n61746), 
            .I3(n61900), .O(n25552));
    defparam i1_4_lut_adj_1014.LUT_INIT = 16'hfffe;
    SB_LUT4 i49983_4_lut (.I0(n29_adj_4495), .I1(n17_adj_4494), .I2(n15_adj_4493), 
            .I3(n13_adj_4492), .O(n65669));
    defparam i49983_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50943_4_lut (.I0(n11_adj_4496), .I1(n9_adj_4491), .I2(n3171), 
            .I3(baudrate[2]), .O(n66629));
    defparam i50943_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i51617_4_lut (.I0(n17_adj_4494), .I1(n15_adj_4493), .I2(n13_adj_4492), 
            .I3(n66629), .O(n67303));
    defparam i51617_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51615_4_lut (.I0(n23_adj_4488), .I1(n21_adj_4487), .I2(n19_adj_4497), 
            .I3(n67303), .O(n67301));
    defparam i51615_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i49996_4_lut (.I0(n29_adj_4495), .I1(n27_adj_4490), .I2(n25_adj_4489), 
            .I3(n67301), .O(n65682));
    defparam i49996_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2141_i6_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3172), .I3(GND_net), .O(n6_adj_4499));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52135_3_lut (.I0(n6_adj_4499), .I1(baudrate[13]), .I2(n29_adj_4495), 
            .I3(GND_net), .O(n67821));   // verilog/uart_rx.v(119[33:55])
    defparam i52135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i32_3_lut (.I0(n14_adj_4500), .I1(baudrate[17]), 
            .I2(n37_adj_4485), .I3(GND_net), .O(n32));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52136_3_lut (.I0(n67821), .I1(baudrate[14]), .I2(n31_adj_4484), 
            .I3(GND_net), .O(n67822));   // verilog/uart_rx.v(119[33:55])
    defparam i52136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49976_4_lut (.I0(n35_adj_4486), .I1(n33_adj_4483), .I2(n31_adj_4484), 
            .I3(n65669), .O(n65662));
    defparam i49976_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52481_4_lut (.I0(n32), .I1(n12_adj_4501), .I2(n37_adj_4485), 
            .I3(n65660), .O(n68167));   // verilog/uart_rx.v(119[33:55])
    defparam i52481_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52058_3_lut (.I0(n67822), .I1(baudrate[15]), .I2(n33_adj_4483), 
            .I3(GND_net), .O(n67744));   // verilog/uart_rx.v(119[33:55])
    defparam i52058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1015 (.I0(n60822), .I1(n62350), .I2(n8165[11]), 
            .I3(n48_adj_4502), .O(n2110));
    defparam i1_3_lut_4_lut_adj_1015.LUT_INIT = 16'h0010;
    SB_LUT4 i52309_3_lut (.I0(n8_adj_4503), .I1(baudrate[10]), .I2(n23_adj_4488), 
            .I3(GND_net), .O(n67995));   // verilog/uart_rx.v(119[33:55])
    defparam i52309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52310_3_lut (.I0(n67995), .I1(baudrate[11]), .I2(n25_adj_4489), 
            .I3(GND_net), .O(n67996));   // verilog/uart_rx.v(119[33:55])
    defparam i52310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Clock_Count_1951_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n50546), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1951_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n50545), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_8 (.CI(n50545), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n50546));
    SB_LUT4 r_Clock_Count_1951_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n50544), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50929_4_lut (.I0(n25_adj_4489), .I1(n23_adj_4488), .I2(n21_adj_4487), 
            .I3(n65696), .O(n66615));
    defparam i50929_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51707_3_lut (.I0(n10_adj_4507), .I1(baudrate[9]), .I2(n21_adj_4487), 
            .I3(GND_net), .O(n67393));   // verilog/uart_rx.v(119[33:55])
    defparam i51707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52056_3_lut (.I0(n67996), .I1(baudrate[12]), .I2(n27_adj_4490), 
            .I3(GND_net), .O(n67742));   // verilog/uart_rx.v(119[33:55])
    defparam i52056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51914_4_lut (.I0(n35_adj_4486), .I1(n33_adj_4483), .I2(n31_adj_4484), 
            .I3(n65682), .O(n67600));
    defparam i51914_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY r_Clock_Count_1951_add_4_7 (.CI(n50544), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n50545));
    SB_LUT4 i52607_4_lut (.I0(n67744), .I1(n68167), .I2(n37_adj_4485), 
            .I3(n65662), .O(n68293));   // verilog/uart_rx.v(119[33:55])
    defparam i52607_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52131_4_lut (.I0(n67742), .I1(n67393), .I2(n27_adj_4490), 
            .I3(n66615), .O(n67817));   // verilog/uart_rx.v(119[33:55])
    defparam i52131_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52629_4_lut (.I0(n67817), .I1(n68293), .I2(n37_adj_4485), 
            .I3(n67600), .O(n68315));   // verilog/uart_rx.v(119[33:55])
    defparam i52629_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52630_3_lut (.I0(n68315), .I1(baudrate[18]), .I2(n3155), 
            .I3(GND_net), .O(n68316));   // verilog/uart_rx.v(119[33:55])
    defparam i52630_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 r_Clock_Count_1951_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n50543), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_6 (.CI(n50543), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n50544));
    SB_LUT4 i52620_3_lut (.I0(n68316), .I1(baudrate[19]), .I2(n3154), 
            .I3(GND_net), .O(n68306));   // verilog/uart_rx.v(119[33:55])
    defparam i52620_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52421_3_lut (.I0(n68306), .I1(baudrate[20]), .I2(n3153), 
            .I3(GND_net), .O(n68107));   // verilog/uart_rx.v(119[33:55])
    defparam i52421_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 r_Clock_Count_1951_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n50542), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_5 (.CI(n50542), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n50543));
    SB_LUT4 i52422_3_lut (.I0(n68107), .I1(baudrate[21]), .I2(n3152), 
            .I3(GND_net), .O(n68108));   // verilog/uart_rx.v(119[33:55])
    defparam i52422_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 r_Clock_Count_1951_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n50541), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52064_3_lut (.I0(n68108), .I1(baudrate[22]), .I2(n3151), 
            .I3(GND_net), .O(n48_adj_4480));   // verilog/uart_rx.v(119[33:55])
    defparam i52064_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY r_Clock_Count_1951_add_4_4 (.CI(n50541), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n50542));
    SB_LUT4 r_Clock_Count_1951_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n50540), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_3 (.CI(n50540), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n50541));
    SB_LUT4 r_Clock_Count_1951_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1951_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1951_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n50540));
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n27966), 
            .D(n479[1]), .R(n58000));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n27966), 
            .D(n479[2]), .R(n58000));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFESR r_Clock_Count_1951__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n27767), .D(n1[1]), .R(n29148));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1951__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n27767), .D(n1[2]), .R(n29148));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1951__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n27767), .D(n1[3]), .R(n29148));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1951__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n27767), .D(n1[4]), .R(n29148));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1951__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n27767), .D(n1[5]), .R(n29148));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1951__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n27767), .D(n1[6]), .R(n29148));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1951__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n27767), .D(n1[7]), .R(n29148));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_1951__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n27767), .D(n1[0]), .R(n29148));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 div_37_i2047_3_lut (.I0(n2938), .I1(n8373[23]), .I2(n294[3]), 
            .I3(GND_net), .O(n3046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2055_3_lut (.I0(n2946), .I1(n8373[15]), .I2(n294[3]), 
            .I3(GND_net), .O(n3054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2048_3_lut (.I0(n2939), .I1(n8373[22]), .I2(n294[3]), 
            .I3(GND_net), .O(n3047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2049_3_lut (.I0(n2940), .I1(n8373[21]), .I2(n294[3]), 
            .I3(GND_net), .O(n3048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2050_3_lut (.I0(n2941), .I1(n8373[20]), .I2(n294[3]), 
            .I3(GND_net), .O(n3049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2053_3_lut (.I0(n2944), .I1(n8373[17]), .I2(n294[3]), 
            .I3(GND_net), .O(n3052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i35_2_lut (.I0(n3052), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4513));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2051_3_lut (.I0(n2942), .I1(n8373[19]), .I2(n294[3]), 
            .I3(GND_net), .O(n3050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i39_2_lut (.I0(n3050), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4514));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2054_3_lut (.I0(n2945), .I1(n8373[16]), .I2(n294[3]), 
            .I3(GND_net), .O(n3053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i33_2_lut (.I0(n3053), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4515));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2052_3_lut (.I0(n2943), .I1(n8373[18]), .I2(n294[3]), 
            .I3(GND_net), .O(n3051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i37_2_lut (.I0(n3051), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4516));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2056_3_lut (.I0(n2947), .I1(n8373[14]), .I2(n294[3]), 
            .I3(GND_net), .O(n3055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2057_3_lut (.I0(n2948), .I1(n8373[13]), .I2(n294[3]), 
            .I3(GND_net), .O(n3056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i27_2_lut (.I0(n3056), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4517));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i29_2_lut (.I0(n3055), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4518));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2058_3_lut (.I0(n2949), .I1(n8373[12]), .I2(n294[3]), 
            .I3(GND_net), .O(n3057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2059_3_lut (.I0(n2950), .I1(n8373[11]), .I2(n294[3]), 
            .I3(GND_net), .O(n3058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i23_2_lut (.I0(n3058), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4519));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i25_2_lut (.I0(n3057), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4520));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2065_3_lut (.I0(n2956), .I1(n8373[5]), .I2(n294[3]), 
            .I3(GND_net), .O(n3064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2066_3_lut (.I0(n2957), .I1(n8373[4]), .I2(n294[3]), 
            .I3(GND_net), .O(n3065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2802_25_lut (.I0(GND_net), .I1(n3151), .I2(n3186), .I3(n50386), 
            .O(n8425[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2802_24_lut (.I0(GND_net), .I1(n3152), .I2(n3082), .I3(n50385), 
            .O(n8425[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_24 (.CI(n50385), .I0(n3152), .I1(n3082), .CO(n50386));
    SB_LUT4 add_2802_23_lut (.I0(GND_net), .I1(n3153), .I2(n3188), .I3(n50384), 
            .O(n8425[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_23 (.CI(n50384), .I0(n3153), .I1(n3188), .CO(n50385));
    SB_LUT4 add_2802_22_lut (.I0(GND_net), .I1(n3154), .I2(n3084), .I3(n50383), 
            .O(n8425[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_22 (.CI(n50383), .I0(n3154), .I1(n3084), .CO(n50384));
    SB_LUT4 add_2802_21_lut (.I0(GND_net), .I1(n3155), .I2(n2977), .I3(n50382), 
            .O(n8425[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_21 (.CI(n50382), .I0(n3155), .I1(n2977), .CO(n50383));
    SB_LUT4 add_2802_20_lut (.I0(GND_net), .I1(n3156), .I2(n2867), .I3(n50381), 
            .O(n8425[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_20 (.CI(n50381), .I0(n3156), .I1(n2867), .CO(n50382));
    SB_LUT4 add_2802_19_lut (.I0(GND_net), .I1(n3157), .I2(n2754), .I3(n50380), 
            .O(n8425[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_19 (.CI(n50380), .I0(n3157), .I1(n2754), .CO(n50381));
    SB_LUT4 add_2802_18_lut (.I0(GND_net), .I1(n3158), .I2(n2638), .I3(n50379), 
            .O(n8425[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_18 (.CI(n50379), .I0(n3158), .I1(n2638), .CO(n50380));
    SB_LUT4 add_2802_17_lut (.I0(GND_net), .I1(n3159), .I2(n2519), .I3(n50378), 
            .O(n8425[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_17 (.CI(n50378), .I0(n3159), .I1(n2519), .CO(n50379));
    SB_LUT4 add_2802_16_lut (.I0(GND_net), .I1(n3160), .I2(n2397), .I3(n50377), 
            .O(n8425[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2070_i11_2_lut (.I0(n3064), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4521));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2802_16 (.CI(n50377), .I0(n3160), .I1(n2397), .CO(n50378));
    SB_LUT4 add_2802_15_lut (.I0(GND_net), .I1(n3161), .I2(n2272), .I3(n50376), 
            .O(n8425[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_15 (.CI(n50376), .I0(n3161), .I1(n2272), .CO(n50377));
    SB_LUT4 add_2802_14_lut (.I0(GND_net), .I1(n3162), .I2(n2144), .I3(n50375), 
            .O(n8425[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_14 (.CI(n50375), .I0(n3162), .I1(n2144), .CO(n50376));
    SB_LUT4 add_2802_13_lut (.I0(GND_net), .I1(n3163), .I2(n2013), .I3(n50374), 
            .O(n8425[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_13 (.CI(n50374), .I0(n3163), .I1(n2013), .CO(n50375));
    SB_LUT4 add_2802_12_lut (.I0(GND_net), .I1(n3164), .I2(n1879), .I3(n50373), 
            .O(n8425[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_12 (.CI(n50373), .I0(n3164), .I1(n1879), .CO(n50374));
    SB_LUT4 add_2802_11_lut (.I0(GND_net), .I1(n3165), .I2(n1742), .I3(n50372), 
            .O(n8425[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_11 (.CI(n50372), .I0(n3165), .I1(n1742), .CO(n50373));
    SB_LUT4 add_2802_10_lut (.I0(GND_net), .I1(n3166), .I2(n1602), .I3(n50371), 
            .O(n8425[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_10 (.CI(n50371), .I0(n3166), .I1(n1602), .CO(n50372));
    SB_LUT4 add_2802_9_lut (.I0(GND_net), .I1(n3167), .I2(n1459), .I3(n50370), 
            .O(n8425[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_9 (.CI(n50370), .I0(n3167), .I1(n1459), .CO(n50371));
    SB_LUT4 add_2802_8_lut (.I0(GND_net), .I1(n3168), .I2(n1460), .I3(n50369), 
            .O(n8425[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_8 (.CI(n50369), .I0(n3168), .I1(n1460), .CO(n50370));
    SB_LUT4 add_2802_7_lut (.I0(GND_net), .I1(n3169), .I2(n1011), .I3(n50368), 
            .O(n8425[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_7 (.CI(n50368), .I0(n3169), .I1(n1011), .CO(n50369));
    SB_LUT4 add_2802_6_lut (.I0(GND_net), .I1(n3170), .I2(n856), .I3(n50367), 
            .O(n8425[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_6 (.CI(n50367), .I0(n3170), .I1(n856), .CO(n50368));
    SB_LUT4 add_2802_5_lut (.I0(GND_net), .I1(n3171), .I2(n698), .I3(n50366), 
            .O(n8425[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_5 (.CI(n50366), .I0(n3171), .I1(n698), .CO(n50367));
    SB_LUT4 add_2802_4_lut (.I0(GND_net), .I1(n3172), .I2(n858), .I3(n50365), 
            .O(n8425[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2802_4 (.CI(n50365), .I0(n3172), .I1(n858), .CO(n50366));
    SB_LUT4 add_2802_3_lut (.I0(n58062), .I1(GND_net), .I2(n538), .I3(n50364), 
            .O(n60336)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2802_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2802_3 (.CI(n50364), .I0(GND_net), .I1(n538), .CO(n50365));
    SB_CARRY add_2802_2 (.CI(VCC_net), .I0(GND_net), .I1(VCC_net), .CO(n50364));
    SB_LUT4 add_2801_23_lut (.I0(GND_net), .I1(n3046), .I2(n3082), .I3(n50363), 
            .O(n8399[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2801_22_lut (.I0(GND_net), .I1(n3047), .I2(n3188), .I3(n50362), 
            .O(n8399[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_22 (.CI(n50362), .I0(n3047), .I1(n3188), .CO(n50363));
    SB_LUT4 div_37_i2064_3_lut (.I0(n2955), .I1(n8373[6]), .I2(n294[3]), 
            .I3(GND_net), .O(n3063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2801_21_lut (.I0(GND_net), .I1(n3048), .I2(n3084), .I3(n50361), 
            .O(n8399[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_21 (.CI(n50361), .I0(n3048), .I1(n3084), .CO(n50362));
    SB_LUT4 add_2801_20_lut (.I0(GND_net), .I1(n3049), .I2(n2977), .I3(n50360), 
            .O(n8399[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_20 (.CI(n50360), .I0(n3049), .I1(n2977), .CO(n50361));
    SB_LUT4 add_2801_19_lut (.I0(GND_net), .I1(n3050), .I2(n2867), .I3(n50359), 
            .O(n8399[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_19 (.CI(n50359), .I0(n3050), .I1(n2867), .CO(n50360));
    SB_LUT4 add_2801_18_lut (.I0(GND_net), .I1(n3051), .I2(n2754), .I3(n50358), 
            .O(n8399[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_18 (.CI(n50358), .I0(n3051), .I1(n2754), .CO(n50359));
    SB_LUT4 add_2801_17_lut (.I0(GND_net), .I1(n3052), .I2(n2638), .I3(n50357), 
            .O(n8399[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_17 (.CI(n50357), .I0(n3052), .I1(n2638), .CO(n50358));
    SB_LUT4 add_2801_16_lut (.I0(GND_net), .I1(n3053), .I2(n2519), .I3(n50356), 
            .O(n8399[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_16 (.CI(n50356), .I0(n3053), .I1(n2519), .CO(n50357));
    SB_LUT4 add_2801_15_lut (.I0(GND_net), .I1(n3054), .I2(n2397), .I3(n50355), 
            .O(n8399[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_15 (.CI(n50355), .I0(n3054), .I1(n2397), .CO(n50356));
    SB_LUT4 add_2801_14_lut (.I0(GND_net), .I1(n3055), .I2(n2272), .I3(n50354), 
            .O(n8399[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_14 (.CI(n50354), .I0(n3055), .I1(n2272), .CO(n50355));
    SB_LUT4 add_2801_13_lut (.I0(GND_net), .I1(n3056), .I2(n2144), .I3(n50353), 
            .O(n8399[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_13 (.CI(n50353), .I0(n3056), .I1(n2144), .CO(n50354));
    SB_LUT4 add_2801_12_lut (.I0(GND_net), .I1(n3057), .I2(n2013), .I3(n50352), 
            .O(n8399[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_12 (.CI(n50352), .I0(n3057), .I1(n2013), .CO(n50353));
    SB_LUT4 add_2801_11_lut (.I0(GND_net), .I1(n3058), .I2(n1879), .I3(n50351), 
            .O(n8399[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_11 (.CI(n50351), .I0(n3058), .I1(n1879), .CO(n50352));
    SB_LUT4 add_2801_10_lut (.I0(GND_net), .I1(n3059), .I2(n1742), .I3(n50350), 
            .O(n8399[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_10 (.CI(n50350), .I0(n3059), .I1(n1742), .CO(n50351));
    SB_LUT4 add_2801_9_lut (.I0(GND_net), .I1(n3060), .I2(n1602), .I3(n50349), 
            .O(n8399[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_9 (.CI(n50349), .I0(n3060), .I1(n1602), .CO(n50350));
    SB_LUT4 add_2801_8_lut (.I0(GND_net), .I1(n3061), .I2(n1459), .I3(n50348), 
            .O(n8399[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_8 (.CI(n50348), .I0(n3061), .I1(n1459), .CO(n50349));
    SB_LUT4 add_2801_7_lut (.I0(GND_net), .I1(n3062), .I2(n1460), .I3(n50347), 
            .O(n8399[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_7 (.CI(n50347), .I0(n3062), .I1(n1460), .CO(n50348));
    SB_LUT4 add_2801_6_lut (.I0(GND_net), .I1(n3063), .I2(n1011), .I3(n50346), 
            .O(n8399[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_6 (.CI(n50346), .I0(n3063), .I1(n1011), .CO(n50347));
    SB_LUT4 add_2801_5_lut (.I0(GND_net), .I1(n3064), .I2(n856), .I3(n50345), 
            .O(n8399[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_5 (.CI(n50345), .I0(n3064), .I1(n856), .CO(n50346));
    SB_LUT4 add_2801_4_lut (.I0(GND_net), .I1(n3065), .I2(n698), .I3(n50344), 
            .O(n8399[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_4 (.CI(n50344), .I0(n3065), .I1(n698), .CO(n50345));
    SB_LUT4 add_2801_3_lut (.I0(GND_net), .I1(n3066), .I2(n858), .I3(n50343), 
            .O(n8399[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2801_3 (.CI(n50343), .I0(n3066), .I1(n858), .CO(n50344));
    SB_LUT4 add_2801_2_lut (.I0(n58066), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60334)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2801_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2801_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50343));
    SB_LUT4 add_2800_22_lut (.I0(GND_net), .I1(n2938), .I2(n3188), .I3(n50342), 
            .O(n8373[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2800_21_lut (.I0(GND_net), .I1(n2939), .I2(n3084), .I3(n50341), 
            .O(n8373[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_21 (.CI(n50341), .I0(n2939), .I1(n3084), .CO(n50342));
    SB_LUT4 add_2800_20_lut (.I0(GND_net), .I1(n2940), .I2(n2977), .I3(n50340), 
            .O(n8373[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2060_3_lut (.I0(n2951), .I1(n8373[10]), .I2(n294[3]), 
            .I3(GND_net), .O(n3059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2800_20 (.CI(n50340), .I0(n2940), .I1(n2977), .CO(n50341));
    SB_LUT4 add_2800_19_lut (.I0(GND_net), .I1(n2941), .I2(n2867), .I3(n50339), 
            .O(n8373[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_19 (.CI(n50339), .I0(n2941), .I1(n2867), .CO(n50340));
    SB_LUT4 add_2800_18_lut (.I0(GND_net), .I1(n2942), .I2(n2754), .I3(n50338), 
            .O(n8373[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_18 (.CI(n50338), .I0(n2942), .I1(n2754), .CO(n50339));
    SB_LUT4 add_2800_17_lut (.I0(GND_net), .I1(n2943), .I2(n2638), .I3(n50337), 
            .O(n8373[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_17 (.CI(n50337), .I0(n2943), .I1(n2638), .CO(n50338));
    SB_LUT4 add_2800_16_lut (.I0(GND_net), .I1(n2944), .I2(n2519), .I3(n50336), 
            .O(n8373[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_16 (.CI(n50336), .I0(n2944), .I1(n2519), .CO(n50337));
    SB_LUT4 add_2800_15_lut (.I0(GND_net), .I1(n2945), .I2(n2397), .I3(n50335), 
            .O(n8373[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_15 (.CI(n50335), .I0(n2945), .I1(n2397), .CO(n50336));
    SB_LUT4 add_2800_14_lut (.I0(GND_net), .I1(n2946), .I2(n2272), .I3(n50334), 
            .O(n8373[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_14 (.CI(n50334), .I0(n2946), .I1(n2272), .CO(n50335));
    SB_LUT4 add_2800_13_lut (.I0(GND_net), .I1(n2947), .I2(n2144), .I3(n50333), 
            .O(n8373[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_13 (.CI(n50333), .I0(n2947), .I1(n2144), .CO(n50334));
    SB_LUT4 add_2800_12_lut (.I0(GND_net), .I1(n2948), .I2(n2013), .I3(n50332), 
            .O(n8373[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_12 (.CI(n50332), .I0(n2948), .I1(n2013), .CO(n50333));
    SB_LUT4 add_2800_11_lut (.I0(GND_net), .I1(n2949), .I2(n1879), .I3(n50331), 
            .O(n8373[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_11 (.CI(n50331), .I0(n2949), .I1(n1879), .CO(n50332));
    SB_LUT4 add_2800_10_lut (.I0(GND_net), .I1(n2950), .I2(n1742), .I3(n50330), 
            .O(n8373[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_10 (.CI(n50330), .I0(n2950), .I1(n1742), .CO(n50331));
    SB_LUT4 add_2800_9_lut (.I0(GND_net), .I1(n2951), .I2(n1602), .I3(n50329), 
            .O(n8373[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_9 (.CI(n50329), .I0(n2951), .I1(n1602), .CO(n50330));
    SB_LUT4 add_2800_8_lut (.I0(GND_net), .I1(n2952), .I2(n1459), .I3(n50328), 
            .O(n8373[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_8 (.CI(n50328), .I0(n2952), .I1(n1459), .CO(n50329));
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk16MHz), .D(n30502));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2800_7_lut (.I0(GND_net), .I1(n2953), .I2(n1460), .I3(n50327), 
            .O(n8373[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFE r_Rx_DV_58 (.Q(rx_data_ready), .C(clk16MHz), .E(VCC_net), 
            .D(n52851));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFFE r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .E(VCC_net), 
            .D(n30498));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_2070_i13_2_lut (.I0(n3063), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4522));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2800_7 (.CI(n50327), .I0(n2953), .I1(n1460), .CO(n50328));
    SB_LUT4 add_2800_6_lut (.I0(GND_net), .I1(n2954), .I2(n1011), .I3(n50326), 
            .O(n8373[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_6 (.CI(n50326), .I0(n2954), .I1(n1011), .CO(n50327));
    SB_LUT4 add_2800_5_lut (.I0(GND_net), .I1(n2955), .I2(n856), .I3(n50325), 
            .O(n8373[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_5 (.CI(n50325), .I0(n2955), .I1(n856), .CO(n50326));
    SB_LUT4 add_2800_4_lut (.I0(GND_net), .I1(n2956), .I2(n698), .I3(n50324), 
            .O(n8373[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_4 (.CI(n50324), .I0(n2956), .I1(n698), .CO(n50325));
    SB_LUT4 add_2800_3_lut (.I0(GND_net), .I1(n2957), .I2(n858), .I3(n50323), 
            .O(n8373[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2800_3 (.CI(n50323), .I0(n2957), .I1(n858), .CO(n50324));
    SB_LUT4 add_2800_2_lut (.I0(n58070), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60332)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2800_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2800_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50323));
    SB_LUT4 i1_3_lut_4_lut_adj_1016 (.I0(baudrate[2]), .I1(n42_adj_4462), 
            .I2(baudrate[3]), .I3(n20921), .O(n58597));   // verilog/uart_rx.v(119[33:55])
    defparam i1_3_lut_4_lut_adj_1016.LUT_INIT = 16'hff4f;
    SB_LUT4 add_2799_21_lut (.I0(GND_net), .I1(n2827), .I2(n3084), .I3(n50322), 
            .O(n8347[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2070_i21_2_lut (.I0(n3059), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4523));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2799_20_lut (.I0(GND_net), .I1(n2828), .I2(n2977), .I3(n50321), 
            .O(n8347[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i2061_3_lut (.I0(n2952), .I1(n8373[9]), .I2(n294[3]), 
            .I3(GND_net), .O(n3060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2799_20 (.CI(n50321), .I0(n2828), .I1(n2977), .CO(n50322));
    SB_LUT4 add_2799_19_lut (.I0(GND_net), .I1(n2829), .I2(n2867), .I3(n50320), 
            .O(n8347[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_19 (.CI(n50320), .I0(n2829), .I1(n2867), .CO(n50321));
    SB_LUT4 add_2799_18_lut (.I0(GND_net), .I1(n2830), .I2(n2754), .I3(n50319), 
            .O(n8347[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_18 (.CI(n50319), .I0(n2830), .I1(n2754), .CO(n50320));
    SB_LUT4 i5585_2_lut_3_lut (.I0(baudrate[2]), .I1(n42_adj_4462), .I2(n20921), 
            .I3(GND_net), .O(n44_adj_4463));   // verilog/uart_rx.v(119[33:55])
    defparam i5585_2_lut_3_lut.LUT_INIT = 16'hf4f4;
    SB_LUT4 div_37_i2062_3_lut (.I0(n2953), .I1(n8373[8]), .I2(n294[3]), 
            .I3(GND_net), .O(n3061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2063_3_lut (.I0(n2954), .I1(n8373[7]), .I2(n294[3]), 
            .I3(GND_net), .O(n3062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2799_17_lut (.I0(GND_net), .I1(n2831), .I2(n2638), .I3(n50318), 
            .O(n8347[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_17 (.CI(n50318), .I0(n2831), .I1(n2638), .CO(n50319));
    SB_LUT4 add_2799_16_lut (.I0(GND_net), .I1(n2832), .I2(n2519), .I3(n50317), 
            .O(n8347[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2070_i15_2_lut (.I0(n3062), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4524));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2799_16 (.CI(n50317), .I0(n2832), .I1(n2519), .CO(n50318));
    SB_LUT4 add_2799_15_lut (.I0(GND_net), .I1(n2833), .I2(n2397), .I3(n50316), 
            .O(n8347[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_15 (.CI(n50316), .I0(n2833), .I1(n2397), .CO(n50317));
    SB_LUT4 div_37_LessThan_2070_i17_2_lut (.I0(n3061), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4525));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2799_14_lut (.I0(GND_net), .I1(n2834), .I2(n2272), .I3(n50315), 
            .O(n8347[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_14 (.CI(n50315), .I0(n2834), .I1(n2272), .CO(n50316));
    SB_LUT4 add_2799_13_lut (.I0(GND_net), .I1(n2835), .I2(n2144), .I3(n50314), 
            .O(n8347[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_13 (.CI(n50314), .I0(n2835), .I1(n2144), .CO(n50315));
    SB_LUT4 add_2799_12_lut (.I0(GND_net), .I1(n2836), .I2(n2013), .I3(n50313), 
            .O(n8347[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_2070_i19_2_lut (.I0(n3060), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4526));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i31_2_lut (.I0(n3054), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4527));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2799_12 (.CI(n50313), .I0(n2836), .I1(n2013), .CO(n50314));
    SB_LUT4 add_2799_11_lut (.I0(GND_net), .I1(n2837), .I2(n1879), .I3(n50312), 
            .O(n8347[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_11 (.CI(n50312), .I0(n2837), .I1(n1879), .CO(n50313));
    SB_LUT4 add_2799_10_lut (.I0(GND_net), .I1(n2838), .I2(n1742), .I3(n50311), 
            .O(n8347[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_10 (.CI(n50311), .I0(n2838), .I1(n1742), .CO(n50312));
    SB_LUT4 add_2799_9_lut (.I0(GND_net), .I1(n2839), .I2(n1602), .I3(n50310), 
            .O(n8347[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_9 (.CI(n50310), .I0(n2839), .I1(n1602), .CO(n50311));
    SB_LUT4 add_2799_8_lut (.I0(GND_net), .I1(n2840), .I2(n1459), .I3(n50309), 
            .O(n8347[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_8 (.CI(n50309), .I0(n2840), .I1(n1459), .CO(n50310));
    SB_LUT4 i50056_4_lut (.I0(n31_adj_4527), .I1(n19_adj_4526), .I2(n17_adj_4525), 
            .I3(n15_adj_4524), .O(n65742));
    defparam i50056_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2799_7_lut (.I0(GND_net), .I1(n2841), .I2(n1460), .I3(n50308), 
            .O(n8347[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_7 (.CI(n50308), .I0(n2841), .I1(n1460), .CO(n50309));
    SB_LUT4 add_2799_6_lut (.I0(GND_net), .I1(n2842), .I2(n1011), .I3(n50307), 
            .O(n8347[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_6 (.CI(n50307), .I0(n2842), .I1(n1011), .CO(n50308));
    SB_LUT4 add_2799_5_lut (.I0(GND_net), .I1(n2843), .I2(n856), .I3(n50306), 
            .O(n8347[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut_adj_1017 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n60776));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1017.LUT_INIT = 16'hfffd;
    SB_CARRY add_2799_5 (.CI(n50306), .I0(n2843), .I1(n856), .CO(n50307));
    SB_LUT4 add_2799_4_lut (.I0(GND_net), .I1(n2844), .I2(n698), .I3(n50305), 
            .O(n8347[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_4 (.CI(n50305), .I0(n2844), .I1(n698), .CO(n50306));
    SB_LUT4 add_2799_3_lut (.I0(GND_net), .I1(n2845), .I2(n858), .I3(n50304), 
            .O(n8347[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2799_3 (.CI(n50304), .I0(n2845), .I1(n858), .CO(n50305));
    SB_LUT4 add_2799_2_lut (.I0(n58074), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60330)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2799_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2799_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50304));
    SB_LUT4 add_2798_20_lut (.I0(GND_net), .I1(n2713), .I2(n2977), .I3(n50303), 
            .O(n8321[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50983_4_lut (.I0(n13_adj_4522), .I1(n11_adj_4521), .I2(n3065), 
            .I3(baudrate[2]), .O(n66669));
    defparam i50983_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 add_2798_19_lut (.I0(GND_net), .I1(n2714), .I2(n2867), .I3(n50302), 
            .O(n8321[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_19 (.CI(n50302), .I0(n2714), .I1(n2867), .CO(n50303));
    SB_LUT4 add_2798_18_lut (.I0(GND_net), .I1(n2715), .I2(n2754), .I3(n50301), 
            .O(n8321[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_18 (.CI(n50301), .I0(n2715), .I1(n2754), .CO(n50302));
    SB_LUT4 i51637_4_lut (.I0(n19_adj_4526), .I1(n17_adj_4525), .I2(n15_adj_4524), 
            .I3(n66669), .O(n67323));
    defparam i51637_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51635_4_lut (.I0(n25_adj_4520), .I1(n23_adj_4519), .I2(n21_adj_4523), 
            .I3(n67323), .O(n67321));
    defparam i51635_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50058_4_lut (.I0(n31_adj_4527), .I1(n29_adj_4518), .I2(n27_adj_4517), 
            .I3(n67321), .O(n65744));
    defparam i50058_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2798_17_lut (.I0(GND_net), .I1(n2716), .I2(n2638), .I3(n50300), 
            .O(n8321[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_17 (.CI(n50300), .I0(n2716), .I1(n2638), .CO(n50301));
    SB_LUT4 add_2798_16_lut (.I0(GND_net), .I1(n2717), .I2(n2519), .I3(n50299), 
            .O(n8321[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_16 (.CI(n50299), .I0(n2717), .I1(n2519), .CO(n50300));
    SB_LUT4 add_2798_15_lut (.I0(GND_net), .I1(n2718), .I2(n2397), .I3(n50298), 
            .O(n8321[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_15 (.CI(n50298), .I0(n2718), .I1(n2397), .CO(n50299));
    SB_LUT4 div_37_LessThan_2070_i8_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3066), .I3(GND_net), .O(n8_adj_4528));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2798_14_lut (.I0(GND_net), .I1(n2719), .I2(n2272), .I3(n50297), 
            .O(n8321[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52139_3_lut (.I0(n8_adj_4528), .I1(baudrate[13]), .I2(n31_adj_4527), 
            .I3(GND_net), .O(n67825));   // verilog/uart_rx.v(119[33:55])
    defparam i52139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52140_3_lut (.I0(n67825), .I1(baudrate[14]), .I2(n33_adj_4515), 
            .I3(GND_net), .O(n67826));   // verilog/uart_rx.v(119[33:55])
    defparam i52140_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2798_14 (.CI(n50297), .I0(n2719), .I1(n2272), .CO(n50298));
    SB_LUT4 add_2798_13_lut (.I0(GND_net), .I1(n2720), .I2(n2144), .I3(n50296), 
            .O(n8321[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_13 (.CI(n50296), .I0(n2720), .I1(n2144), .CO(n50297));
    SB_LUT4 add_2798_12_lut (.I0(GND_net), .I1(n2721), .I2(n2013), .I3(n50295), 
            .O(n8321[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk16MHz), .D(n30201));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk16MHz), .D(n30200));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2798_12 (.CI(n50295), .I0(n2721), .I1(n2013), .CO(n50296));
    SB_LUT4 add_2798_11_lut (.I0(GND_net), .I1(n2722), .I2(n1879), .I3(n50294), 
            .O(n8321[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_11 (.CI(n50294), .I0(n2722), .I1(n1879), .CO(n50295));
    SB_LUT4 add_2798_10_lut (.I0(GND_net), .I1(n2723), .I2(n1742), .I3(n50293), 
            .O(n8321[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_10 (.CI(n50293), .I0(n2723), .I1(n1742), .CO(n50294));
    SB_LUT4 add_2798_9_lut (.I0(GND_net), .I1(n2724), .I2(n1602), .I3(n50292), 
            .O(n8321[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_9 (.CI(n50292), .I0(n2724), .I1(n1602), .CO(n50293));
    SB_LUT4 add_2798_8_lut (.I0(GND_net), .I1(n2725), .I2(n1459), .I3(n50291), 
            .O(n8321[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_8 (.CI(n50291), .I0(n2725), .I1(n1459), .CO(n50292));
    SB_LUT4 add_2798_7_lut (.I0(GND_net), .I1(n2726), .I2(n1460), .I3(n50290), 
            .O(n8321[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_7 (.CI(n50290), .I0(n2726), .I1(n1460), .CO(n50291));
    SB_LUT4 add_2798_6_lut (.I0(GND_net), .I1(n2727), .I2(n1011), .I3(n50289), 
            .O(n8321[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_6 (.CI(n50289), .I0(n2727), .I1(n1011), .CO(n50290));
    SB_LUT4 add_2798_5_lut (.I0(GND_net), .I1(n2728), .I2(n856), .I3(n50288), 
            .O(n8321[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_5 (.CI(n50288), .I0(n2728), .I1(n856), .CO(n50289));
    SB_LUT4 add_2798_4_lut (.I0(GND_net), .I1(n2729), .I2(n698), .I3(n50287), 
            .O(n8321[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_4 (.CI(n50287), .I0(n2729), .I1(n698), .CO(n50288));
    SB_LUT4 add_2798_3_lut (.I0(GND_net), .I1(n2730), .I2(n858), .I3(n50286), 
            .O(n8321[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2798_3 (.CI(n50286), .I0(n2730), .I1(n858), .CO(n50287));
    SB_LUT4 div_37_LessThan_2070_i34_3_lut (.I0(n16_adj_4529), .I1(baudrate[17]), 
            .I2(n39_adj_4514), .I3(GND_net), .O(n34_adj_4530));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2798_2_lut (.I0(n58078), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60328)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2798_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2798_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50286));
    SB_LUT4 add_2797_19_lut (.I0(GND_net), .I1(n2596), .I2(n2867), .I3(n50285), 
            .O(n8295[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2797_18_lut (.I0(GND_net), .I1(n2597), .I2(n2754), .I3(n50284), 
            .O(n8295[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_18 (.CI(n50284), .I0(n2597), .I1(n2754), .CO(n50285));
    SB_LUT4 add_2797_17_lut (.I0(GND_net), .I1(n2598), .I2(n2638), .I3(n50283), 
            .O(n8295[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_17 (.CI(n50283), .I0(n2598), .I1(n2638), .CO(n50284));
    SB_LUT4 add_2797_16_lut (.I0(GND_net), .I1(n2599), .I2(n2519), .I3(n50282), 
            .O(n8295[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_16 (.CI(n50282), .I0(n2599), .I1(n2519), .CO(n50283));
    SB_LUT4 add_2797_15_lut (.I0(GND_net), .I1(n2600), .I2(n2397), .I3(n50281), 
            .O(n8295[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_15 (.CI(n50281), .I0(n2600), .I1(n2397), .CO(n50282));
    SB_LUT4 add_2797_14_lut (.I0(GND_net), .I1(n2601), .I2(n2272), .I3(n50280), 
            .O(n8295[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_14 (.CI(n50280), .I0(n2601), .I1(n2272), .CO(n50281));
    SB_LUT4 add_2797_13_lut (.I0(GND_net), .I1(n2602), .I2(n2144), .I3(n50279), 
            .O(n8295[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_13 (.CI(n50279), .I0(n2602), .I1(n2144), .CO(n50280));
    SB_LUT4 add_2797_12_lut (.I0(GND_net), .I1(n2603), .I2(n2013), .I3(n50278), 
            .O(n8295[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i50048_4_lut (.I0(n37_adj_4516), .I1(n35_adj_4513), .I2(n33_adj_4515), 
            .I3(n65742), .O(n65734));
    defparam i50048_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2797_12 (.CI(n50278), .I0(n2603), .I1(n2013), .CO(n50279));
    SB_LUT4 add_2797_11_lut (.I0(GND_net), .I1(n2604), .I2(n1879), .I3(n50277), 
            .O(n8295[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_11 (.CI(n50277), .I0(n2604), .I1(n1879), .CO(n50278));
    SB_LUT4 add_2797_10_lut (.I0(GND_net), .I1(n2605), .I2(n1742), .I3(n50276), 
            .O(n8295[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52479_4_lut (.I0(n34_adj_4530), .I1(n14_adj_4531), .I2(n39_adj_4514), 
            .I3(n65728), .O(n68165));   // verilog/uart_rx.v(119[33:55])
    defparam i52479_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2797_10 (.CI(n50276), .I0(n2605), .I1(n1742), .CO(n50277));
    SB_LUT4 i52052_3_lut (.I0(n67826), .I1(baudrate[15]), .I2(n35_adj_4513), 
            .I3(GND_net), .O(n67738));   // verilog/uart_rx.v(119[33:55])
    defparam i52052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2797_9_lut (.I0(GND_net), .I1(n2606), .I2(n1602), .I3(n50275), 
            .O(n8295[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_9 (.CI(n50275), .I0(n2606), .I1(n1602), .CO(n50276));
    SB_LUT4 i52141_3_lut (.I0(n10_adj_4532), .I1(baudrate[10]), .I2(n25_adj_4520), 
            .I3(GND_net), .O(n67827));   // verilog/uart_rx.v(119[33:55])
    defparam i52141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52142_3_lut (.I0(n67827), .I1(baudrate[11]), .I2(n27_adj_4517), 
            .I3(GND_net), .O(n67828));   // verilog/uart_rx.v(119[33:55])
    defparam i52142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2797_8_lut (.I0(GND_net), .I1(n2607), .I2(n1459), .I3(n50274), 
            .O(n8295[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_8 (.CI(n50274), .I0(n2607), .I1(n1459), .CO(n50275));
    SB_LUT4 i50971_4_lut (.I0(n27_adj_4517), .I1(n25_adj_4520), .I2(n23_adj_4519), 
            .I3(n65757), .O(n66657));
    defparam i50971_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_2797_7_lut (.I0(GND_net), .I1(n2608), .I2(n1460), .I3(n50273), 
            .O(n8295[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_7 (.CI(n50273), .I0(n2608), .I1(n1460), .CO(n50274));
    SB_LUT4 div_37_LessThan_2070_i20_3_lut (.I0(n12_adj_4533), .I1(baudrate[9]), 
            .I2(n23_adj_4519), .I3(GND_net), .O(n20));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2797_6_lut (.I0(GND_net), .I1(n2609), .I2(n1011), .I3(n50272), 
            .O(n8295[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_6 (.CI(n50272), .I0(n2609), .I1(n1011), .CO(n50273));
    SB_LUT4 add_2797_5_lut (.I0(GND_net), .I1(n2610), .I2(n856), .I3(n50271), 
            .O(n8295[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_5 (.CI(n50271), .I0(n2610), .I1(n856), .CO(n50272));
    SB_LUT4 add_2797_4_lut (.I0(GND_net), .I1(n2611), .I2(n698), .I3(n50270), 
            .O(n8295[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2797_4 (.CI(n50270), .I0(n2611), .I1(n698), .CO(n50271));
    SB_LUT4 i52050_3_lut (.I0(n67828), .I1(baudrate[12]), .I2(n29_adj_4518), 
            .I3(GND_net), .O(n26));   // verilog/uart_rx.v(119[33:55])
    defparam i52050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2797_3_lut (.I0(GND_net), .I1(n2612), .I2(n858), .I3(n50269), 
            .O(n8295[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51948_4_lut (.I0(n37_adj_4516), .I1(n35_adj_4513), .I2(n33_adj_4515), 
            .I3(n65744), .O(n67634));
    defparam i51948_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_2797_3 (.CI(n50269), .I0(n2612), .I1(n858), .CO(n50270));
    SB_LUT4 i52605_4_lut (.I0(n67738), .I1(n68165), .I2(n39_adj_4514), 
            .I3(n65734), .O(n68291));   // verilog/uart_rx.v(119[33:55])
    defparam i52605_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2797_2_lut (.I0(n58082), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60326)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2797_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2797_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50269));
    SB_LUT4 add_2796_18_lut (.I0(GND_net), .I1(n2476), .I2(n2754), .I3(n50268), 
            .O(n8269[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2796_17_lut (.I0(GND_net), .I1(n2477), .I2(n2638), .I3(n50267), 
            .O(n8269[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_17 (.CI(n50267), .I0(n2477), .I1(n2638), .CO(n50268));
    SB_LUT4 i51703_4_lut (.I0(n26), .I1(n20), .I2(n29_adj_4518), .I3(n66657), 
            .O(n67389));   // verilog/uart_rx.v(119[33:55])
    defparam i51703_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2796_16_lut (.I0(GND_net), .I1(n2478), .I2(n2519), .I3(n50266), 
            .O(n8269[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_16 (.CI(n50266), .I0(n2478), .I1(n2519), .CO(n50267));
    SB_LUT4 add_2796_15_lut (.I0(GND_net), .I1(n2479), .I2(n2397), .I3(n50265), 
            .O(n8269[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_15 (.CI(n50265), .I0(n2479), .I1(n2397), .CO(n50266));
    SB_LUT4 add_2796_14_lut (.I0(GND_net), .I1(n2480), .I2(n2272), .I3(n50264), 
            .O(n8269[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_14 (.CI(n50264), .I0(n2480), .I1(n2272), .CO(n50265));
    SB_LUT4 add_2796_13_lut (.I0(GND_net), .I1(n2481), .I2(n2144), .I3(n50263), 
            .O(n8269[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_13 (.CI(n50263), .I0(n2481), .I1(n2144), .CO(n50264));
    SB_LUT4 add_2796_12_lut (.I0(GND_net), .I1(n2482), .I2(n2013), .I3(n50262), 
            .O(n8269[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_12 (.CI(n50262), .I0(n2482), .I1(n2013), .CO(n50263));
    SB_LUT4 i52631_4_lut (.I0(n67389), .I1(n68291), .I2(n39_adj_4514), 
            .I3(n67634), .O(n68317));   // verilog/uart_rx.v(119[33:55])
    defparam i52631_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2796_11_lut (.I0(GND_net), .I1(n2483), .I2(n1879), .I3(n50261), 
            .O(n8269[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_11 (.CI(n50261), .I0(n2483), .I1(n1879), .CO(n50262));
    SB_LUT4 add_2796_10_lut (.I0(GND_net), .I1(n2484), .I2(n1742), .I3(n50260), 
            .O(n8269[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_10 (.CI(n50260), .I0(n2484), .I1(n1742), .CO(n50261));
    SB_LUT4 add_2796_9_lut (.I0(GND_net), .I1(n2485), .I2(n1602), .I3(n50259), 
            .O(n8269[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_9 (.CI(n50259), .I0(n2485), .I1(n1602), .CO(n50260));
    SB_LUT4 add_2796_8_lut (.I0(GND_net), .I1(n2486), .I2(n1459), .I3(n50258), 
            .O(n8269[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_8 (.CI(n50258), .I0(n2486), .I1(n1459), .CO(n50259));
    SB_LUT4 add_2796_7_lut (.I0(GND_net), .I1(n2487), .I2(n1460), .I3(n50257), 
            .O(n8269[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_7 (.CI(n50257), .I0(n2487), .I1(n1460), .CO(n50258));
    SB_LUT4 add_2796_6_lut (.I0(GND_net), .I1(n2488), .I2(n1011), .I3(n50256), 
            .O(n8269[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_6 (.CI(n50256), .I0(n2488), .I1(n1011), .CO(n50257));
    SB_LUT4 add_2796_5_lut (.I0(GND_net), .I1(n2489), .I2(n856), .I3(n50255), 
            .O(n8269[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_5 (.CI(n50255), .I0(n2489), .I1(n856), .CO(n50256));
    SB_LUT4 add_2796_4_lut (.I0(GND_net), .I1(n2490), .I2(n698), .I3(n50254), 
            .O(n8269[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_4 (.CI(n50254), .I0(n2490), .I1(n698), .CO(n50255));
    SB_LUT4 add_2796_3_lut (.I0(GND_net), .I1(n2491), .I2(n858), .I3(n50253), 
            .O(n8269[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2796_3 (.CI(n50253), .I0(n2491), .I1(n858), .CO(n50254));
    SB_LUT4 add_2796_2_lut (.I0(n58086), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60324)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2796_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2796_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50253));
    SB_LUT4 add_2795_17_lut (.I0(GND_net), .I1(n2353), .I2(n2638), .I3(n50252), 
            .O(n8243[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2795_16_lut (.I0(GND_net), .I1(n2354), .I2(n2519), .I3(n50251), 
            .O(n8243[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_16 (.CI(n50251), .I0(n2354), .I1(n2519), .CO(n50252));
    SB_LUT4 add_2795_15_lut (.I0(GND_net), .I1(n2355), .I2(n2397), .I3(n50250), 
            .O(n8243[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_15 (.CI(n50250), .I0(n2355), .I1(n2397), .CO(n50251));
    SB_LUT4 add_2795_14_lut (.I0(GND_net), .I1(n2356), .I2(n2272), .I3(n50249), 
            .O(n8243[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_14 (.CI(n50249), .I0(n2356), .I1(n2272), .CO(n50250));
    SB_LUT4 add_2795_13_lut (.I0(GND_net), .I1(n2357), .I2(n2144), .I3(n50248), 
            .O(n8243[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_13 (.CI(n50248), .I0(n2357), .I1(n2144), .CO(n50249));
    SB_LUT4 add_2795_12_lut (.I0(GND_net), .I1(n2358), .I2(n2013), .I3(n50247), 
            .O(n8243[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_12 (.CI(n50247), .I0(n2358), .I1(n2013), .CO(n50248));
    SB_LUT4 add_2795_11_lut (.I0(GND_net), .I1(n2359), .I2(n1879), .I3(n50246), 
            .O(n8243[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_11 (.CI(n50246), .I0(n2359), .I1(n1879), .CO(n50247));
    SB_LUT4 add_2795_10_lut (.I0(GND_net), .I1(n2360), .I2(n1742), .I3(n50245), 
            .O(n8243[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_10 (.CI(n50245), .I0(n2360), .I1(n1742), .CO(n50246));
    SB_LUT4 add_2795_9_lut (.I0(GND_net), .I1(n2361), .I2(n1602), .I3(n50244), 
            .O(n8243[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_9 (.CI(n50244), .I0(n2361), .I1(n1602), .CO(n50245));
    SB_LUT4 add_2795_8_lut (.I0(GND_net), .I1(n2362), .I2(n1459), .I3(n50243), 
            .O(n8243[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_8 (.CI(n50243), .I0(n2362), .I1(n1459), .CO(n50244));
    SB_LUT4 add_2795_7_lut (.I0(GND_net), .I1(n2363), .I2(n1460), .I3(n50242), 
            .O(n8243[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_7 (.CI(n50242), .I0(n2363), .I1(n1460), .CO(n50243));
    SB_LUT4 add_2795_6_lut (.I0(GND_net), .I1(n2364), .I2(n1011), .I3(n50241), 
            .O(n8243[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_6 (.CI(n50241), .I0(n2364), .I1(n1011), .CO(n50242));
    SB_LUT4 add_2795_5_lut (.I0(GND_net), .I1(n2365), .I2(n856), .I3(n50240), 
            .O(n8243[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_5 (.CI(n50240), .I0(n2365), .I1(n856), .CO(n50241));
    SB_LUT4 add_2795_4_lut (.I0(GND_net), .I1(n2366), .I2(n698), .I3(n50239), 
            .O(n8243[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_4 (.CI(n50239), .I0(n2366), .I1(n698), .CO(n50240));
    SB_LUT4 i52632_3_lut (.I0(n68317), .I1(baudrate[18]), .I2(n3049), 
            .I3(GND_net), .O(n68318));   // verilog/uart_rx.v(119[33:55])
    defparam i52632_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52618_3_lut (.I0(n68318), .I1(baudrate[19]), .I2(n3048), 
            .I3(GND_net), .O(n68304));   // verilog/uart_rx.v(119[33:55])
    defparam i52618_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51705_3_lut (.I0(n68304), .I1(baudrate[20]), .I2(n3047), 
            .I3(GND_net), .O(n67391));   // verilog/uart_rx.v(119[33:55])
    defparam i51705_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2795_3_lut (.I0(GND_net), .I1(n2367), .I2(n858), .I3(n50238), 
            .O(n8243[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2795_3 (.CI(n50238), .I0(n2367), .I1(n858), .CO(n50239));
    SB_LUT4 add_2795_2_lut (.I0(n58090), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60322)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2795_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2795_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50238));
    SB_LUT4 add_2794_16_lut (.I0(GND_net), .I1(n2227), .I2(n2519), .I3(n50237), 
            .O(n8217[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2794_15_lut (.I0(GND_net), .I1(n2228), .I2(n2397), .I3(n50236), 
            .O(n8217[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_15 (.CI(n50236), .I0(n2228), .I1(n2397), .CO(n50237));
    SB_LUT4 add_2794_14_lut (.I0(GND_net), .I1(n2229), .I2(n2272), .I3(n50235), 
            .O(n8217[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_14 (.CI(n50235), .I0(n2229), .I1(n2272), .CO(n50236));
    SB_LUT4 div_37_i1974_3_lut (.I0(n2827), .I1(n8347[23]), .I2(n294[4]), 
            .I3(GND_net), .O(n2938));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2794_13_lut (.I0(GND_net), .I1(n2230), .I2(n2144), .I3(n50234), 
            .O(n8217[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_13 (.CI(n50234), .I0(n2230), .I1(n2144), .CO(n50235));
    SB_LUT4 div_37_i1975_3_lut (.I0(n2828), .I1(n8347[22]), .I2(n294[4]), 
            .I3(GND_net), .O(n2939));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1990_3_lut (.I0(n2843), .I1(n8347[7]), .I2(n294[4]), 
            .I3(GND_net), .O(n2954));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2794_12_lut (.I0(GND_net), .I1(n2231), .I2(n2013), .I3(n50233), 
            .O(n8217[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1976_3_lut (.I0(n2829), .I1(n8347[21]), .I2(n294[4]), 
            .I3(GND_net), .O(n2940));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1976_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2794_12 (.CI(n50233), .I0(n2231), .I1(n2013), .CO(n50234));
    SB_LUT4 div_37_i1979_3_lut (.I0(n2832), .I1(n8347[18]), .I2(n294[4]), 
            .I3(GND_net), .O(n2943));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i37_2_lut (.I0(n2943), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4534));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2794_11_lut (.I0(GND_net), .I1(n2232), .I2(n1879), .I3(n50232), 
            .O(n8217[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_11 (.CI(n50232), .I0(n2232), .I1(n1879), .CO(n50233));
    SB_LUT4 div_37_i1977_3_lut (.I0(n2830), .I1(n8347[20]), .I2(n294[4]), 
            .I3(GND_net), .O(n2941));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2794_10_lut (.I0(GND_net), .I1(n2233), .I2(n1742), .I3(n50231), 
            .O(n8217[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_10 (.CI(n50231), .I0(n2233), .I1(n1742), .CO(n50232));
    SB_LUT4 add_2794_9_lut (.I0(GND_net), .I1(n2234), .I2(n1602), .I3(n50230), 
            .O(n8217[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_9 (.CI(n50230), .I0(n2234), .I1(n1602), .CO(n50231));
    SB_LUT4 add_2794_8_lut (.I0(GND_net), .I1(n2235), .I2(n1459), .I3(n50229), 
            .O(n8217[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i41_2_lut (.I0(n2941), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4535));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2794_8 (.CI(n50229), .I0(n2235), .I1(n1459), .CO(n50230));
    SB_LUT4 add_2794_7_lut (.I0(GND_net), .I1(n2236), .I2(n1460), .I3(n50228), 
            .O(n8217[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_7 (.CI(n50228), .I0(n2236), .I1(n1460), .CO(n50229));
    SB_LUT4 add_2794_6_lut (.I0(GND_net), .I1(n2237), .I2(n1011), .I3(n50227), 
            .O(n8217[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_6 (.CI(n50227), .I0(n2237), .I1(n1011), .CO(n50228));
    SB_LUT4 add_2794_5_lut (.I0(GND_net), .I1(n2238), .I2(n856), .I3(n50226), 
            .O(n8217[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_5 (.CI(n50226), .I0(n2238), .I1(n856), .CO(n50227));
    SB_LUT4 add_2794_4_lut (.I0(GND_net), .I1(n2239), .I2(n698), .I3(n50225), 
            .O(n8217[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_4 (.CI(n50225), .I0(n2239), .I1(n698), .CO(n50226));
    SB_LUT4 add_2794_3_lut (.I0(GND_net), .I1(n2240), .I2(n858), .I3(n50224), 
            .O(n8217[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2794_3 (.CI(n50224), .I0(n2240), .I1(n858), .CO(n50225));
    SB_LUT4 add_2794_2_lut (.I0(n58094), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60320)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2794_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2794_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50224));
    SB_LUT4 add_2793_14_lut (.I0(GND_net), .I1(n2098), .I2(n2397), .I3(n50223), 
            .O(n8191[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2793_13_lut (.I0(GND_net), .I1(n2099), .I2(n2272), .I3(n50222), 
            .O(n8191[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_13 (.CI(n50222), .I0(n2099), .I1(n2272), .CO(n50223));
    SB_LUT4 add_2793_12_lut (.I0(GND_net), .I1(n2100), .I2(n2144), .I3(n50221), 
            .O(n8191[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_12 (.CI(n50221), .I0(n2100), .I1(n2144), .CO(n50222));
    SB_LUT4 add_2793_11_lut (.I0(GND_net), .I1(n2101), .I2(n2013), .I3(n50220), 
            .O(n8191[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_11 (.CI(n50220), .I0(n2101), .I1(n2013), .CO(n50221));
    SB_LUT4 add_2793_10_lut (.I0(GND_net), .I1(n2102), .I2(n1879), .I3(n50219), 
            .O(n8191[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut_adj_1018 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n60744));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1018.LUT_INIT = 16'hffdf;
    SB_CARRY add_2793_10 (.CI(n50219), .I0(n2102), .I1(n1879), .CO(n50220));
    SB_LUT4 add_2793_9_lut (.I0(GND_net), .I1(n2103), .I2(n1742), .I3(n50218), 
            .O(n8191[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_9 (.CI(n50218), .I0(n2103), .I1(n1742), .CO(n50219));
    SB_LUT4 div_37_i1980_3_lut (.I0(n2833), .I1(n8347[17]), .I2(n294[4]), 
            .I3(GND_net), .O(n2944));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i35_2_lut (.I0(n2944), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4536));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2793_8_lut (.I0(GND_net), .I1(n2104), .I2(n1602), .I3(n50217), 
            .O(n8191[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1978_3_lut (.I0(n2831), .I1(n8347[19]), .I2(n294[4]), 
            .I3(GND_net), .O(n2942));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i39_2_lut (.I0(n2942), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4537));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1982_3_lut (.I0(n2835), .I1(n8347[15]), .I2(n294[4]), 
            .I3(GND_net), .O(n2946));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1983_3_lut (.I0(n2836), .I1(n8347[14]), .I2(n294[4]), 
            .I3(GND_net), .O(n2947));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i29_2_lut (.I0(n2947), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4538));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2793_8 (.CI(n50217), .I0(n2104), .I1(n1602), .CO(n50218));
    SB_LUT4 add_2793_7_lut (.I0(GND_net), .I1(n2105), .I2(n1459), .I3(n50216), 
            .O(n8191[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_7 (.CI(n50216), .I0(n2105), .I1(n1459), .CO(n50217));
    SB_LUT4 add_2793_6_lut (.I0(GND_net), .I1(n2106), .I2(n1460), .I3(n50215), 
            .O(n8191[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_6 (.CI(n50215), .I0(n2106), .I1(n1460), .CO(n50216));
    SB_LUT4 add_2793_5_lut (.I0(GND_net), .I1(n2107), .I2(n1011), .I3(n50214), 
            .O(n8191[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_5 (.CI(n50214), .I0(n2107), .I1(n1011), .CO(n50215));
    SB_LUT4 add_2793_4_lut (.I0(GND_net), .I1(n2108), .I2(n856), .I3(n50213), 
            .O(n8191[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut_adj_1019 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n60728));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1019.LUT_INIT = 16'hffef;
    SB_CARRY add_2793_4 (.CI(n50213), .I0(n2108), .I1(n856), .CO(n50214));
    SB_LUT4 i1_3_lut_4_lut_adj_1020 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n60760));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1020.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1997_i31_2_lut (.I0(n2946), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4539));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2793_3_lut (.I0(GND_net), .I1(n2109), .I2(n698), .I3(n50212), 
            .O(n8191[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_3 (.CI(n50212), .I0(n2109), .I1(n698), .CO(n50213));
    SB_LUT4 add_2793_2_lut (.I0(GND_net), .I1(n2110), .I2(n858), .I3(VCC_net), 
            .O(n8191[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2793_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2793_2 (.CI(VCC_net), .I0(n2110), .I1(n858), .CO(n50212));
    SB_LUT4 add_2792_14_lut (.I0(GND_net), .I1(n1966), .I2(n2272), .I3(n50211), 
            .O(n8165[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2792_13_lut (.I0(GND_net), .I1(n1967), .I2(n2144), .I3(n50210), 
            .O(n8165[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_13 (.CI(n50210), .I0(n1967), .I1(n2144), .CO(n50211));
    SB_LUT4 add_2792_12_lut (.I0(GND_net), .I1(n1968), .I2(n2013), .I3(n50209), 
            .O(n8165[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_12 (.CI(n50209), .I0(n1968), .I1(n2013), .CO(n50210));
    SB_LUT4 add_2792_11_lut (.I0(GND_net), .I1(n1969), .I2(n1879), .I3(n50208), 
            .O(n8165[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_11 (.CI(n50208), .I0(n1969), .I1(n1879), .CO(n50209));
    SB_LUT4 add_2792_10_lut (.I0(GND_net), .I1(n1970), .I2(n1742), .I3(n50207), 
            .O(n8165[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_10 (.CI(n50207), .I0(n1970), .I1(n1742), .CO(n50208));
    SB_LUT4 div_37_i1984_3_lut (.I0(n2837), .I1(n8347[13]), .I2(n294[4]), 
            .I3(GND_net), .O(n2948));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1985_3_lut (.I0(n2838), .I1(n8347[12]), .I2(n294[4]), 
            .I3(GND_net), .O(n2949));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1986_3_lut (.I0(n2839), .I1(n8347[11]), .I2(n294[4]), 
            .I3(GND_net), .O(n2950));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i23_2_lut (.I0(n2950), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4540));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2792_9_lut (.I0(GND_net), .I1(n1971), .I2(n1602), .I3(n50206), 
            .O(n8165[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_9 (.CI(n50206), .I0(n1971), .I1(n1602), .CO(n50207));
    SB_LUT4 add_2792_8_lut (.I0(GND_net), .I1(n1972), .I2(n1459), .I3(n50205), 
            .O(n8165[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR r_SM_Main_i1 (.Q(\r_SM_Main[1] ), .C(clk16MHz), .D(n3_adj_4541), 
            .R(\r_SM_Main[2] ));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2792_8 (.CI(n50205), .I0(n1972), .I1(n1459), .CO(n50206));
    SB_LUT4 add_2792_7_lut (.I0(GND_net), .I1(n1973), .I2(n1460), .I3(n50204), 
            .O(n8165[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i25_2_lut (.I0(n2949), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4542));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2792_7 (.CI(n50204), .I0(n1973), .I1(n1460), .CO(n50205));
    SB_LUT4 div_37_LessThan_1997_i27_2_lut (.I0(n2948), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4543));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2792_6_lut (.I0(GND_net), .I1(n1974), .I2(n1011), .I3(n50203), 
            .O(n8165[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1988_3_lut (.I0(n2841), .I1(n8347[9]), .I2(n294[4]), 
            .I3(GND_net), .O(n2952));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1987_3_lut (.I0(n2840), .I1(n8347[10]), .I2(n294[4]), 
            .I3(GND_net), .O(n2951));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1989_3_lut (.I0(n2842), .I1(n8347[8]), .I2(n294[4]), 
            .I3(GND_net), .O(n2953));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1981_3_lut (.I0(n2834), .I1(n8347[16]), .I2(n294[4]), 
            .I3(GND_net), .O(n2945));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1981_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2792_6 (.CI(n50203), .I0(n1974), .I1(n1011), .CO(n50204));
    SB_LUT4 add_2792_5_lut (.I0(GND_net), .I1(n1975), .I2(n856), .I3(n50202), 
            .O(n8165[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_5 (.CI(n50202), .I0(n1975), .I1(n856), .CO(n50203));
    SB_LUT4 add_2792_4_lut (.I0(GND_net), .I1(n1976), .I2(n698), .I3(n50201), 
            .O(n8165[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i17_2_lut (.I0(n2953), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4544));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2792_4 (.CI(n50201), .I0(n1976), .I1(n698), .CO(n50202));
    SB_LUT4 add_2792_3_lut (.I0(GND_net), .I1(n1977), .I2(n858), .I3(n50200), 
            .O(n8165[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i19_2_lut (.I0(n2952), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4545));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i19_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2792_3 (.CI(n50200), .I0(n1977), .I1(n858), .CO(n50201));
    SB_LUT4 add_2792_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n8165[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2792_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2792_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50200));
    SB_LUT4 add_2791_13_lut (.I0(GND_net), .I1(n1831), .I2(n2144), .I3(n50199), 
            .O(n8139[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2791_12_lut (.I0(GND_net), .I1(n1832), .I2(n2013), .I3(n50198), 
            .O(n8139[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52929_2_lut_4_lut (.I0(n67903), .I1(baudrate[10]), .I2(n1693), 
            .I3(n25639), .O(n294[13]));   // verilog/uart_rx.v(119[33:55])
    defparam i52929_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_CARRY add_2791_12 (.CI(n50198), .I0(n1832), .I1(n2013), .CO(n50199));
    SB_LUT4 add_2791_11_lut (.I0(GND_net), .I1(n1833), .I2(n1879), .I3(n50197), 
            .O(n8139[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_11 (.CI(n50197), .I0(n1833), .I1(n1879), .CO(n50198));
    SB_LUT4 add_2791_10_lut (.I0(GND_net), .I1(n1834), .I2(n1742), .I3(n50196), 
            .O(n8139[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_10 (.CI(n50196), .I0(n1834), .I1(n1742), .CO(n50197));
    SB_LUT4 add_2791_9_lut (.I0(GND_net), .I1(n1835), .I2(n1602), .I3(n50195), 
            .O(n8139[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_9 (.CI(n50195), .I0(n1835), .I1(n1602), .CO(n50196));
    SB_LUT4 add_2791_8_lut (.I0(GND_net), .I1(n1836), .I2(n1459), .I3(n50194), 
            .O(n8139[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i21_2_lut (.I0(n2951), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4546));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2791_8 (.CI(n50194), .I0(n1836), .I1(n1459), .CO(n50195));
    SB_LUT4 add_2791_7_lut (.I0(GND_net), .I1(n1837), .I2(n1460), .I3(n50193), 
            .O(n8139[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i33_2_lut (.I0(n2945), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4547));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1991_3_lut (.I0(n2844), .I1(n8347[6]), .I2(n294[4]), 
            .I3(GND_net), .O(n2955));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1992_3_lut (.I0(n2845), .I1(n8347[5]), .I2(n294[4]), 
            .I3(GND_net), .O(n2956));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i13_2_lut (.I0(n2955), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4548));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2791_7 (.CI(n50193), .I0(n1837), .I1(n1460), .CO(n50194));
    SB_LUT4 add_2791_6_lut (.I0(GND_net), .I1(n1838), .I2(n1011), .I3(n50192), 
            .O(n8139[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_6 (.CI(n50192), .I0(n1838), .I1(n1011), .CO(n50193));
    SB_LUT4 add_2791_5_lut (.I0(GND_net), .I1(n1839), .I2(n856), .I3(n50191), 
            .O(n8139[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_5 (.CI(n50191), .I0(n1839), .I1(n856), .CO(n50192));
    SB_LUT4 add_2791_4_lut (.I0(GND_net), .I1(n1840), .I2(n698), .I3(n50190), 
            .O(n8139[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_4 (.CI(n50190), .I0(n1840), .I1(n698), .CO(n50191));
    SB_LUT4 add_2791_3_lut (.I0(GND_net), .I1(n1841), .I2(n858), .I3(n50189), 
            .O(n8139[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2791_3 (.CI(n50189), .I0(n1841), .I1(n858), .CO(n50190));
    SB_LUT4 add_2791_2_lut (.I0(n58103), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60318)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2791_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2791_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50189));
    SB_LUT4 add_2790_11_lut (.I0(GND_net), .I1(n1693), .I2(n2013), .I3(n50188), 
            .O(n8113[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2790_10_lut (.I0(GND_net), .I1(n1694), .I2(n1879), .I3(n50187), 
            .O(n8113[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_10 (.CI(n50187), .I0(n1694), .I1(n1879), .CO(n50188));
    SB_LUT4 add_2790_9_lut (.I0(GND_net), .I1(n1695), .I2(n1742), .I3(n50186), 
            .O(n8113[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_9 (.CI(n50186), .I0(n1695), .I1(n1742), .CO(n50187));
    SB_LUT4 add_2790_8_lut (.I0(GND_net), .I1(n1696), .I2(n1602), .I3(n50185), 
            .O(n8113[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_8 (.CI(n50185), .I0(n1696), .I1(n1602), .CO(n50186));
    SB_LUT4 add_2790_7_lut (.I0(GND_net), .I1(n1697), .I2(n1459), .I3(n50184), 
            .O(n8113[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_7 (.CI(n50184), .I0(n1697), .I1(n1459), .CO(n50185));
    SB_LUT4 add_2790_6_lut (.I0(GND_net), .I1(n1698), .I2(n1460), .I3(n50183), 
            .O(n8113[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_6 (.CI(n50183), .I0(n1698), .I1(n1460), .CO(n50184));
    SB_LUT4 add_2790_5_lut (.I0(GND_net), .I1(n1699), .I2(n1011), .I3(n50182), 
            .O(n8113[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_5 (.CI(n50182), .I0(n1699), .I1(n1011), .CO(n50183));
    SB_LUT4 div_37_LessThan_1997_i15_2_lut (.I0(n2954), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4549));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50106_4_lut (.I0(n33_adj_4547), .I1(n21_adj_4546), .I2(n19_adj_4545), 
            .I3(n17_adj_4544), .O(n65792));
    defparam i50106_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2790_4_lut (.I0(GND_net), .I1(n1700), .I2(n856), .I3(n50181), 
            .O(n8113[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_4 (.CI(n50181), .I0(n1700), .I1(n856), .CO(n50182));
    SB_LUT4 add_2790_3_lut (.I0(GND_net), .I1(n1701), .I2(n698), .I3(n50180), 
            .O(n8113[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_3 (.CI(n50180), .I0(n1701), .I1(n698), .CO(n50181));
    SB_LUT4 add_2790_2_lut (.I0(GND_net), .I1(n1702), .I2(n858), .I3(VCC_net), 
            .O(n8113[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2790_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2790_2 (.CI(VCC_net), .I0(n1702), .I1(n858), .CO(n50180));
    SB_LUT4 add_2789_11_lut (.I0(GND_net), .I1(n1552), .I2(n1879), .I3(n50179), 
            .O(n8087[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51017_4_lut (.I0(n15_adj_4549), .I1(n13_adj_4548), .I2(n2956), 
            .I3(baudrate[2]), .O(n66703));
    defparam i51017_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i51651_4_lut (.I0(n21_adj_4546), .I1(n19_adj_4545), .I2(n17_adj_4544), 
            .I3(n66703), .O(n67337));
    defparam i51651_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 add_2789_10_lut (.I0(GND_net), .I1(n1553), .I2(n1742), .I3(n50178), 
            .O(n8087[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_10 (.CI(n50178), .I0(n1553), .I1(n1742), .CO(n50179));
    SB_LUT4 add_2789_9_lut (.I0(GND_net), .I1(n1554), .I2(n1602), .I3(n50177), 
            .O(n8087[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_9 (.CI(n50177), .I0(n1554), .I1(n1602), .CO(n50178));
    SB_LUT4 add_2789_8_lut (.I0(GND_net), .I1(n1555), .I2(n1459), .I3(n50176), 
            .O(n8087[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_8 (.CI(n50176), .I0(n1555), .I1(n1459), .CO(n50177));
    SB_LUT4 add_2789_7_lut (.I0(GND_net), .I1(n1556), .I2(n1460), .I3(n50175), 
            .O(n8087[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_7 (.CI(n50175), .I0(n1556), .I1(n1460), .CO(n50176));
    SB_LUT4 add_2789_6_lut (.I0(GND_net), .I1(n1557), .I2(n1011), .I3(n50174), 
            .O(n8087[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_6 (.CI(n50174), .I0(n1557), .I1(n1011), .CO(n50175));
    SB_LUT4 add_2789_5_lut (.I0(GND_net), .I1(n1558), .I2(n856), .I3(n50173), 
            .O(n8087[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_5 (.CI(n50173), .I0(n1558), .I1(n856), .CO(n50174));
    SB_LUT4 add_2789_4_lut (.I0(GND_net), .I1(n1559), .I2(n698), .I3(n50172), 
            .O(n8087[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_4 (.CI(n50172), .I0(n1559), .I1(n698), .CO(n50173));
    SB_LUT4 add_2789_3_lut (.I0(GND_net), .I1(n1560), .I2(n858), .I3(n50171), 
            .O(n8087[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_3 (.CI(n50171), .I0(n1560), .I1(n858), .CO(n50172));
    SB_LUT4 add_2789_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n8087[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2789_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2789_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50171));
    SB_LUT4 add_2788_10_lut (.I0(GND_net), .I1(n1408), .I2(n1742), .I3(n50170), 
            .O(n8061[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2788_9_lut (.I0(GND_net), .I1(n1409), .I2(n1602), .I3(n50169), 
            .O(n8061[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_9 (.CI(n50169), .I0(n1409), .I1(n1602), .CO(n50170));
    SB_LUT4 add_2788_8_lut (.I0(GND_net), .I1(n1410), .I2(n1459), .I3(n50168), 
            .O(n8061[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_8 (.CI(n50168), .I0(n1410), .I1(n1459), .CO(n50169));
    SB_LUT4 add_2788_7_lut (.I0(GND_net), .I1(n1411), .I2(n1460), .I3(n50167), 
            .O(n8061[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_7 (.CI(n50167), .I0(n1411), .I1(n1460), .CO(n50168));
    SB_LUT4 add_2788_6_lut (.I0(GND_net), .I1(n1412), .I2(n1011), .I3(n50166), 
            .O(n8061[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_6 (.CI(n50166), .I0(n1412), .I1(n1011), .CO(n50167));
    SB_LUT4 add_2788_5_lut (.I0(GND_net), .I1(n1413), .I2(n856), .I3(n50165), 
            .O(n8061[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_5 (.CI(n50165), .I0(n1413), .I1(n856), .CO(n50166));
    SB_LUT4 add_2788_4_lut (.I0(GND_net), .I1(n1414), .I2(n698), .I3(n50164), 
            .O(n8061[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2788_4 (.CI(n50164), .I0(n1414), .I1(n698), .CO(n50165));
    SB_LUT4 add_2788_3_lut (.I0(GND_net), .I1(n1415), .I2(n858), .I3(n50163), 
            .O(n8061[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i51649_4_lut (.I0(n27_adj_4543), .I1(n25_adj_4542), .I2(n23_adj_4540), 
            .I3(n67337), .O(n67335));
    defparam i51649_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY add_2788_3 (.CI(n50163), .I0(n1415), .I1(n858), .CO(n50164));
    SB_LUT4 add_2788_2_lut (.I0(n58112), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60316)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2788_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2788_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50163));
    SB_LUT4 add_2787_9_lut (.I0(GND_net), .I1(n1261), .I2(n1602), .I3(n50162), 
            .O(n8035[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2787_8_lut (.I0(GND_net), .I1(n1262), .I2(n1459), .I3(n50161), 
            .O(n8035[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_8 (.CI(n50161), .I0(n1262), .I1(n1459), .CO(n50162));
    SB_LUT4 add_2787_7_lut (.I0(GND_net), .I1(n1263), .I2(n1460), .I3(n50160), 
            .O(n8035[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_7 (.CI(n50160), .I0(n1263), .I1(n1460), .CO(n50161));
    SB_LUT4 add_2787_6_lut (.I0(GND_net), .I1(n1264), .I2(n1011), .I3(n50159), 
            .O(n8035[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_6 (.CI(n50159), .I0(n1264), .I1(n1011), .CO(n50160));
    SB_LUT4 add_2787_5_lut (.I0(GND_net), .I1(n1265), .I2(n856), .I3(n50158), 
            .O(n8035[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_5 (.CI(n50158), .I0(n1265), .I1(n856), .CO(n50159));
    SB_LUT4 i50108_4_lut (.I0(n33_adj_4547), .I1(n31_adj_4539), .I2(n29_adj_4538), 
            .I3(n67335), .O(n65794));
    defparam i50108_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2787_4_lut (.I0(GND_net), .I1(n1266), .I2(n698), .I3(n50157), 
            .O(n8035[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_4 (.CI(n50157), .I0(n1266), .I1(n698), .CO(n50158));
    SB_LUT4 add_2787_3_lut (.I0(GND_net), .I1(n1267), .I2(n858), .I3(n50156), 
            .O(n8035[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2787_3 (.CI(n50156), .I0(n1267), .I1(n858), .CO(n50157));
    SB_LUT4 add_2787_2_lut (.I0(n58116), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60314)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2787_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2787_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50156));
    SB_LUT4 add_2786_8_lut (.I0(GND_net), .I1(n1111), .I2(n1459), .I3(n50155), 
            .O(n8009[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2786_7_lut (.I0(GND_net), .I1(n1112), .I2(n1460), .I3(n50154), 
            .O(n8009[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_7 (.CI(n50154), .I0(n1112), .I1(n1460), .CO(n50155));
    SB_LUT4 add_2786_6_lut (.I0(GND_net), .I1(n1113), .I2(n1011), .I3(n50153), 
            .O(n8009[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2786_6 (.CI(n50153), .I0(n1113), .I1(n1011), .CO(n50154));
    SB_LUT4 add_2786_5_lut (.I0(GND_net), .I1(n1114), .I2(n856), .I3(n50152), 
            .O(n8009[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i10_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2957), .I3(GND_net), .O(n10_adj_4550));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2786_5 (.CI(n50152), .I0(n1114), .I1(n856), .CO(n50153));
    SB_LUT4 add_2786_4_lut (.I0(GND_net), .I1(n1115), .I2(n698), .I3(n50151), 
            .O(n8009[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i52145_3_lut (.I0(n10_adj_4550), .I1(baudrate[13]), .I2(n33_adj_4547), 
            .I3(GND_net), .O(n67831));   // verilog/uart_rx.v(119[33:55])
    defparam i52145_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2786_4 (.CI(n50151), .I0(n1115), .I1(n698), .CO(n50152));
    SB_LUT4 i52146_3_lut (.I0(n67831), .I1(baudrate[14]), .I2(n35_adj_4536), 
            .I3(GND_net), .O(n67832));   // verilog/uart_rx.v(119[33:55])
    defparam i52146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2786_3_lut (.I0(GND_net), .I1(n1116), .I2(n858), .I3(n50150), 
            .O(n8009[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1997_i36_3_lut (.I0(n18), .I1(baudrate[17]), 
            .I2(n41_adj_4535), .I3(GND_net), .O(n36_adj_4551));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i36_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2786_3 (.CI(n50150), .I0(n1116), .I1(n858), .CO(n50151));
    SB_LUT4 add_2786_2_lut (.I0(n58120), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n60312)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2786_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2786_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n50150));
    SB_LUT4 i50102_4_lut (.I0(n39_adj_4537), .I1(n37_adj_4534), .I2(n35_adj_4536), 
            .I3(n65792), .O(n65788));
    defparam i50102_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52477_4_lut (.I0(n36_adj_4551), .I1(n16_adj_4552), .I2(n41_adj_4535), 
            .I3(n65786), .O(n68163));   // verilog/uart_rx.v(119[33:55])
    defparam i52477_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52046_3_lut (.I0(n67832), .I1(baudrate[15]), .I2(n37_adj_4534), 
            .I3(GND_net), .O(n67732));   // verilog/uart_rx.v(119[33:55])
    defparam i52046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i22_3_lut (.I0(n14_adj_4553), .I1(baudrate[9]), 
            .I2(n25_adj_4542), .I3(GND_net), .O(n22));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53406_2_lut_4_lut (.I0(n68060), .I1(baudrate[6]), .I2(n1111), 
            .I3(n62572), .O(n294[17]));   // verilog/uart_rx.v(119[33:55])
    defparam i53406_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_1021 (.I0(baudrate[30]), .I1(baudrate[25]), 
            .I2(baudrate[31]), .I3(baudrate[26]), .O(n61766));
    defparam i1_2_lut_4_lut_adj_1021.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1022 (.I0(n68060), .I1(baudrate[6]), .I2(n1111), 
            .I3(n60312), .O(n1267));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1022.LUT_INIT = 16'h7100;
    SB_LUT4 i52475_4_lut (.I0(n22), .I1(n12_adj_4554), .I2(n25_adj_4542), 
            .I3(n65800), .O(n68161));   // verilog/uart_rx.v(119[33:55])
    defparam i52475_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52476_3_lut (.I0(n68161), .I1(baudrate[10]), .I2(n27_adj_4543), 
            .I3(GND_net), .O(n68162));   // verilog/uart_rx.v(119[33:55])
    defparam i52476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52360_3_lut (.I0(n68162), .I1(baudrate[11]), .I2(n29_adj_4538), 
            .I3(GND_net), .O(n68046));   // verilog/uart_rx.v(119[33:55])
    defparam i52360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_765_i40_3_lut_3_lut (.I0(n1114), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n40_adj_4460));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i40_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i51960_4_lut (.I0(n39_adj_4537), .I1(n37_adj_4534), .I2(n35_adj_4536), 
            .I3(n65794), .O(n67646));
    defparam i51960_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52603_4_lut (.I0(n67732), .I1(n68163), .I2(n41_adj_4535), 
            .I3(n65788), .O(n68289));   // verilog/uart_rx.v(119[33:55])
    defparam i52603_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52304_3_lut (.I0(n68046), .I1(baudrate[12]), .I2(n31_adj_4539), 
            .I3(GND_net), .O(n67990));   // verilog/uart_rx.v(119[33:55])
    defparam i52304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52627_4_lut (.I0(n67990), .I1(n68289), .I2(n41_adj_4535), 
            .I3(n67646), .O(n68313));   // verilog/uart_rx.v(119[33:55])
    defparam i52627_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52628_3_lut (.I0(n68313), .I1(baudrate[18]), .I2(n2940), 
            .I3(GND_net), .O(n68314));   // verilog/uart_rx.v(119[33:55])
    defparam i52628_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52624_3_lut (.I0(n68314), .I1(baudrate[19]), .I2(n2939), 
            .I3(GND_net), .O(n68310));   // verilog/uart_rx.v(119[33:55])
    defparam i52624_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50473_3_lut_4_lut (.I0(n1114), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1115), .O(n66159));   // verilog/uart_rx.v(119[33:55])
    defparam i50473_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1250_i30_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1839), .I3(GND_net), .O(n30_adj_4555));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50408_2_lut_4_lut (.I0(n1834), .I1(baudrate[8]), .I2(n1838), 
            .I3(baudrate[4]), .O(n66094));
    defparam i50408_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_3_lut_4_lut_adj_1023 (.I0(baudrate[3]), .I1(n42), .I2(baudrate[4]), 
            .I3(n20931), .O(n58551));   // verilog/uart_rx.v(119[33:55])
    defparam i1_3_lut_4_lut_adj_1023.LUT_INIT = 16'hff4f;
    SB_LUT4 div_37_i1899_3_lut (.I0(n2713), .I1(n8321[23]), .I2(n294[5]), 
            .I3(GND_net), .O(n2827));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1900_3_lut (.I0(n2714), .I1(n8321[22]), .I2(n294[5]), 
            .I3(GND_net), .O(n2828));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5756_2_lut_3_lut (.I0(baudrate[3]), .I1(n42), .I2(n20931), 
            .I3(GND_net), .O(n44));   // verilog/uart_rx.v(119[33:55])
    defparam i5756_2_lut_3_lut.LUT_INIT = 16'hf4f4;
    SB_LUT4 div_37_i1905_3_lut (.I0(n2719), .I1(n8321[17]), .I2(n294[5]), 
            .I3(GND_net), .O(n2833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1901_3_lut (.I0(n2715), .I1(n8321[21]), .I2(n294[5]), 
            .I3(GND_net), .O(n2829));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i43_2_lut (.I0(n2829), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4556));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1903_3_lut (.I0(n2717), .I1(n8321[19]), .I2(n294[5]), 
            .I3(GND_net), .O(n2831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i32_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1834), .I3(GND_net), .O(n32_adj_4557));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i32_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1904_3_lut (.I0(n2718), .I1(n8321[18]), .I2(n294[5]), 
            .I3(GND_net), .O(n2832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i37_2_lut (.I0(n2832), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4558));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i39_2_lut (.I0(n2831), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4559));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1902_3_lut (.I0(n2716), .I1(n8321[20]), .I2(n294[5]), 
            .I3(GND_net), .O(n2830));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i41_2_lut (.I0(n2830), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4560));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1906_3_lut (.I0(n2720), .I1(n8321[16]), .I2(n294[5]), 
            .I3(GND_net), .O(n2834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53411_2_lut_4_lut (.I0(n67909), .I1(baudrate[7]), .I2(n1261), 
            .I3(n62570), .O(n294[16]));   // verilog/uart_rx.v(119[33:55])
    defparam i53411_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_1024 (.I0(n67909), .I1(baudrate[7]), .I2(n1261), 
            .I3(n60314), .O(n1415));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1024.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_i1907_3_lut (.I0(n2721), .I1(n8321[15]), .I2(n294[5]), 
            .I3(GND_net), .O(n2835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i31_2_lut (.I0(n2835), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4561));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i33_2_lut (.I0(n2834), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4562));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1908_3_lut (.I0(n2722), .I1(n8321[14]), .I2(n294[5]), 
            .I3(GND_net), .O(n2836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1910_3_lut (.I0(n2724), .I1(n8321[12]), .I2(n294[5]), 
            .I3(GND_net), .O(n2838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1909_3_lut (.I0(n2723), .I1(n8321[13]), .I2(n294[5]), 
            .I3(GND_net), .O(n2837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i25_2_lut (.I0(n2838), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4563));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i27_2_lut (.I0(n2837), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4564));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i29_2_lut (.I0(n2836), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4565));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1914_3_lut (.I0(n2728), .I1(n8321[8]), .I2(n294[5]), 
            .I3(GND_net), .O(n2842));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1915_3_lut (.I0(n2729), .I1(n8321[7]), .I2(n294[5]), 
            .I3(GND_net), .O(n2843));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1916_3_lut (.I0(n2730), .I1(n8321[6]), .I2(n294[5]), 
            .I3(GND_net), .O(n2844));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i15_2_lut (.I0(n2843), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4566));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i17_2_lut (.I0(n2842), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4567));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1912_3_lut (.I0(n2726), .I1(n8321[10]), .I2(n294[5]), 
            .I3(GND_net), .O(n2840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1911_3_lut (.I0(n2725), .I1(n8321[11]), .I2(n294[5]), 
            .I3(GND_net), .O(n2839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1913_3_lut (.I0(n2727), .I1(n8321[9]), .I2(n294[5]), 
            .I3(GND_net), .O(n2841));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i19_2_lut (.I0(n2841), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4568));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i21_2_lut (.I0(n2840), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4569));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i23_2_lut (.I0(n2839), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4570));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_866_i38_3_lut_3_lut (.I0(n1265), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n38_adj_4456));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i38_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i46896_1_lut (.I0(n62572), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n58120));
    defparam i46896_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i46892_1_lut (.I0(n62568), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n58112));
    defparam i46892_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1922_i35_2_lut (.I0(n2833), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4571));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46870_1_lut (.I0(n62546), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n58103));
    defparam i46870_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i50163_4_lut (.I0(n35_adj_4571), .I1(n23_adj_4570), .I2(n21_adj_4569), 
            .I3(n19_adj_4568), .O(n65849));
    defparam i50163_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51077_4_lut (.I0(n17_adj_4567), .I1(n15_adj_4566), .I2(n2844), 
            .I3(baudrate[2]), .O(n66763));
    defparam i51077_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i51675_4_lut (.I0(n23_adj_4570), .I1(n21_adj_4569), .I2(n19_adj_4568), 
            .I3(n66763), .O(n67361));
    defparam i51675_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51671_4_lut (.I0(n29_adj_4565), .I1(n27_adj_4564), .I2(n25_adj_4563), 
            .I3(n67361), .O(n67357));
    defparam i51671_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50167_4_lut (.I0(n35_adj_4571), .I1(n33_adj_4562), .I2(n31_adj_4561), 
            .I3(n67357), .O(n65853));
    defparam i50167_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1922_i12_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2845), .I3(GND_net), .O(n12_adj_4572));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52151_3_lut (.I0(n12_adj_4572), .I1(baudrate[13]), .I2(n35_adj_4571), 
            .I3(GND_net), .O(n67837));   // verilog/uart_rx.v(119[33:55])
    defparam i52151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i38_3_lut (.I0(n20_adj_4573), .I1(baudrate[17]), 
            .I2(n43_adj_4556), .I3(GND_net), .O(n38_adj_4574));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52152_3_lut (.I0(n67837), .I1(baudrate[14]), .I2(n37_adj_4558), 
            .I3(GND_net), .O(n67838));   // verilog/uart_rx.v(119[33:55])
    defparam i52152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50155_4_lut (.I0(n41_adj_4560), .I1(n39_adj_4559), .I2(n37_adj_4558), 
            .I3(n65849), .O(n65841));
    defparam i50155_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52149_4_lut (.I0(n38_adj_4574), .I1(n18_adj_4575), .I2(n43_adj_4556), 
            .I3(n65834), .O(n67835));   // verilog/uart_rx.v(119[33:55])
    defparam i52149_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52038_3_lut (.I0(n67838), .I1(baudrate[15]), .I2(n39_adj_4559), 
            .I3(GND_net), .O(n67724));   // verilog/uart_rx.v(119[33:55])
    defparam i52038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i24_3_lut (.I0(n16_adj_4576), .I1(baudrate[9]), 
            .I2(n27_adj_4564), .I3(GND_net), .O(n24_adj_4577));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52473_4_lut (.I0(n24_adj_4577), .I1(n14_adj_4578), .I2(n27_adj_4564), 
            .I3(n65861), .O(n68159));   // verilog/uart_rx.v(119[33:55])
    defparam i52473_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52474_3_lut (.I0(n68159), .I1(baudrate[10]), .I2(n29_adj_4565), 
            .I3(GND_net), .O(n68160));   // verilog/uart_rx.v(119[33:55])
    defparam i52474_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52362_3_lut (.I0(n68160), .I1(baudrate[11]), .I2(n31_adj_4561), 
            .I3(GND_net), .O(n68048));   // verilog/uart_rx.v(119[33:55])
    defparam i52362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51988_4_lut (.I0(n41_adj_4560), .I1(n39_adj_4559), .I2(n37_adj_4558), 
            .I3(n65853), .O(n67674));
    defparam i51988_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52464_4_lut (.I0(n67724), .I1(n67835), .I2(n43_adj_4556), 
            .I3(n65841), .O(n68150));   // verilog/uart_rx.v(119[33:55])
    defparam i52464_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52302_3_lut (.I0(n68048), .I1(baudrate[12]), .I2(n33_adj_4562), 
            .I3(GND_net), .O(n67988));   // verilog/uart_rx.v(119[33:55])
    defparam i52302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52611_4_lut (.I0(n67988), .I1(n68150), .I2(n43_adj_4556), 
            .I3(n67674), .O(n68297));   // verilog/uart_rx.v(119[33:55])
    defparam i52611_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52612_3_lut (.I0(n68297), .I1(baudrate[18]), .I2(n2828), 
            .I3(GND_net), .O(n68298));   // verilog/uart_rx.v(119[33:55])
    defparam i52612_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50513_4_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n4937), .I3(\o_Rx_DV_N_3488[8] ), .O(n65381));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i50513_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i50599_4_lut (.I0(r_Rx_Data), .I1(\o_Rx_DV_N_3488[12] ), .I2(n56722), 
            .I3(r_SM_Main[0]), .O(n65387));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i50599_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i50510_4_lut (.I0(n65381), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n65378));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i50510_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50516_4_lut (.I0(n65387), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n65384));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i50516_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_1_i3_4_lut (.I0(n65384), .I1(n65378), 
            .I2(\r_SM_Main[1] ), .I3(n27), .O(n3_adj_4541));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_1_i3_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 i50465_3_lut_4_lut (.I0(n1265), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1266), .O(n66151));   // verilog/uart_rx.v(119[33:55])
    defparam i50465_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i53414_2_lut_4_lut (.I0(n67696), .I1(baudrate[8]), .I2(n1408), 
            .I3(n62568), .O(n294[15]));   // verilog/uart_rx.v(119[33:55])
    defparam i53414_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1822_3_lut (.I0(n2596), .I1(n8295[23]), .I2(n294[6]), 
            .I3(GND_net), .O(n2713));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1827_3_lut (.I0(n2601), .I1(n8295[18]), .I2(n294[6]), 
            .I3(GND_net), .O(n2718));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1823_3_lut (.I0(n2597), .I1(n8295[22]), .I2(n294[6]), 
            .I3(GND_net), .O(n2714));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i45_2_lut (.I0(n2714), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4579));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1826_3_lut (.I0(n2600), .I1(n8295[19]), .I2(n294[6]), 
            .I3(GND_net), .O(n2717));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1025 (.I0(n67696), .I1(baudrate[8]), .I2(n1408), 
            .I3(n60316), .O(n1560));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1025.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_i1825_3_lut (.I0(n2599), .I1(n8295[20]), .I2(n294[6]), 
            .I3(GND_net), .O(n2716));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i39_2_lut (.I0(n2717), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4580));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i41_2_lut (.I0(n2716), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4581));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1828_3_lut (.I0(n2602), .I1(n8295[17]), .I2(n294[6]), 
            .I3(GND_net), .O(n2719));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1829_3_lut (.I0(n2603), .I1(n8295[16]), .I2(n294[6]), 
            .I3(GND_net), .O(n2720));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i33_2_lut (.I0(n2720), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4582));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i35_2_lut (.I0(n2719), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4583));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1830_3_lut (.I0(n2604), .I1(n8295[15]), .I2(n294[6]), 
            .I3(GND_net), .O(n2721));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1831_3_lut (.I0(n2605), .I1(n8295[14]), .I2(n294[6]), 
            .I3(GND_net), .O(n2722));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1832_3_lut (.I0(n2606), .I1(n8295[13]), .I2(n294[6]), 
            .I3(GND_net), .O(n2723));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i27_2_lut (.I0(n2723), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4584));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i29_2_lut (.I0(n2722), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4585));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i31_2_lut (.I0(n2721), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4586));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1824_3_lut (.I0(n2598), .I1(n8295[21]), .I2(n294[6]), 
            .I3(GND_net), .O(n2715));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i43_2_lut (.I0(n2715), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4587));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1837_3_lut (.I0(n2611), .I1(n8295[8]), .I2(n294[6]), 
            .I3(GND_net), .O(n2728));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1836_3_lut (.I0(n2610), .I1(n8295[9]), .I2(n294[6]), 
            .I3(GND_net), .O(n2727));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1838_3_lut (.I0(n2612), .I1(n8295[7]), .I2(n294[6]), 
            .I3(GND_net), .O(n2729));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i17_2_lut (.I0(n2728), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4588));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i19_2_lut (.I0(n2727), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4589));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1833_3_lut (.I0(n2607), .I1(n8295[12]), .I2(n294[6]), 
            .I3(GND_net), .O(n2724));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1834_3_lut (.I0(n2608), .I1(n8295[11]), .I2(n294[6]), 
            .I3(GND_net), .O(n2725));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1835_3_lut (.I0(n2609), .I1(n8295[10]), .I2(n294[6]), 
            .I3(GND_net), .O(n2726));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i21_2_lut (.I0(n2726), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4590));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i23_2_lut (.I0(n2725), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4591));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i25_2_lut (.I0(n2724), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4592));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i28_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1975), .I3(GND_net), .O(n28));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50394_2_lut_4_lut (.I0(n1970), .I1(baudrate[8]), .I2(n1974), 
            .I3(baudrate[4]), .O(n66080));
    defparam i50394_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1845_i37_2_lut (.I0(n2718), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4593));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50203_4_lut (.I0(n37_adj_4593), .I1(n25_adj_4592), .I2(n23_adj_4591), 
            .I3(n21_adj_4590), .O(n65889));
    defparam i50203_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51163_4_lut (.I0(n19_adj_4589), .I1(n17_adj_4588), .I2(n2729), 
            .I3(baudrate[2]), .O(n66849));
    defparam i51163_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i51709_4_lut (.I0(n25_adj_4592), .I1(n23_adj_4591), .I2(n21_adj_4590), 
            .I3(n66849), .O(n67395));
    defparam i51709_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i51695_4_lut (.I0(n31_adj_4586), .I1(n29_adj_4585), .I2(n27_adj_4584), 
            .I3(n67395), .O(n67381));
    defparam i51695_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i50207_4_lut (.I0(n37_adj_4593), .I1(n35_adj_4583), .I2(n33_adj_4582), 
            .I3(n67381), .O(n65893));
    defparam i50207_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1845_i14_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2730), .I3(GND_net), .O(n14_adj_4594));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i14_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52157_3_lut (.I0(n14_adj_4594), .I1(baudrate[13]), .I2(n37_adj_4593), 
            .I3(GND_net), .O(n67843));   // verilog/uart_rx.v(119[33:55])
    defparam i52157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52158_3_lut (.I0(n67843), .I1(baudrate[14]), .I2(n39_adj_4580), 
            .I3(GND_net), .O(n67844));   // verilog/uart_rx.v(119[33:55])
    defparam i52158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i40_3_lut (.I0(n22_adj_4595), .I1(baudrate[17]), 
            .I2(n45_adj_4579), .I3(GND_net), .O(n40_adj_4596));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50196_4_lut (.I0(n43_adj_4587), .I1(n41_adj_4581), .I2(n39_adj_4580), 
            .I3(n65889), .O(n65882));
    defparam i50196_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51699_4_lut (.I0(n40_adj_4596), .I1(n20_adj_4597), .I2(n45_adj_4579), 
            .I3(n65880), .O(n67385));   // verilog/uart_rx.v(119[33:55])
    defparam i51699_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52034_3_lut (.I0(n67844), .I1(baudrate[15]), .I2(n41_adj_4581), 
            .I3(GND_net), .O(n67720));   // verilog/uart_rx.v(119[33:55])
    defparam i52034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i26_3_lut (.I0(n18_adj_4598), .I1(baudrate[9]), 
            .I2(n29_adj_4585), .I3(GND_net), .O(n26_adj_4599));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52471_4_lut (.I0(n26_adj_4599), .I1(n16_adj_4600), .I2(n29_adj_4585), 
            .I3(n65902), .O(n68157));   // verilog/uart_rx.v(119[33:55])
    defparam i52471_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52472_3_lut (.I0(n68157), .I1(baudrate[10]), .I2(n31_adj_4586), 
            .I3(GND_net), .O(n68158));   // verilog/uart_rx.v(119[33:55])
    defparam i52472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52364_3_lut (.I0(n68158), .I1(baudrate[11]), .I2(n33_adj_4582), 
            .I3(GND_net), .O(n68050));   // verilog/uart_rx.v(119[33:55])
    defparam i52364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52014_4_lut (.I0(n43_adj_4587), .I1(n41_adj_4581), .I2(n39_adj_4580), 
            .I3(n65893), .O(n67700));
    defparam i52014_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52298_4_lut (.I0(n67720), .I1(n67385), .I2(n45_adj_4579), 
            .I3(n65882), .O(n67984));   // verilog/uart_rx.v(119[33:55])
    defparam i52298_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_LessThan_1341_i30_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1970), .I3(GND_net), .O(n30_adj_4601));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52297_3_lut (.I0(n68050), .I1(baudrate[12]), .I2(n35_adj_4583), 
            .I3(GND_net), .O(n67983));   // verilog/uart_rx.v(119[33:55])
    defparam i52297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52300_4_lut (.I0(n67983), .I1(n67984), .I2(n45_adj_4579), 
            .I3(n67700), .O(n67986));   // verilog/uart_rx.v(119[33:55])
    defparam i52300_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1743_3_lut (.I0(n2476), .I1(n8269[23]), .I2(n294[7]), 
            .I3(GND_net), .O(n2596));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1744_3_lut (.I0(n2477), .I1(n8269[22]), .I2(n294[7]), 
            .I3(GND_net), .O(n2597));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1748_3_lut (.I0(n2481), .I1(n8269[18]), .I2(n294[7]), 
            .I3(GND_net), .O(n2601));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i37_2_lut (.I0(n2601), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1745_3_lut (.I0(n2478), .I1(n8269[21]), .I2(n294[7]), 
            .I3(GND_net), .O(n2598));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i43_2_lut (.I0(n2598), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4603));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1746_3_lut (.I0(n2479), .I1(n8269[20]), .I2(n294[7]), 
            .I3(GND_net), .O(n2599));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1747_3_lut (.I0(n2480), .I1(n8269[19]), .I2(n294[7]), 
            .I3(GND_net), .O(n2600));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i39_2_lut (.I0(n2600), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4604));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i41_2_lut (.I0(n2599), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4605));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1749_3_lut (.I0(n2482), .I1(n8269[17]), .I2(n294[7]), 
            .I3(GND_net), .O(n2602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1751_3_lut (.I0(n2484), .I1(n8269[15]), .I2(n294[7]), 
            .I3(GND_net), .O(n2604));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1750_3_lut (.I0(n2483), .I1(n8269[16]), .I2(n294[7]), 
            .I3(GND_net), .O(n2603));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i31_2_lut (.I0(n2604), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4606));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i33_2_lut (.I0(n2603), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4607));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i35_2_lut (.I0(n2602), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4608));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1752_3_lut (.I0(n2485), .I1(n8269[14]), .I2(n294[7]), 
            .I3(GND_net), .O(n2605));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1753_3_lut (.I0(n2486), .I1(n8269[13]), .I2(n294[7]), 
            .I3(GND_net), .O(n2606));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i27_2_lut (.I0(n2606), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4609));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i29_2_lut (.I0(n2605), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4610));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1757_3_lut (.I0(n2490), .I1(n8269[9]), .I2(n294[7]), 
            .I3(GND_net), .O(n2610));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1756_3_lut (.I0(n2489), .I1(n8269[10]), .I2(n294[7]), 
            .I3(GND_net), .O(n2609));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i19_2_lut (.I0(n2610), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4611));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i21_2_lut (.I0(n2609), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4612));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1755_3_lut (.I0(n2488), .I1(n8269[11]), .I2(n294[7]), 
            .I3(GND_net), .O(n2608));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1754_3_lut (.I0(n2487), .I1(n8269[12]), .I2(n294[7]), 
            .I3(GND_net), .O(n2607));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i23_2_lut (.I0(n2608), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4613));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i25_2_lut (.I0(n2607), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4614));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1758_3_lut (.I0(n2491), .I1(n8269[8]), .I2(n294[7]), 
            .I3(GND_net), .O(n2611));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i17_2_lut (.I0(n2611), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4615));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50261_4_lut (.I0(n23_adj_4613), .I1(n21_adj_4612), .I2(n19_adj_4611), 
            .I3(n17_adj_4615), .O(n65947));
    defparam i50261_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50255_4_lut (.I0(n29_adj_4610), .I1(n27_adj_4609), .I2(n25_adj_4614), 
            .I3(n65947), .O(n65941));
    defparam i50255_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52081_4_lut (.I0(n35_adj_4608), .I1(n33_adj_4607), .I2(n31_adj_4606), 
            .I3(n65941), .O(n67767));
    defparam i52081_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i16_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2612), .I3(GND_net), .O(n16_adj_4616));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51874_3_lut (.I0(n16_adj_4616), .I1(baudrate[13]), .I2(n39_adj_4604), 
            .I3(GND_net), .O(n67560));   // verilog/uart_rx.v(119[33:55])
    defparam i51874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51875_3_lut (.I0(n67560), .I1(baudrate[14]), .I2(n41_adj_4605), 
            .I3(GND_net), .O(n67561));   // verilog/uart_rx.v(119[33:55])
    defparam i51875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51173_4_lut (.I0(n41_adj_4605), .I1(n39_adj_4604), .I2(n27_adj_4609), 
            .I3(n65943), .O(n66859));
    defparam i51173_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52029_3_lut (.I0(n22_adj_4617), .I1(baudrate[7]), .I2(n27_adj_4609), 
            .I3(GND_net), .O(n67715));   // verilog/uart_rx.v(119[33:55])
    defparam i52029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51150_3_lut (.I0(n67561), .I1(baudrate[15]), .I2(n43_adj_4603), 
            .I3(GND_net), .O(n66836));   // verilog/uart_rx.v(119[33:55])
    defparam i51150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1026 (.I0(n23), .I1(\o_Rx_DV_N_3488[12] ), .I2(n4940), 
            .I3(GND_net), .O(n60348));   // verilog/uart_rx.v(69[17:62])
    defparam i1_3_lut_adj_1026.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1027 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n27), .I2(n29), 
            .I3(n60348), .O(\r_SM_Main_2__N_3536[1] ));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1027.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i28_3_lut (.I0(n20_adj_4618), .I1(baudrate[9]), 
            .I2(n31_adj_4606), .I3(GND_net), .O(n28_adj_4619));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52409_4_lut (.I0(n28_adj_4619), .I1(n18_adj_4620), .I2(n31_adj_4606), 
            .I3(n65939), .O(n68095));   // verilog/uart_rx.v(119[33:55])
    defparam i52409_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52410_3_lut (.I0(n68095), .I1(baudrate[10]), .I2(n33_adj_4607), 
            .I3(GND_net), .O(n68096));   // verilog/uart_rx.v(119[33:55])
    defparam i52410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52193_3_lut (.I0(n68096), .I1(baudrate[11]), .I2(n35_adj_4608), 
            .I3(GND_net), .O(n67879));   // verilog/uart_rx.v(119[33:55])
    defparam i52193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51175_4_lut (.I0(n41_adj_4605), .I1(n39_adj_4604), .I2(n37_adj_4602), 
            .I3(n67767), .O(n66861));
    defparam i51175_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52188_4_lut (.I0(n66836), .I1(n67715), .I2(n43_adj_4603), 
            .I3(n66859), .O(n67874));   // verilog/uart_rx.v(119[33:55])
    defparam i52188_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51148_3_lut (.I0(n67879), .I1(baudrate[12]), .I2(n37_adj_4602), 
            .I3(GND_net), .O(n66834));   // verilog/uart_rx.v(119[33:55])
    defparam i51148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52499_4_lut (.I0(n66834), .I1(n67874), .I2(n43_adj_4603), 
            .I3(n66861), .O(n68185));   // verilog/uart_rx.v(119[33:55])
    defparam i52499_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52500_3_lut (.I0(n68185), .I1(baudrate[16]), .I2(n2597), 
            .I3(GND_net), .O(n68186));   // verilog/uart_rx.v(119[33:55])
    defparam i52500_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46680_1_lut (.I0(n62350), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n58094));
    defparam i46680_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52963_2_lut_4_lut (.I0(n68188), .I1(baudrate[13]), .I2(n2098), 
            .I3(n25607), .O(n294[10]));   // verilog/uart_rx.v(119[33:55])
    defparam i52963_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1430_i28_3_lut_3_lut (.I0(baudrate[3]), .I1(baudrate[4]), 
            .I2(n2107), .I3(GND_net), .O(n28_adj_4621));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50378_2_lut_4_lut (.I0(n2102), .I1(baudrate[9]), .I2(n2106), 
            .I3(baudrate[5]), .O(n66064));
    defparam i50378_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1430_i30_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[9]), 
            .I2(n2102), .I3(GND_net), .O(n30_adj_4622));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i42443_1_lut (.I0(n25619), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n58082));
    defparam i42443_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i42439_1_lut (.I0(n25622), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n58078));
    defparam i42439_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1028 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4937), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n60696), .O(n60702));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1028.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1029 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n60702), .O(n60708));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1029.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1030 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4937), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n60680), .O(n60686));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1030.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1031 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n60686), .O(n60692));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1031.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1662_3_lut (.I0(n2353), .I1(n8243[23]), .I2(n294[8]), 
            .I3(GND_net), .O(n2476));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1672_3_lut (.I0(n2363), .I1(n8243[13]), .I2(n294[8]), 
            .I3(GND_net), .O(n2486));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1666_3_lut (.I0(n2357), .I1(n8243[19]), .I2(n294[8]), 
            .I3(GND_net), .O(n2480));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i39_2_lut (.I0(n2480), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4623));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1663_3_lut (.I0(n2354), .I1(n8243[22]), .I2(n294[8]), 
            .I3(GND_net), .O(n2477));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i45_2_lut (.I0(n2477), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4624));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1664_3_lut (.I0(n2355), .I1(n8243[21]), .I2(n294[8]), 
            .I3(GND_net), .O(n2478));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i43_2_lut (.I0(n2478), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4625));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1032 (.I0(n60322), .I1(n48_adj_4626), .I2(GND_net), 
            .I3(GND_net), .O(n2491));
    defparam i1_2_lut_adj_1032.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i1667_3_lut (.I0(n2358), .I1(n8243[18]), .I2(n294[8]), 
            .I3(GND_net), .O(n2481));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1668_3_lut (.I0(n2359), .I1(n8243[17]), .I2(n294[8]), 
            .I3(GND_net), .O(n2482));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1669_3_lut (.I0(n2360), .I1(n8243[16]), .I2(n294[8]), 
            .I3(GND_net), .O(n2483));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i33_2_lut (.I0(n2483), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4627));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i35_2_lut (.I0(n2482), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4628));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i37_2_lut (.I0(n2481), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4629));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1665_3_lut (.I0(n2356), .I1(n8243[20]), .I2(n294[8]), 
            .I3(GND_net), .O(n2479));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i41_2_lut (.I0(n2479), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4630));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1671_3_lut (.I0(n2362), .I1(n8243[14]), .I2(n294[8]), 
            .I3(GND_net), .O(n2485));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1670_3_lut (.I0(n2361), .I1(n8243[15]), .I2(n294[8]), 
            .I3(GND_net), .O(n2484));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i29_2_lut (.I0(n2485), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4631));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i31_2_lut (.I0(n2484), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4632));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1676_3_lut (.I0(n2367), .I1(n8243[9]), .I2(n294[8]), 
            .I3(GND_net), .O(n2490));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1674_3_lut (.I0(n2365), .I1(n8243[11]), .I2(n294[8]), 
            .I3(GND_net), .O(n2488));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1675_3_lut (.I0(n2366), .I1(n8243[10]), .I2(n294[8]), 
            .I3(GND_net), .O(n2489));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i21_2_lut (.I0(n2489), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4633));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i23_2_lut (.I0(n2488), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4634));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1673_3_lut (.I0(n2364), .I1(n8243[12]), .I2(n294[8]), 
            .I3(GND_net), .O(n2487));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i25_2_lut (.I0(n2487), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4635));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i27_2_lut (.I0(n2486), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4636));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i19_2_lut (.I0(n2490), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4637));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50319_4_lut (.I0(n25_adj_4635), .I1(n23_adj_4634), .I2(n21_adj_4633), 
            .I3(n19_adj_4637), .O(n66005));
    defparam i50319_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50313_4_lut (.I0(n31_adj_4632), .I1(n29_adj_4631), .I2(n27_adj_4636), 
            .I3(n66005), .O(n65999));
    defparam i50313_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52087_4_lut (.I0(n37_adj_4629), .I1(n35_adj_4628), .I2(n33_adj_4627), 
            .I3(n65999), .O(n67773));
    defparam i52087_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51886_3_lut (.I0(n18_adj_4638), .I1(baudrate[13]), .I2(n41_adj_4630), 
            .I3(GND_net), .O(n67572));   // verilog/uart_rx.v(119[33:55])
    defparam i51886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51887_3_lut (.I0(n67572), .I1(baudrate[14]), .I2(n43_adj_4625), 
            .I3(GND_net), .O(n67573));   // verilog/uart_rx.v(119[33:55])
    defparam i51887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51193_4_lut (.I0(n43_adj_4625), .I1(n41_adj_4630), .I2(n29_adj_4631), 
            .I3(n66003), .O(n66879));
    defparam i51193_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_1685_i26_3_lut (.I0(n24_adj_4639), .I1(baudrate[7]), 
            .I2(n29_adj_4631), .I3(GND_net), .O(n26_adj_4640));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51144_3_lut (.I0(n67573), .I1(baudrate[15]), .I2(n45_adj_4624), 
            .I3(GND_net), .O(n66830));   // verilog/uart_rx.v(119[33:55])
    defparam i51144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i30_3_lut (.I0(n22_adj_4641), .I1(baudrate[9]), 
            .I2(n33_adj_4627), .I3(GND_net), .O(n30_adj_4642));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52407_4_lut (.I0(n30_adj_4642), .I1(n20_adj_4643), .I2(n33_adj_4627), 
            .I3(n65992), .O(n68093));   // verilog/uart_rx.v(119[33:55])
    defparam i52407_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52408_3_lut (.I0(n68093), .I1(baudrate[10]), .I2(n35_adj_4628), 
            .I3(GND_net), .O(n68094));   // verilog/uart_rx.v(119[33:55])
    defparam i52408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52199_3_lut (.I0(n68094), .I1(baudrate[11]), .I2(n37_adj_4629), 
            .I3(GND_net), .O(n67885));   // verilog/uart_rx.v(119[33:55])
    defparam i52199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51197_4_lut (.I0(n43_adj_4625), .I1(n41_adj_4630), .I2(n39_adj_4623), 
            .I3(n67773), .O(n66883));
    defparam i51197_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52026_4_lut (.I0(n66830), .I1(n26_adj_4640), .I2(n45_adj_4624), 
            .I3(n66879), .O(n67712));   // verilog/uart_rx.v(119[33:55])
    defparam i52026_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51142_3_lut (.I0(n67885), .I1(baudrate[12]), .I2(n39_adj_4623), 
            .I3(GND_net), .O(n66828));   // verilog/uart_rx.v(119[33:55])
    defparam i51142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52028_4_lut (.I0(n66828), .I1(n67712), .I2(n45_adj_4624), 
            .I3(n66883), .O(n67714));   // verilog/uart_rx.v(119[33:55])
    defparam i52028_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1579_3_lut (.I0(n2227), .I1(n8217[23]), .I2(n294[9]), 
            .I3(GND_net), .O(n2353));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1580_3_lut (.I0(n2228), .I1(n8217[22]), .I2(n294[9]), 
            .I3(GND_net), .O(n2354));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1581_3_lut (.I0(n2229), .I1(n8217[21]), .I2(n294[9]), 
            .I3(GND_net), .O(n2355));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1582_3_lut (.I0(n2230), .I1(n8217[20]), .I2(n294[9]), 
            .I3(GND_net), .O(n2356));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i41_2_lut (.I0(n2356), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4644));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1583_3_lut (.I0(n2231), .I1(n8217[19]), .I2(n294[9]), 
            .I3(GND_net), .O(n2357));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i39_2_lut (.I0(n2357), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4645));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1584_3_lut (.I0(n2232), .I1(n8217[18]), .I2(n294[9]), 
            .I3(GND_net), .O(n2358));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i37_2_lut (.I0(n2358), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4646));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1585_3_lut (.I0(n2233), .I1(n8217[17]), .I2(n294[9]), 
            .I3(GND_net), .O(n2359));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i35_2_lut (.I0(n2359), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4647));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1586_3_lut (.I0(n2234), .I1(n8217[16]), .I2(n294[9]), 
            .I3(GND_net), .O(n2360));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1588_3_lut (.I0(n2236), .I1(n8217[14]), .I2(n294[9]), 
            .I3(GND_net), .O(n2362));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1587_3_lut (.I0(n2235), .I1(n8217[15]), .I2(n294[9]), 
            .I3(GND_net), .O(n2361));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i29_2_lut (.I0(n2362), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4648));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i31_2_lut (.I0(n2361), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4649));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i42423_1_lut_4_lut (.I0(n61902), .I1(n61904), .I2(n61746), 
            .I3(n61900), .O(n58062));
    defparam i42423_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i50452_3_lut_4_lut (.I0(n1413), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1414), .O(n66138));   // verilog/uart_rx.v(119[33:55])
    defparam i50452_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i33_2_lut (.I0(n2360), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4650));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i24_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2238), .I3(GND_net), .O(n24_adj_4651));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1589_3_lut (.I0(n2237), .I1(n8217[13]), .I2(n294[9]), 
            .I3(GND_net), .O(n2363));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1590_3_lut (.I0(n2238), .I1(n8217[12]), .I2(n294[9]), 
            .I3(GND_net), .O(n2364));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1591_3_lut (.I0(n2239), .I1(n8217[11]), .I2(n294[9]), 
            .I3(GND_net), .O(n2365));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i23_2_lut (.I0(n2365), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4652));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i25_2_lut (.I0(n2364), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4653));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i27_2_lut (.I0(n2363), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4654));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1592_3_lut (.I0(n2240), .I1(n8217[10]), .I2(n294[9]), 
            .I3(GND_net), .O(n2366));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i21_2_lut (.I0(n2366), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4655));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50358_2_lut_4_lut (.I0(n2233), .I1(baudrate[8]), .I2(n2237), 
            .I3(baudrate[4]), .O(n66044));
    defparam i50358_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i50344_4_lut (.I0(n27_adj_4654), .I1(n25_adj_4653), .I2(n23_adj_4652), 
            .I3(n21_adj_4655), .O(n66030));
    defparam i50344_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50340_4_lut (.I0(n33_adj_4650), .I1(n31_adj_4649), .I2(n29_adj_4648), 
            .I3(n66030), .O(n66026));
    defparam i50340_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1517_i26_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2233), .I3(GND_net), .O(n26_adj_4656));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i20_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2367), .I3(GND_net), .O(n20_adj_4657));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i20_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i28_3_lut (.I0(n26_adj_4658), .I1(baudrate[7]), 
            .I2(n31_adj_4649), .I3(GND_net), .O(n28_adj_4659));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i32_3_lut (.I0(n24_adj_4660), .I1(baudrate[9]), 
            .I2(n35_adj_4647), .I3(GND_net), .O(n32_adj_4661));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52405_4_lut (.I0(n32_adj_4661), .I1(n22_adj_4662), .I2(n35_adj_4647), 
            .I3(n66024), .O(n68091));   // verilog/uart_rx.v(119[33:55])
    defparam i52405_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52406_3_lut (.I0(n68091), .I1(baudrate[10]), .I2(n37_adj_4646), 
            .I3(GND_net), .O(n68092));   // verilog/uart_rx.v(119[33:55])
    defparam i52406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52201_3_lut (.I0(n68092), .I1(baudrate[11]), .I2(n39_adj_4645), 
            .I3(GND_net), .O(n67887));   // verilog/uart_rx.v(119[33:55])
    defparam i52201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52089_4_lut (.I0(n39_adj_4645), .I1(n37_adj_4646), .I2(n35_adj_4647), 
            .I3(n66026), .O(n67775));
    defparam i52089_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52469_4_lut (.I0(n28_adj_4659), .I1(n20_adj_4657), .I2(n31_adj_4649), 
            .I3(n66028), .O(n68155));   // verilog/uart_rx.v(119[33:55])
    defparam i52469_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51138_3_lut (.I0(n67887), .I1(baudrate[12]), .I2(n41_adj_4644), 
            .I3(GND_net), .O(n66824));   // verilog/uart_rx.v(119[33:55])
    defparam i51138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52555_4_lut (.I0(n66824), .I1(n68155), .I2(n41_adj_4644), 
            .I3(n67775), .O(n68241));   // verilog/uart_rx.v(119[33:55])
    defparam i52555_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52556_3_lut (.I0(n68241), .I1(baudrate[13]), .I2(n2355), 
            .I3(GND_net), .O(n68242));   // verilog/uart_rx.v(119[33:55])
    defparam i52556_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50366_2_lut_4_lut (.I0(n2235), .I1(baudrate[6]), .I2(n2236), 
            .I3(baudrate[5]), .O(n66052));
    defparam i50366_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i28_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2235), .I3(GND_net), .O(n28_adj_4663));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_965_i36_3_lut_3_lut (.I0(n1413), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n36));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i36_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i52532_3_lut (.I0(n68242), .I1(baudrate[14]), .I2(n2354), 
            .I3(GND_net), .O(n68218));   // verilog/uart_rx.v(119[33:55])
    defparam i52532_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52456_3_lut (.I0(n68218), .I1(baudrate[15]), .I2(n2353), 
            .I3(GND_net), .O(n48_adj_4626));   // verilog/uart_rx.v(119[33:55])
    defparam i52456_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1494_3_lut (.I0(n2098), .I1(n8191[23]), .I2(n294[10]), 
            .I3(GND_net), .O(n2227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1495_3_lut (.I0(n2099), .I1(n8191[22]), .I2(n294[10]), 
            .I3(GND_net), .O(n2228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1496_3_lut (.I0(n2100), .I1(n8191[21]), .I2(n294[10]), 
            .I3(GND_net), .O(n2229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i43_2_lut (.I0(n2229), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4664));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1497_3_lut (.I0(n2101), .I1(n8191[20]), .I2(n294[10]), 
            .I3(GND_net), .O(n2230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i41_2_lut (.I0(n2230), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4665));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1498_3_lut (.I0(n2102), .I1(n8191[19]), .I2(n294[10]), 
            .I3(GND_net), .O(n2231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i39_2_lut (.I0(n2231), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4666));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1499_3_lut (.I0(n2103), .I1(n8191[18]), .I2(n294[10]), 
            .I3(GND_net), .O(n2232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i37_2_lut (.I0(n2232), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4667));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1033 (.I0(n25607), .I1(n48_adj_4668), .I2(baudrate[0]), 
            .I3(GND_net), .O(n2240));
    defparam i1_3_lut_adj_1033.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i1500_3_lut (.I0(n2104), .I1(n8191[17]), .I2(n294[10]), 
            .I3(GND_net), .O(n2233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1502_3_lut (.I0(n2106), .I1(n8191[15]), .I2(n294[10]), 
            .I3(GND_net), .O(n2235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1501_3_lut (.I0(n2105), .I1(n8191[16]), .I2(n294[10]), 
            .I3(GND_net), .O(n2234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i31_2_lut (.I0(n2235), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4669));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i33_2_lut (.I0(n2234), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4670));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i35_2_lut (.I0(n2233), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4671));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1503_3_lut (.I0(n2107), .I1(n8191[14]), .I2(n294[10]), 
            .I3(GND_net), .O(n2236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1504_3_lut (.I0(n2108), .I1(n8191[13]), .I2(n294[10]), 
            .I3(GND_net), .O(n2237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1505_3_lut (.I0(n2109), .I1(n8191[12]), .I2(n294[10]), 
            .I3(GND_net), .O(n2238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i25_2_lut (.I0(n2238), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4672));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i27_2_lut (.I0(n2237), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4673));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i29_2_lut (.I0(n2236), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4674));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1506_3_lut (.I0(n2110), .I1(n8191[11]), .I2(n294[10]), 
            .I3(GND_net), .O(n2239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i23_2_lut (.I0(n2239), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4675));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50368_4_lut (.I0(n29_adj_4674), .I1(n27_adj_4673), .I2(n25_adj_4672), 
            .I3(n23_adj_4675), .O(n66054));
    defparam i50368_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50360_4_lut (.I0(n35_adj_4671), .I1(n33_adj_4670), .I2(n31_adj_4669), 
            .I3(n66054), .O(n66046));
    defparam i50360_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1517_i22_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2240), .I3(GND_net), .O(n22_adj_4676));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i22_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i30_3_lut (.I0(n28_adj_4663), .I1(baudrate[7]), 
            .I2(n33_adj_4670), .I3(GND_net), .O(n30_adj_4677));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i22_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2365), .I3(GND_net), .O(n22_adj_4662));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i42435_1_lut (.I0(n25644), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n58074));
    defparam i42435_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1517_i34_3_lut (.I0(n26_adj_4656), .I1(baudrate[9]), 
            .I2(n37_adj_4667), .I3(GND_net), .O(n34_adj_4678));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52403_4_lut (.I0(n34_adj_4678), .I1(n24_adj_4651), .I2(n37_adj_4667), 
            .I3(n66044), .O(n68089));   // verilog/uart_rx.v(119[33:55])
    defparam i52403_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50338_2_lut_4_lut (.I0(n2360), .I1(baudrate[8]), .I2(n2364), 
            .I3(baudrate[4]), .O(n66024));
    defparam i50338_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i52404_3_lut (.I0(n68089), .I1(baudrate[10]), .I2(n39_adj_4666), 
            .I3(GND_net), .O(n68090));   // verilog/uart_rx.v(119[33:55])
    defparam i52404_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52205_3_lut (.I0(n68090), .I1(baudrate[11]), .I2(n41_adj_4665), 
            .I3(GND_net), .O(n67891));   // verilog/uart_rx.v(119[33:55])
    defparam i52205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i24_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2360), .I3(GND_net), .O(n24_adj_4660));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52093_4_lut (.I0(n41_adj_4665), .I1(n39_adj_4666), .I2(n37_adj_4667), 
            .I3(n66046), .O(n67779));
    defparam i52093_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50342_2_lut_4_lut (.I0(n2362), .I1(baudrate[6]), .I2(n2363), 
            .I3(baudrate[5]), .O(n66028));
    defparam i50342_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i52286_4_lut (.I0(n30_adj_4677), .I1(n22_adj_4676), .I2(n33_adj_4670), 
            .I3(n66052), .O(n67972));   // verilog/uart_rx.v(119[33:55])
    defparam i52286_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51132_3_lut (.I0(n67891), .I1(baudrate[12]), .I2(n43_adj_4664), 
            .I3(GND_net), .O(n66818));   // verilog/uart_rx.v(119[33:55])
    defparam i51132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52369_4_lut (.I0(n66818), .I1(n67972), .I2(n43_adj_4664), 
            .I3(n67779), .O(n68055));   // verilog/uart_rx.v(119[33:55])
    defparam i52369_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52370_3_lut (.I0(n68055), .I1(baudrate[13]), .I2(n2228), 
            .I3(GND_net), .O(n68056));   // verilog/uart_rx.v(119[33:55])
    defparam i52370_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i26_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2362), .I3(GND_net), .O(n26_adj_4658));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1685_i20_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2489), .I3(GND_net), .O(n20_adj_4643));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50306_2_lut_4_lut (.I0(n2484), .I1(baudrate[8]), .I2(n2488), 
            .I3(baudrate[4]), .O(n65992));
    defparam i50306_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1685_i22_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2484), .I3(GND_net), .O(n22_adj_4641));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1685_i24_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2486), .I3(GND_net), .O(n24_adj_4639));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1685_i18_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n60322), .I3(n48_adj_4626), .O(n18_adj_4638));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i18_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i50317_2_lut_4_lut (.I0(n2486), .I1(baudrate[6]), .I2(n2487), 
            .I3(baudrate[5]), .O(n66003));
    defparam i50317_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_4_lut_adj_1034 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4937), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n60792), .O(n60798));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1034.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1035 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n60798), .O(n60804));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1035.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1407_3_lut (.I0(n1966), .I1(n8165[23]), .I2(n294[11]), 
            .I3(GND_net), .O(n2098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1407_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1408_3_lut (.I0(n1967), .I1(n8165[22]), .I2(n294[11]), 
            .I3(GND_net), .O(n2099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1409_3_lut (.I0(n1968), .I1(n8165[21]), .I2(n294[11]), 
            .I3(GND_net), .O(n2100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1413_3_lut (.I0(n1972), .I1(n8165[17]), .I2(n294[11]), 
            .I3(GND_net), .O(n2104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1412_3_lut (.I0(n1971), .I1(n8165[18]), .I2(n294[11]), 
            .I3(GND_net), .O(n2103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i35_2_lut (.I0(n2104), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4679));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i37_2_lut (.I0(n2103), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4680));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1418_3_lut (.I0(n1977), .I1(n8165[12]), .I2(n294[11]), 
            .I3(GND_net), .O(n2109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1410_3_lut (.I0(n1969), .I1(n8165[20]), .I2(n294[11]), 
            .I3(GND_net), .O(n2101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i41_2_lut (.I0(n2101), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4681));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1411_3_lut (.I0(n1970), .I1(n8165[19]), .I2(n294[11]), 
            .I3(GND_net), .O(n2102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i39_2_lut (.I0(n2102), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4682));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1415_3_lut (.I0(n1974), .I1(n8165[15]), .I2(n294[11]), 
            .I3(GND_net), .O(n2106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1414_3_lut (.I0(n1973), .I1(n8165[16]), .I2(n294[11]), 
            .I3(GND_net), .O(n2105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1416_3_lut (.I0(n1975), .I1(n8165[14]), .I2(n294[11]), 
            .I3(GND_net), .O(n2107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46649_1_lut_2_lut (.I0(baudrate[17]), .I1(n25619), .I2(GND_net), 
            .I3(GND_net), .O(n58086));
    defparam i46649_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_37_LessThan_1430_i29_2_lut (.I0(n2107), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4683));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i31_2_lut (.I0(n2106), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4684));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i33_2_lut (.I0(n2105), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4685));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1417_3_lut (.I0(n1976), .I1(n8165[13]), .I2(n294[11]), 
            .I3(GND_net), .O(n2108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1036 (.I0(baudrate[27]), .I1(baudrate[24]), .I2(baudrate[29]), 
            .I3(baudrate[30]), .O(n61800));
    defparam i1_4_lut_adj_1036.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1037 (.I0(n61750), .I1(n61798), .I2(n60848), 
            .I3(GND_net), .O(n61808));
    defparam i1_3_lut_adj_1037.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1038 (.I0(n61808), .I1(n61804), .I2(n61806), 
            .I3(n61800), .O(n25607));
    defparam i1_4_lut_adj_1038.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1430_i27_2_lut (.I0(n2108), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4686));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1039 (.I0(n23), .I1(\o_Rx_DV_N_3488[12] ), .I2(n4937), 
            .I3(\o_Rx_DV_N_3488[8] ), .O(n60306));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1039.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1040 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n27), .I2(n29), 
            .I3(n60306), .O(r_SM_Main_2__N_3446[1]));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1040.LUT_INIT = 16'hfffe;
    SB_LUT4 i50386_4_lut (.I0(n33_adj_4685), .I1(n31_adj_4684), .I2(n29_adj_4683), 
            .I3(n27_adj_4686), .O(n66072));
    defparam i50386_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_4_lut_adj_1041 (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), 
            .I2(\o_Rx_DV_N_3488[2] ), .I3(\o_Rx_DV_N_3488[1] ), .O(n61386));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1041.LUT_INIT = 16'h7bde;
    SB_LUT4 equal_267_i3_2_lut (.I0(r_Clock_Count[2]), .I1(\o_Rx_DV_N_3488[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4687));   // verilog/uart_rx.v(69[17:62])
    defparam equal_267_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i38_3_lut (.I0(n30_adj_4622), .I1(baudrate[10]), 
            .I2(n41_adj_4681), .I3(GND_net), .O(n38_adj_4688));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28992_rep_4_2_lut (.I0(n8165[11]), .I1(n294[11]), .I2(GND_net), 
            .I3(GND_net), .O(n58097));   // verilog/uart_rx.v(119[33:55])
    defparam i28992_rep_4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1042 (.I0(r_Clock_Count[3]), .I1(n3_adj_4687), 
            .I2(\o_Rx_DV_N_3488[4] ), .I3(n61386), .O(n61390));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1042.LUT_INIT = 16'hffde;
    SB_LUT4 equal_267_i5_2_lut (.I0(r_Clock_Count[4]), .I1(\o_Rx_DV_N_3488[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/uart_rx.v(69[17:62])
    defparam equal_267_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i26_4_lut (.I0(n58097), .I1(baudrate[2]), 
            .I2(n2109), .I3(baudrate[1]), .O(n26_adj_4689));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i26_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i51902_3_lut (.I0(n26_adj_4689), .I1(baudrate[6]), .I2(n33_adj_4685), 
            .I3(GND_net), .O(n67588));   // verilog/uart_rx.v(119[33:55])
    defparam i51902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1043 (.I0(r_Clock_Count[5]), .I1(n5), .I2(\o_Rx_DV_N_3488[6] ), 
            .I3(n61390), .O(n61394));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1043.LUT_INIT = 16'hffde;
    SB_LUT4 equal_267_i8_2_lut (.I0(r_Clock_Count[7]), .I1(\o_Rx_DV_N_3488[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4690));   // verilog/uart_rx.v(69[17:62])
    defparam equal_267_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i51903_3_lut (.I0(n67588), .I1(baudrate[7]), .I2(n35_adj_4679), 
            .I3(GND_net), .O(n67589));   // verilog/uart_rx.v(119[33:55])
    defparam i51903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50380_4_lut (.I0(n39_adj_4682), .I1(n37_adj_4680), .I2(n35_adj_4679), 
            .I3(n66072), .O(n66066));
    defparam i50380_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52401_4_lut (.I0(n38_adj_4688), .I1(n28_adj_4621), .I2(n41_adj_4681), 
            .I3(n66064), .O(n68087));   // verilog/uart_rx.v(119[33:55])
    defparam i52401_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51118_3_lut (.I0(n67589), .I1(baudrate[8]), .I2(n37_adj_4680), 
            .I3(GND_net), .O(n66804));   // verilog/uart_rx.v(119[33:55])
    defparam i51118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1044 (.I0(r_Clock_Count[6]), .I1(n8_adj_4690), 
            .I2(n61394), .I3(\o_Rx_DV_N_3488[7] ), .O(n56722));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1044.LUT_INIT = 16'hfdfe;
    SB_LUT4 i52567_4_lut (.I0(n66804), .I1(n68087), .I2(n41_adj_4681), 
            .I3(n66066), .O(n68253));   // verilog/uart_rx.v(119[33:55])
    defparam i52567_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52568_3_lut (.I0(n68253), .I1(baudrate[11]), .I2(n2100), 
            .I3(GND_net), .O(n68254));   // verilog/uart_rx.v(119[33:55])
    defparam i52568_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52502_3_lut (.I0(n68254), .I1(baudrate[12]), .I2(n2099), 
            .I3(GND_net), .O(n68188));   // verilog/uart_rx.v(119[33:55])
    defparam i52502_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51124_3_lut (.I0(n68188), .I1(baudrate[13]), .I2(n2098), 
            .I3(GND_net), .O(n48_adj_4668));   // verilog/uart_rx.v(119[33:55])
    defparam i51124_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n58912));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 div_37_i1318_3_lut (.I0(n1831), .I1(n8139[23]), .I2(n294[12]), 
            .I3(GND_net), .O(n1966));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1319_3_lut (.I0(n1832), .I1(n8139[22]), .I2(n294[12]), 
            .I3(GND_net), .O(n1967));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1320_3_lut (.I0(n1833), .I1(n8139[21]), .I2(n294[12]), 
            .I3(GND_net), .O(n1968));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1323_3_lut (.I0(n1836), .I1(n8139[18]), .I2(n294[12]), 
            .I3(GND_net), .O(n1971));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i37_2_lut (.I0(n1971), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4691));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1324_3_lut (.I0(n1837), .I1(n8139[17]), .I2(n294[12]), 
            .I3(GND_net), .O(n1972));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i35_2_lut (.I0(n1972), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4692));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1321_3_lut (.I0(n1834), .I1(n8139[20]), .I2(n294[12]), 
            .I3(GND_net), .O(n1969));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i41_2_lut (.I0(n1969), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4693));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1325_3_lut (.I0(n1838), .I1(n8139[16]), .I2(n294[12]), 
            .I3(GND_net), .O(n1973));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1327_3_lut (.I0(n1840), .I1(n8139[14]), .I2(n294[12]), 
            .I3(GND_net), .O(n1975));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i29_2_lut (.I0(n1975), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4694));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i33_2_lut (.I0(n1973), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4695));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1322_3_lut (.I0(n1835), .I1(n8139[19]), .I2(n294[12]), 
            .I3(GND_net), .O(n1970));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1326_3_lut (.I0(n1839), .I1(n8139[15]), .I2(n294[12]), 
            .I3(GND_net), .O(n1974));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i31_2_lut (.I0(n1974), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4696));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i39_2_lut (.I0(n1970), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4697));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1328_3_lut (.I0(n1841), .I1(n8139[13]), .I2(n294[12]), 
            .I3(GND_net), .O(n1976));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i27_2_lut (.I0(n1976), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50400_4_lut (.I0(n33_adj_4695), .I1(n31_adj_4696), .I2(n29_adj_4694), 
            .I3(n27_adj_4698), .O(n66086));
    defparam i50400_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1341_i38_3_lut (.I0(n30_adj_4601), .I1(baudrate[9]), 
            .I2(n41_adj_4693), .I3(GND_net), .O(n38_adj_4699));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i26_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1977), .I3(GND_net), .O(n26_adj_4700));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51906_3_lut (.I0(n26_adj_4700), .I1(baudrate[5]), .I2(n33_adj_4695), 
            .I3(GND_net), .O(n67592));   // verilog/uart_rx.v(119[33:55])
    defparam i51906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51907_3_lut (.I0(n67592), .I1(baudrate[6]), .I2(n35_adj_4692), 
            .I3(GND_net), .O(n67593));   // verilog/uart_rx.v(119[33:55])
    defparam i51907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50396_4_lut (.I0(n39_adj_4697), .I1(n37_adj_4691), .I2(n35_adj_4692), 
            .I3(n66086), .O(n66082));
    defparam i50396_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1766_i18_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2610), .I3(GND_net), .O(n18_adj_4620));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52399_4_lut (.I0(n38_adj_4699), .I1(n28), .I2(n41_adj_4693), 
            .I3(n66080), .O(n68085));   // verilog/uart_rx.v(119[33:55])
    defparam i52399_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i51106_3_lut (.I0(n67593), .I1(baudrate[7]), .I2(n37_adj_4691), 
            .I3(GND_net), .O(n66792));   // verilog/uart_rx.v(119[33:55])
    defparam i51106_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52565_4_lut (.I0(n66792), .I1(n68085), .I2(n41_adj_4693), 
            .I3(n66082), .O(n68251));   // verilog/uart_rx.v(119[33:55])
    defparam i52565_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52566_3_lut (.I0(n68251), .I1(baudrate[10]), .I2(n1968), 
            .I3(GND_net), .O(n68252));   // verilog/uart_rx.v(119[33:55])
    defparam i52566_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52508_3_lut (.I0(n68252), .I1(baudrate[11]), .I2(n1967), 
            .I3(GND_net), .O(n68194));   // verilog/uart_rx.v(119[33:55])
    defparam i52508_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50253_2_lut_4_lut (.I0(n2605), .I1(baudrate[8]), .I2(n2609), 
            .I3(baudrate[4]), .O(n65939));
    defparam i50253_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51112_3_lut (.I0(n68194), .I1(baudrate[12]), .I2(n1966), 
            .I3(GND_net), .O(n48_adj_4502));   // verilog/uart_rx.v(119[33:55])
    defparam i51112_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1766_i20_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2605), .I3(GND_net), .O(n20_adj_4618));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1045 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4937), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n58912), .O(n60440));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1045.LUT_INIT = 16'hfeff;
    SB_LUT4 div_37_LessThan_1766_i22_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2607), .I3(GND_net), .O(n22_adj_4617));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1046 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n60440), .O(n60446));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1046.LUT_INIT = 16'hfffe;
    SB_LUT4 i46823_2_lut (.I0(\o_Rx_DV_N_3488[12] ), .I1(n56722), .I2(GND_net), 
            .I3(GND_net), .O(n62500));
    defparam i46823_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i46919_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n62500), .O(n62596));
    defparam i46919_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i2_4_lut (.I0(n60446), .I1(r_SM_Main_2__N_3446[1]), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n2));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i2_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 i50257_2_lut_4_lut (.I0(n2607), .I1(baudrate[6]), .I2(n2608), 
            .I3(baudrate[5]), .O(n65943));
    defparam i50257_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1227_3_lut (.I0(n1693), .I1(n8113[23]), .I2(n294[13]), 
            .I3(GND_net), .O(n1831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1233_3_lut (.I0(n1699), .I1(n8113[17]), .I2(n294[13]), 
            .I3(GND_net), .O(n1837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1228_3_lut (.I0(n1694), .I1(n8113[22]), .I2(n294[13]), 
            .I3(GND_net), .O(n1832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1231_3_lut (.I0(n1697), .I1(n8113[19]), .I2(n294[13]), 
            .I3(GND_net), .O(n1835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1232_3_lut (.I0(n1698), .I1(n8113[18]), .I2(n294[13]), 
            .I3(GND_net), .O(n1836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i1_4_lut (.I0(r_Rx_Data), .I1(n62596), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n11645));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i3_3_lut (.I0(n11645), .I1(n2), .I2(\r_SM_Main[1] ), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i3_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 div_37_LessThan_1250_i37_2_lut (.I0(n1836), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4701));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i39_2_lut (.I0(n1835), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4702));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1229_3_lut (.I0(n1695), .I1(n8113[21]), .I2(n294[13]), 
            .I3(GND_net), .O(n1833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i43_2_lut (.I0(n1833), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4703));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1047 (.I0(n25639), .I1(n48_adj_4704), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1841));
    defparam i1_3_lut_adj_1047.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i1236_3_lut (.I0(n1702), .I1(n8113[14]), .I2(n294[13]), 
            .I3(GND_net), .O(n1840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1230_3_lut (.I0(n1696), .I1(n8113[20]), .I2(n294[13]), 
            .I3(GND_net), .O(n1834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i41_2_lut (.I0(n1834), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4705));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1234_3_lut (.I0(n1700), .I1(n8113[16]), .I2(n294[13]), 
            .I3(GND_net), .O(n1838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1235_3_lut (.I0(n1701), .I1(n8113[15]), .I2(n294[13]), 
            .I3(GND_net), .O(n1839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i31_2_lut (.I0(n1839), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4706));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i33_2_lut (.I0(n1838), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4707));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i35_2_lut (.I0(n1837), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4708));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i29_2_lut (.I0(n1840), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4709));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50416_4_lut (.I0(n35_adj_4708), .I1(n33_adj_4707), .I2(n31_adj_4706), 
            .I3(n29_adj_4709), .O(n66102));
    defparam i50416_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1845_i16_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2728), .I3(GND_net), .O(n16_adj_4600));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50216_2_lut_4_lut (.I0(n2723), .I1(baudrate[8]), .I2(n2727), 
            .I3(baudrate[4]), .O(n65902));
    defparam i50216_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1250_i40_3_lut (.I0(n32_adj_4557), .I1(baudrate[9]), 
            .I2(n43_adj_4703), .I3(GND_net), .O(n40_adj_4710));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i28_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1841), .I3(GND_net), .O(n28_adj_4711));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i28_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51908_3_lut (.I0(n28_adj_4711), .I1(baudrate[5]), .I2(n35_adj_4708), 
            .I3(GND_net), .O(n67594));   // verilog/uart_rx.v(119[33:55])
    defparam i51908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51909_3_lut (.I0(n67594), .I1(baudrate[6]), .I2(n37_adj_4701), 
            .I3(GND_net), .O(n67595));   // verilog/uart_rx.v(119[33:55])
    defparam i51909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50412_4_lut (.I0(n41_adj_4705), .I1(n39_adj_4702), .I2(n37_adj_4701), 
            .I3(n66102), .O(n66098));
    defparam i50412_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52371_4_lut (.I0(n40_adj_4710), .I1(n30_adj_4555), .I2(n43_adj_4703), 
            .I3(n66094), .O(n68057));   // verilog/uart_rx.v(119[33:55])
    defparam i52371_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_1845_i18_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2723), .I3(GND_net), .O(n18_adj_4598));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i20_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2725), .I3(GND_net), .O(n20_adj_4597));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51104_3_lut (.I0(n67595), .I1(baudrate[7]), .I2(n39_adj_4702), 
            .I3(GND_net), .O(n66790));   // verilog/uart_rx.v(119[33:55])
    defparam i51104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52595_4_lut (.I0(n66790), .I1(n68057), .I2(n43_adj_4703), 
            .I3(n66098), .O(n68281));   // verilog/uart_rx.v(119[33:55])
    defparam i52595_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52596_3_lut (.I0(n68281), .I1(baudrate[10]), .I2(n1832), 
            .I3(GND_net), .O(n68282));   // verilog/uart_rx.v(119[33:55])
    defparam i52596_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50194_2_lut_4_lut (.I0(n2715), .I1(baudrate[16]), .I2(n2724), 
            .I3(baudrate[7]), .O(n65880));
    defparam i50194_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1845_i22_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2715), .I3(GND_net), .O(n22_adj_4595));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1922_i14_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2843), .I3(GND_net), .O(n14_adj_4578));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50175_2_lut_4_lut (.I0(n2838), .I1(baudrate[8]), .I2(n2842), 
            .I3(baudrate[4]), .O(n65861));
    defparam i50175_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1134_3_lut (.I0(n1552), .I1(n8087[23]), .I2(n294[14]), 
            .I3(GND_net), .O(n1693));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i16_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2838), .I3(GND_net), .O(n16_adj_4576));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1135_3_lut (.I0(n1553), .I1(n8087[22]), .I2(n294[14]), 
            .I3(GND_net), .O(n1694));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1136_3_lut (.I0(n1554), .I1(n8087[21]), .I2(n294[14]), 
            .I3(GND_net), .O(n1695));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i18_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2840), .I3(GND_net), .O(n18_adj_4575));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50148_2_lut_4_lut (.I0(n2830), .I1(baudrate[16]), .I2(n2839), 
            .I3(baudrate[7]), .O(n65834));
    defparam i50148_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1157_i43_2_lut (.I0(n1695), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4712));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1139_3_lut (.I0(n1557), .I1(n8087[18]), .I2(n294[14]), 
            .I3(GND_net), .O(n1698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1137_3_lut (.I0(n1555), .I1(n8087[20]), .I2(n294[14]), 
            .I3(GND_net), .O(n1696));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i37_2_lut (.I0(n1698), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4713));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i20_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2830), .I3(GND_net), .O(n20_adj_4573));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46894_1_lut_2_lut (.I0(baudrate[8]), .I1(n62568), .I2(GND_net), 
            .I3(GND_net), .O(n58116));
    defparam i46894_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_37_LessThan_1157_i41_2_lut (.I0(n1696), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4714));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1142_3_lut (.I0(n1560), .I1(n8087[15]), .I2(n294[14]), 
            .I3(GND_net), .O(n1701));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1138_3_lut (.I0(n1556), .I1(n8087[19]), .I2(n294[14]), 
            .I3(GND_net), .O(n1697));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1157_i39_2_lut (.I0(n1697), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4715));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1140_3_lut (.I0(n1558), .I1(n8087[17]), .I2(n294[14]), 
            .I3(GND_net), .O(n1699));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1141_3_lut (.I0(n1559), .I1(n8087[16]), .I2(n294[14]), 
            .I3(GND_net), .O(n1700));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1048 (.I0(baudrate[27]), .I1(baudrate[28]), .I2(GND_net), 
            .I3(GND_net), .O(n61746));
    defparam i1_2_lut_adj_1048.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1049 (.I0(n61790), .I1(n61746), .I2(n61748), 
            .I3(baudrate[11]), .O(n61776));
    defparam i1_4_lut_adj_1049.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1050 (.I0(n61776), .I1(n61778), .I2(n61766), 
            .I3(n61644), .O(n25639));
    defparam i1_4_lut_adj_1050.LUT_INIT = 16'hfffe;
    SB_LUT4 i28985_rep_5_2_lut (.I0(n8087[14]), .I1(n294[14]), .I2(GND_net), 
            .I3(GND_net), .O(n58106));   // verilog/uart_rx.v(119[33:55])
    defparam i28985_rep_5_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1157_i32_4_lut (.I0(n58106), .I1(baudrate[2]), 
            .I2(n1701), .I3(baudrate[1]), .O(n32_adj_4716));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i32_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i51912_3_lut (.I0(n32_adj_4716), .I1(baudrate[6]), .I2(n39_adj_4715), 
            .I3(GND_net), .O(n67598));   // verilog/uart_rx.v(119[33:55])
    defparam i51912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51913_3_lut (.I0(n67598), .I1(baudrate[7]), .I2(n41_adj_4714), 
            .I3(GND_net), .O(n67599));   // verilog/uart_rx.v(119[33:55])
    defparam i51913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51319_4_lut (.I0(n41_adj_4714), .I1(n39_adj_4715), .I2(n37_adj_4713), 
            .I3(n66116), .O(n67005));
    defparam i51319_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52016_3_lut (.I0(n34_adj_4717), .I1(baudrate[5]), .I2(n37_adj_4713), 
            .I3(GND_net), .O(n67702));   // verilog/uart_rx.v(119[33:55])
    defparam i52016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i12_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2955), .I3(GND_net), .O(n12_adj_4554));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50114_2_lut_4_lut (.I0(n2950), .I1(baudrate[8]), .I2(n2954), 
            .I3(baudrate[4]), .O(n65800));
    defparam i50114_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i51099_3_lut (.I0(n67599), .I1(baudrate[8]), .I2(n43_adj_4712), 
            .I3(GND_net), .O(n66785));   // verilog/uart_rx.v(119[33:55])
    defparam i51099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52216_4_lut (.I0(n66785), .I1(n67702), .I2(n43_adj_4712), 
            .I3(n67005), .O(n67902));   // verilog/uart_rx.v(119[33:55])
    defparam i52216_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_1997_i14_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2950), .I3(GND_net), .O(n14_adj_4553));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i52217_3_lut (.I0(n67902), .I1(baudrate[9]), .I2(n1694), .I3(GND_net), 
            .O(n67903));   // verilog/uart_rx.v(119[33:55])
    defparam i52217_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1157_i48_3_lut (.I0(n67903), .I1(baudrate[10]), 
            .I2(n1693), .I3(GND_net), .O(n48_adj_4704));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1997_i16_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2952), .I3(GND_net), .O(n16_adj_4552));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50100_2_lut_4_lut (.I0(n2942), .I1(baudrate[16]), .I2(n2951), 
            .I3(baudrate[7]), .O(n65786));
    defparam i50100_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1997_i18_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2942), .I3(GND_net), .O(n18));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i10_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3064), .I3(GND_net), .O(n10_adj_4532));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i14_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3061), .I3(GND_net), .O(n14_adj_4531));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50042_2_lut_4_lut (.I0(n3051), .I1(baudrate[16]), .I2(n3060), 
            .I3(baudrate[7]), .O(n65728));
    defparam i50042_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2070_i16_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3051), .I3(GND_net), .O(n16_adj_4529));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i12_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3059), .I3(GND_net), .O(n12_adj_4533));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50071_2_lut_4_lut (.I0(n3059), .I1(baudrate[8]), .I2(n3063), 
            .I3(baudrate[4]), .O(n65757));
    defparam i50071_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i46679_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n25619), .I3(baudrate[15]), .O(n62350));
    defparam i46679_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53432_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n25619), .I3(n48_adj_4626), .O(n294[8]));
    defparam i53432_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i46656_1_lut_2_lut_3_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n25619), .I3(GND_net), .O(n58090));
    defparam i46656_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i46869_2_lut_3_lut_4_lut (.I0(baudrate[13]), .I1(baudrate[14]), 
            .I2(n62350), .I3(baudrate[12]), .O(n62546));
    defparam i46869_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i53426_2_lut_3_lut_4_lut (.I0(baudrate[13]), .I1(baudrate[14]), 
            .I2(n62350), .I3(n48_adj_4502), .O(n294[11]));
    defparam i53426_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i46898_1_lut (.I0(n62574), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n58070));
    defparam i46898_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i53470_2_lut_4_lut (.I0(n68108), .I1(baudrate[22]), .I2(n3151), 
            .I3(n25552), .O(n294[1]));
    defparam i53470_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_2141_i8_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3170), .I3(GND_net), .O(n8_adj_4503));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46891_2_lut_3_lut_4_lut (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(n62546), .I3(baudrate[9]), .O(n62568));
    defparam i46891_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2141_i12_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3167), .I3(GND_net), .O(n12_adj_4501));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49974_2_lut_4_lut (.I0(n3157), .I1(baudrate[16]), .I2(n3166), 
            .I3(baudrate[7]), .O(n65660));
    defparam i49974_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2141_i14_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3157), .I3(GND_net), .O(n14_adj_4500));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i10_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3165), .I3(GND_net), .O(n10_adj_4507));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1039_3_lut (.I0(n1408), .I1(n8061[23]), .I2(n294[15]), 
            .I3(GND_net), .O(n1552));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1040_3_lut (.I0(n1409), .I1(n8061[22]), .I2(n294[15]), 
            .I3(GND_net), .O(n1553));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1044_3_lut (.I0(n1413), .I1(n8061[18]), .I2(n294[15]), 
            .I3(GND_net), .O(n1557));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i37_2_lut (.I0(n1557), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4718));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50010_2_lut_4_lut (.I0(n3165), .I1(baudrate[8]), .I2(n3169), 
            .I3(baudrate[4]), .O(n65696));
    defparam i50010_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1045_3_lut (.I0(n1414), .I1(n8061[17]), .I2(n294[15]), 
            .I3(GND_net), .O(n1558));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1043_3_lut (.I0(n1412), .I1(n8061[19]), .I2(n294[15]), 
            .I3(GND_net), .O(n1556));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i53417_2_lut_3_lut_4_lut (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(n62546), .I3(n48_adj_4498), .O(n294[14]));
    defparam i53417_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_3_lut_adj_1051 (.I0(baudrate[26]), .I1(baudrate[30]), 
            .I2(baudrate[23]), .I3(GND_net), .O(n61904));
    defparam i1_2_lut_3_lut_adj_1051.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_LessThan_1062_i39_2_lut (.I0(n1556), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4719));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i53401_2_lut_3_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n62572), .I3(n48_adj_4470), .O(n294[19]));
    defparam i53401_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i46855_2_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), .I2(baudrate[7]), 
            .I3(baudrate[8]), .O(n62532));
    defparam i46855_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1041_3_lut (.I0(n1410), .I1(n8061[21]), .I2(n294[15]), 
            .I3(GND_net), .O(n1554));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i43_2_lut (.I0(n1554), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4720));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1046_3_lut (.I0(n1415), .I1(n8061[16]), .I2(n294[15]), 
            .I3(GND_net), .O(n1559));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1042_3_lut (.I0(n1411), .I1(n8061[20]), .I2(n294[15]), 
            .I3(GND_net), .O(n1555));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1062_i41_2_lut (.I0(n1555), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4721));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i32_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1560), .I3(GND_net), .O(n32_adj_4722));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i32_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i51916_3_lut (.I0(n32_adj_4722), .I1(baudrate[5]), .I2(n39_adj_4719), 
            .I3(GND_net), .O(n67602));   // verilog/uart_rx.v(119[33:55])
    defparam i51916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51917_3_lut (.I0(n67602), .I1(baudrate[6]), .I2(n41_adj_4721), 
            .I3(GND_net), .O(n67603));   // verilog/uart_rx.v(119[33:55])
    defparam i51917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51327_4_lut (.I0(n41_adj_4721), .I1(n39_adj_4719), .I2(n37_adj_4718), 
            .I3(n66128), .O(n67013));
    defparam i51327_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52012_3_lut (.I0(n34_adj_4723), .I1(baudrate[4]), .I2(n37_adj_4718), 
            .I3(GND_net), .O(n67698));   // verilog/uart_rx.v(119[33:55])
    defparam i52012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51094_3_lut (.I0(n67603), .I1(baudrate[7]), .I2(n43_adj_4720), 
            .I3(GND_net), .O(n66780));   // verilog/uart_rx.v(119[33:55])
    defparam i51094_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52218_4_lut (.I0(n66780), .I1(n67698), .I2(n43_adj_4720), 
            .I3(n67013), .O(n67904));   // verilog/uart_rx.v(119[33:55])
    defparam i52218_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i52219_3_lut (.I0(n67904), .I1(baudrate[8]), .I2(n1553), .I3(GND_net), 
            .O(n67905));   // verilog/uart_rx.v(119[33:55])
    defparam i52219_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1062_i48_3_lut (.I0(n67905), .I1(baudrate[9]), 
            .I2(n1552), .I3(GND_net), .O(n48_adj_4498));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i48_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4724));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_4_lut_adj_1052 (.I0(baudrate[28]), .I1(baudrate[25]), 
            .I2(baudrate[26]), .I3(baudrate[29]), .O(n60294));
    defparam i1_3_lut_4_lut_adj_1052.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1053 (.I0(baudrate[20]), .I1(baudrate[21]), 
            .I2(baudrate[22]), .I3(baudrate[23]), .O(n61804));
    defparam i1_2_lut_4_lut_adj_1053.LUT_INIT = 16'hfffe;
    SB_LUT4 i46795_2_lut_3_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(baudrate[4]), 
            .I3(GND_net), .O(n62472));
    defparam i46795_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_4_lut_adj_1054 (.I0(baudrate[12]), .I1(baudrate[13]), 
            .I2(baudrate[14]), .I3(baudrate[15]), .O(n60966));
    defparam i1_2_lut_4_lut_adj_1054.LUT_INIT = 16'hfffe;
    SB_LUT4 i50638_2_lut_3_lut (.I0(n25589), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n65404));   // verilog/uart_rx.v(119[33:55])
    defparam i50638_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_2_lut_4_lut_adj_1055 (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(baudrate[18]), .I3(baudrate[19]), .O(n61806));
    defparam i1_2_lut_4_lut_adj_1055.LUT_INIT = 16'hfffe;
    SB_LUT4 i50028_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_4466), .I2(n25589), 
            .I3(GND_net), .O(n65714));   // verilog/uart_rx.v(119[33:55])
    defparam i50028_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_4_lut_adj_1056 (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(baudrate[12]), .I3(baudrate[13]), .O(n61656));
    defparam i1_2_lut_4_lut_adj_1056.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1057 (.I0(baudrate[6]), .I1(baudrate[7]), 
            .I2(baudrate[8]), .I3(baudrate[9]), .O(n61658));
    defparam i1_2_lut_4_lut_adj_1057.LUT_INIT = 16'hfffe;
    SB_LUT4 i46895_2_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[8]), .I2(n62568), 
            .I3(GND_net), .O(n62572));
    defparam i46895_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_4_lut_adj_1058 (.I0(n25589), .I1(n48_adj_4466), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n44_adj_4467));
    defparam i1_3_lut_4_lut_adj_1058.LUT_INIT = 16'hefff;
    SB_LUT4 i50034_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_4468), .I2(n25632), 
            .I3(GND_net), .O(n65720));   // verilog/uart_rx.v(119[33:55])
    defparam i50034_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i50648_4_lut (.I0(\o_Rx_DV_N_3488[8] ), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n4937), .I3(n56959), .O(n65352));
    defparam i50648_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i50643_4_lut (.I0(n65352), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n65349));
    defparam i50643_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i14_4_lut (.I0(\r_SM_Main[1] ), .I1(n65349), .I2(r_SM_Main[0]), 
            .I3(n27), .O(n27724));
    defparam i14_4_lut.LUT_INIT = 16'h05c5;
    SB_LUT4 i1_4_lut_adj_1059 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n4937), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n60760), .O(n60766));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1059.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1060 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n60766), .O(n60772));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1060.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1061 (.I0(baudrate[9]), .I1(baudrate[10]), .I2(GND_net), 
            .I3(GND_net), .O(n60826));
    defparam i1_2_lut_adj_1061.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1062 (.I0(baudrate[5]), .I1(baudrate[6]), .I2(GND_net), 
            .I3(GND_net), .O(n60830));
    defparam i1_2_lut_adj_1062.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1063 (.I0(baudrate[7]), .I1(baudrate[8]), .I2(GND_net), 
            .I3(GND_net), .O(n60828));
    defparam i1_2_lut_adj_1063.LUT_INIT = 16'heeee;
    SB_LUT4 i46827_2_lut (.I0(baudrate[3]), .I1(baudrate[4]), .I2(GND_net), 
            .I3(GND_net), .O(n62504));
    defparam i46827_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1064 (.I0(baudrate[29]), .I1(baudrate[24]), .I2(GND_net), 
            .I3(GND_net), .O(n61748));
    defparam i1_2_lut_adj_1064.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1065 (.I0(baudrate[20]), .I1(baudrate[21]), .I2(GND_net), 
            .I3(GND_net), .O(n61792));
    defparam i1_2_lut_adj_1065.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1066 (.I0(baudrate[31]), .I1(baudrate[26]), .I2(GND_net), 
            .I3(GND_net), .O(n61750));
    defparam i1_2_lut_adj_1066.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1067 (.I0(baudrate[28]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n60848));
    defparam i1_2_lut_adj_1067.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1068 (.I0(baudrate[27]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n61666));
    defparam i1_2_lut_adj_1068.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1069 (.I0(baudrate[22]), .I1(baudrate[23]), .I2(GND_net), 
            .I3(GND_net), .O(n61790));
    defparam i1_2_lut_adj_1069.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1070 (.I0(n61790), .I1(n61666), .I2(n60848), 
            .I3(baudrate[19]), .O(n60868));
    defparam i1_4_lut_adj_1070.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1071 (.I0(n60868), .I1(n61750), .I2(n61792), 
            .I3(n61748), .O(n25622));
    defparam i1_4_lut_adj_1071.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1072 (.I0(baudrate[17]), .I1(baudrate[18]), .I2(GND_net), 
            .I3(GND_net), .O(n62450));
    defparam i1_2_lut_adj_1072.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1073 (.I0(baudrate[13]), .I1(baudrate[14]), .I2(GND_net), 
            .I3(GND_net), .O(n60822));
    defparam i1_2_lut_adj_1073.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1074 (.I0(baudrate[15]), .I1(baudrate[16]), .I2(GND_net), 
            .I3(GND_net), .O(n60820));
    defparam i1_2_lut_adj_1074.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1075 (.I0(baudrate[11]), .I1(baudrate[12]), .I2(GND_net), 
            .I3(GND_net), .O(n60824));
    defparam i1_2_lut_adj_1075.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1076 (.I0(n60824), .I1(n60820), .I2(n60822), 
            .I3(n62450), .O(n60842));
    defparam i1_4_lut_adj_1076.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1077 (.I0(n62504), .I1(n60828), .I2(n60830), 
            .I3(n60826), .O(n60844));
    defparam i1_4_lut_adj_1077.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1078 (.I0(n60844), .I1(n25622), .I2(n60842), 
            .I3(GND_net), .O(n25589));
    defparam i1_3_lut_adj_1078.LUT_INIT = 16'hfefe;
    SB_LUT4 i52763_3_lut (.I0(n25589), .I1(baudrate[1]), .I2(baudrate[2]), 
            .I3(GND_net), .O(n25530));   // verilog/uart_rx.v(119[33:55])
    defparam i52763_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i42427_1_lut (.I0(n25629), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n58066));
    defparam i42427_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_4_lut_adj_1079 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n60712));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1079.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_3_lut_4_lut_adj_1080 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n60792));   // verilog/uart_rx.v(98[17:39])
    defparam i1_3_lut_4_lut_adj_1080.LUT_INIT = 16'hfffb;
    SB_LUT4 div_37_i2175_1_lut (.I0(baudrate[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n538));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2175_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2174_1_lut (.I0(baudrate[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n858));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2174_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2173_1_lut (.I0(baudrate[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2173_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2172_1_lut (.I0(baudrate[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n856));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2172_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2171_1_lut (.I0(baudrate[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1011));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2171_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2170_1_lut (.I0(baudrate[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1460));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2170_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2169_1_lut (.I0(baudrate[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1459));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2169_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2168_1_lut (.I0(baudrate[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2168_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2167_1_lut (.I0(baudrate[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1742));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2167_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2166_1_lut (.I0(baudrate[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1879));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2166_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2165_1_lut (.I0(baudrate[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2165_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2164_1_lut (.I0(baudrate[11]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2164_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2163_1_lut (.I0(baudrate[12]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2163_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2162_1_lut (.I0(baudrate[13]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2397));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2162_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2161_1_lut (.I0(baudrate[14]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2519));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2161_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2160_1_lut (.I0(baudrate[15]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2638));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2160_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2159_1_lut (.I0(baudrate[16]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2754));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2159_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2158_1_lut (.I0(baudrate[17]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2867));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2158_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2157_1_lut (.I0(baudrate[18]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2977));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2157_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2156_1_lut (.I0(baudrate[19]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2156_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2155_1_lut (.I0(baudrate[20]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2155_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i50442_3_lut_4_lut (.I0(n1558), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1559), .O(n66128));   // verilog/uart_rx.v(119[33:55])
    defparam i50442_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i2083_1_lut (.I0(baudrate[21]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2083_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2153_1_lut (.I0(baudrate[22]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2153_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1062_i34_3_lut_3_lut (.I0(n1558), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n34_adj_4723));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i7236_2_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n20919));   // verilog/uart_rx.v(119[33:55])
    defparam i7236_2_lut_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[24]), .I3(baudrate[31]), .O(n61676));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i46835_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[29]), .I3(baudrate[24]), .O(n62512));
    defparam i46835_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50605_3_lut_4_lut (.I0(n962), .I1(baudrate[1]), .I2(n48), 
            .I3(n25545), .O(n1115));
    defparam i50605_3_lut_4_lut.LUT_INIT = 16'haaa6;
    SB_LUT4 i5749_2_lut_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), 
            .I3(baudrate[1]), .O(n42));   // verilog/uart_rx.v(119[33:55])
    defparam i5749_2_lut_4_lut.LUT_INIT = 16'hb2bb;
    SB_LUT4 i5747_2_lut_3_lut (.I0(baudrate[2]), .I1(n962), .I2(baudrate[1]), 
            .I3(GND_net), .O(n11428));   // verilog/uart_rx.v(119[33:55])
    defparam i5747_2_lut_3_lut.LUT_INIT = 16'h4545;
    SB_LUT4 i50430_3_lut_4_lut (.I0(n1699), .I1(baudrate[4]), .I2(baudrate[3]), 
            .I3(n1700), .O(n66116));   // verilog/uart_rx.v(119[33:55])
    defparam i50430_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1157_i34_3_lut_3_lut (.I0(n1699), .I1(baudrate[4]), 
            .I2(baudrate[3]), .I3(GND_net), .O(n34_adj_4717));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i1_2_lut_4_lut_adj_1081 (.I0(n68282), .I1(baudrate[11]), .I2(n1831), 
            .I3(n60318), .O(n1977));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1081.LUT_INIT = 16'h7100;
    SB_LUT4 i53420_2_lut_4_lut (.I0(n68282), .I1(baudrate[11]), .I2(n1831), 
            .I3(n62546), .O(n294[12]));   // verilog/uart_rx.v(119[33:55])
    defparam i53420_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i1_2_lut_4_lut_adj_1082 (.I0(n68056), .I1(baudrate[14]), .I2(n2227), 
            .I3(n60320), .O(n2367));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1082.LUT_INIT = 16'h7100;
    SB_LUT4 i53429_2_lut_4_lut (.I0(n68056), .I1(baudrate[14]), .I2(n2227), 
            .I3(n62350), .O(n294[9]));   // verilog/uart_rx.v(119[33:55])
    defparam i53429_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i50682_2_lut (.I0(n56722), .I1(r_Rx_Data), .I2(GND_net), .I3(GND_net), 
            .O(n65372));
    defparam i50682_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_adj_1083 (.I0(n67714), .I1(baudrate[16]), .I2(n2476), 
            .I3(n60324), .O(n2612));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1083.LUT_INIT = 16'h7100;
    SB_LUT4 i53435_2_lut_4_lut (.I0(n67714), .I1(baudrate[16]), .I2(n2476), 
            .I3(n62318), .O(n294[7]));   // verilog/uart_rx.v(119[33:55])
    defparam i53435_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i53301_4_lut_4_lut (.I0(r_SM_Main_2__N_3446[1]), .I1(\r_SM_Main[1] ), 
            .I2(n6_adj_4724), .I3(n58912), .O(n58000));
    defparam i53301_4_lut_4_lut.LUT_INIT = 16'h0703;
    SB_LUT4 i50679_4_lut (.I0(n65372), .I1(n29), .I2(n23), .I3(\o_Rx_DV_N_3488[12] ), 
            .O(n65369));
    defparam i50679_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i50099_4_lut (.I0(n65369), .I1(r_SM_Main[0]), .I2(n27), .I3(\o_Rx_DV_N_3488[24] ), 
            .O(n65366));
    defparam i50099_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i53201_4_lut (.I0(\r_SM_Main[2] ), .I1(n65366), .I2(r_SM_Main_2__N_3446[1]), 
            .I3(\r_SM_Main[1] ), .O(n29148));
    defparam i53201_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i1_4_lut_adj_1084 (.I0(n56722), .I1(\r_SM_Main[1] ), .I2(r_Rx_Data), 
            .I3(r_SM_Main[0]), .O(n60400));
    defparam i1_4_lut_adj_1084.LUT_INIT = 16'h1000;
    SB_LUT4 i1_4_lut_adj_1085 (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3488[12] ), 
            .I3(n60400), .O(n60406));
    defparam i1_4_lut_adj_1085.LUT_INIT = 16'h0100;
    SB_LUT4 i52676_4_lut (.I0(\r_SM_Main[2] ), .I1(\o_Rx_DV_N_3488[24] ), 
            .I2(n27), .I3(n60406), .O(n27767));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i52676_4_lut.LUT_INIT = 16'h5455;
    SB_LUT4 i1_3_lut_4_lut_adj_1086 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n60696));
    defparam i1_3_lut_4_lut_adj_1086.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_3_lut_4_lut_adj_1087 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(\r_Bit_Index[0] ), .I3(n4), .O(n60680));
    defparam i1_3_lut_4_lut_adj_1087.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_4_lut_adj_1088 (.I0(n68186), .I1(baudrate[17]), .I2(n2596), 
            .I3(n60326), .O(n2730));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1088.LUT_INIT = 16'h7100;
    SB_LUT4 i53438_2_lut_4_lut (.I0(n68186), .I1(baudrate[17]), .I2(n2596), 
            .I3(n25619), .O(n294[6]));   // verilog/uart_rx.v(119[33:55])
    defparam i53438_2_lut_4_lut.LUT_INIT = 16'h0071;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (n2873, pwm_out, clk32MHz, pwm_setpoint, GND_net, n45, 
            n43, reset, \pwm_counter[22] , \pwm_counter[21] , VCC_net) /* synthesis syn_module_defined=1 */ ;
    input n2873;
    output pwm_out;
    input clk32MHz;
    input [23:0]pwm_setpoint;
    input GND_net;
    input n45;
    input n43;
    input reset;
    output \pwm_counter[22] ;
    output \pwm_counter[21] ;
    input VCC_net;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[16:24])
    
    wire pwm_out_N_577;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n65922, n6, n39, n41, n37, n29, n31, n23, n25, n35, 
        n11, n13, n15, n27, n33, n9, n17, n19, n21, n65876, 
        n65855, n12, n30, n66845, n66782, n67962, n67353, n68133, 
        n67371, n67372, n16, n24, n65761, n8, n65748, n67283, 
        n66555, n4, n67369, n67370, n65843, n10, n65839, n67964, 
        n66557, n68213, n68214, n68138, n65769, n67906, n66563, 
        n68119, n56471, n55503, n55531, n55551, n55579, n55607, 
        n55635, n55663, n55697, n55739, n55773, n55807, n55839, 
        n55867, n55899, n55935, n55963, n55995, n56055, n56179, 
        n56347, n56473, n56475, n56477, n50426, n48, n50425, n50424, 
        n50423, n50422, n50421, n50420, n50419, n50418, n50417, 
        n50416, n50415, n50414, n50413, n50412, n50411, n50410, 
        n50409, n50408, n50407, n50406, n50405, n50404, n60011, 
        n22, n15_adj_4450, n20, n24_adj_4451, n19_adj_4452;
    
    SB_DFFE pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .E(n2873), .D(pwm_out_N_577));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 i50236_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n65922));   // verilog/pwm.v(21[8:24])
    defparam i50236_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i50190_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n65876));
    defparam i50190_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i50169_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11), .O(n65855));
    defparam i50169_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51159_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n65922), 
            .O(n66845));
    defparam i51159_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i51096_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n66845), 
            .O(n66782));
    defparam i51096_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i52276_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n66782), 
            .O(n67962));
    defparam i52276_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51667_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n67962), 
            .O(n67353));
    defparam i51667_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i52447_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n67353), 
            .O(n68133));
    defparam i52447_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i51685_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n67371));   // verilog/pwm.v(21[8:24])
    defparam i51685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51686_3_lut (.I0(n67371), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n67372));   // verilog/pwm.v(21[8:24])
    defparam i51686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50075_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n65876), 
            .O(n65761));
    defparam i50075_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i51597_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n65748), 
            .O(n67283));   // verilog/pwm.v(21[8:24])
    defparam i51597_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50869_3_lut (.I0(n67372), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n66555));   // verilog/pwm.v(21[8:24])
    defparam i50869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_counter[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_setpoint[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i51683_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n67369));   // verilog/pwm.v(21[8:24])
    defparam i51683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i51684_3_lut (.I0(n67369), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n67370));   // verilog/pwm.v(21[8:24])
    defparam i51684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50157_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n65855), 
            .O(n65843));
    defparam i50157_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52278_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n65839), 
            .O(n67964));   // verilog/pwm.v(21[8:24])
    defparam i52278_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i50871_3_lut (.I0(n67370), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n66557));   // verilog/pwm.v(21[8:24])
    defparam i50871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52527_4_lut (.I0(n66557), .I1(n67964), .I2(n35), .I3(n65843), 
            .O(n68213));   // verilog/pwm.v(21[8:24])
    defparam i52527_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52528_3_lut (.I0(n68213), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n68214));   // verilog/pwm.v(21[8:24])
    defparam i52528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52452_3_lut (.I0(n68214), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n68138));   // verilog/pwm.v(21[8:24])
    defparam i52452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i50083_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n68133), 
            .O(n65769));
    defparam i50083_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i52220_4_lut (.I0(n66555), .I1(n67283), .I2(n45), .I3(n65761), 
            .O(n67906));   // verilog/pwm.v(21[8:24])
    defparam i52220_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i50877_3_lut (.I0(n68138), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n66563));   // verilog/pwm.v(21[8:24])
    defparam i50877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i52433_4_lut (.I0(n66563), .I1(n67906), .I2(n45), .I3(n65769), 
            .O(n68119));   // verilog/pwm.v(21[8:24])
    defparam i52433_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i52434_3_lut (.I0(n68119), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_577));   // verilog/pwm.v(21[8:24])
    defparam i52434_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFR pwm_counter_1939__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n56471), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n55503), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i22 (.Q(\pwm_counter[22] ), .C(clk32MHz), 
            .D(n55531), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i21 (.Q(\pwm_counter[21] ), .C(clk32MHz), 
            .D(n55551), .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n55579), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n55607), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n55635), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n55663), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n55697), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n55739), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n55773), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n55807), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n55839), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n55867), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n55899), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n55935), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n55963), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n55995), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n56055), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n56179), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n56347), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n56473), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n56475), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_1939__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n56477), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_LUT4 pwm_counter_1939_add_4_25_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n50426), .O(n55503)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 pwm_counter_1939_add_4_24_lut (.I0(n48), .I1(GND_net), .I2(\pwm_counter[22] ), 
            .I3(n50425), .O(n55531)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_24 (.CI(n50425), .I0(GND_net), .I1(\pwm_counter[22] ), 
            .CO(n50426));
    SB_LUT4 pwm_counter_1939_add_4_23_lut (.I0(n48), .I1(GND_net), .I2(\pwm_counter[21] ), 
            .I3(n50424), .O(n55551)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_23 (.CI(n50424), .I0(GND_net), .I1(\pwm_counter[21] ), 
            .CO(n50425));
    SB_LUT4 pwm_counter_1939_add_4_22_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n50423), .O(n55579)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_22 (.CI(n50423), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n50424));
    SB_LUT4 pwm_counter_1939_add_4_21_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n50422), .O(n55607)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_21 (.CI(n50422), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n50423));
    SB_LUT4 pwm_counter_1939_add_4_20_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n50421), .O(n55635)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_20 (.CI(n50421), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n50422));
    SB_LUT4 pwm_counter_1939_add_4_19_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n50420), .O(n55663)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_19 (.CI(n50420), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n50421));
    SB_LUT4 pwm_counter_1939_add_4_18_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n50419), .O(n55697)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_18 (.CI(n50419), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n50420));
    SB_LUT4 pwm_counter_1939_add_4_17_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n50418), .O(n55739)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_17 (.CI(n50418), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n50419));
    SB_LUT4 pwm_counter_1939_add_4_16_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n50417), .O(n55773)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_16 (.CI(n50417), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n50418));
    SB_LUT4 pwm_counter_1939_add_4_15_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n50416), .O(n55807)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_15 (.CI(n50416), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n50417));
    SB_LUT4 pwm_counter_1939_add_4_14_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n50415), .O(n55839)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_14 (.CI(n50415), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n50416));
    SB_LUT4 pwm_counter_1939_add_4_13_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n50414), .O(n55867)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_13 (.CI(n50414), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n50415));
    SB_LUT4 pwm_counter_1939_add_4_12_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n50413), .O(n55899)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_12 (.CI(n50413), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n50414));
    SB_LUT4 pwm_counter_1939_add_4_11_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n50412), .O(n55935)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_11 (.CI(n50412), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n50413));
    SB_LUT4 pwm_counter_1939_add_4_10_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n50411), .O(n55963)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_10 (.CI(n50411), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n50412));
    SB_LUT4 pwm_counter_1939_add_4_9_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n50410), .O(n55995)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_9 (.CI(n50410), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n50411));
    SB_LUT4 pwm_counter_1939_add_4_8_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n50409), .O(n56055)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_8 (.CI(n50409), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n50410));
    SB_LUT4 pwm_counter_1939_add_4_7_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n50408), .O(n56179)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_7 (.CI(n50408), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n50409));
    SB_LUT4 pwm_counter_1939_add_4_6_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n50407), .O(n56347)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_6 (.CI(n50407), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n50408));
    SB_LUT4 pwm_counter_1939_add_4_5_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n50406), .O(n56473)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_5 (.CI(n50406), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n50407));
    SB_LUT4 pwm_counter_1939_add_4_4_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n50405), .O(n56475)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_4 (.CI(n50405), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n50406));
    SB_LUT4 pwm_counter_1939_add_4_3_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n50404), .O(n56477)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_3 (.CI(n50404), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n50405));
    SB_LUT4 pwm_counter_1939_add_4_2_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n56471)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1939_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_1939_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n50404));
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50062_2_lut_4_lut (.I0(pwm_setpoint[21]), .I1(\pwm_counter[21] ), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n65748));
    defparam i50062_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(\pwm_counter[21] ), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i50153_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n65839));
    defparam i50153_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n60011));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_4_lut (.I0(pwm_counter[18]), .I1(pwm_counter[16]), .I2(pwm_counter[15]), 
            .I3(pwm_counter[19]), .O(n22));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n60011), .I1(pwm_counter[12]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n15_adj_4450));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i7_3_lut (.I0(pwm_counter[20]), .I1(\pwm_counter[22] ), .I2(pwm_counter[11]), 
            .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n15_adj_4450), .I1(n22), .I2(pwm_counter[13]), 
            .I3(\pwm_counter[21] ), .O(n24_adj_4451));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(pwm_counter[14]), .I1(pwm_counter[17]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4452));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(pwm_counter[23]), .I1(n19_adj_4452), .I2(n24_adj_4451), 
            .I3(n20), .O(n48));   // verilog/pwm.v(17[20:33])
    defparam i1_4_lut.LUT_INIT = 16'haaab;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (\state[1] , \state[0] , GND_net, n6, n5, n6_adj_8, 
            n42774, state_7__N_4317, n42779, \data[15] , n27706, clk16MHz, 
            n11, n9, clk_out, n29648, CS_c, n29646, \current[0] , 
            n29643, n29628, \data[12] , n29627, \data[11] , n29626, 
            \data[10] , n29625, \data[9] , n29624, \data[8] , n29617, 
            \data[7] , n29612, \data[6] , n29608, \data[5] , n29607, 
            \data[4] , n29606, \data[3] , n29605, \data[2] , n29604, 
            \data[1] , VCC_net, n30506, \data[0] , n30394, \current[1] , 
            n30393, \current[2] , n30392, \current[3] , n30391, \current[4] , 
            n30390, \current[5] , n30389, \current[6] , n30388, \current[7] , 
            n30387, \current[8] , n30386, \current[9] , n30385, \current[10] , 
            n30383, \current[11] , \current[15] , CS_CLK_c, n6_adj_9, 
            n5_adj_10, n15, n25532, n25571, n25523, n25519, n4, 
            n25527) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \state[1] ;
    output \state[0] ;
    input GND_net;
    output n6;
    output n5;
    output n6_adj_8;
    output n42774;
    output state_7__N_4317;
    output n42779;
    output \data[15] ;
    output n27706;
    input clk16MHz;
    output n11;
    input n9;
    output clk_out;
    input n29648;
    output CS_c;
    input n29646;
    output \current[0] ;
    input n29643;
    input n29628;
    output \data[12] ;
    input n29627;
    output \data[11] ;
    input n29626;
    output \data[10] ;
    input n29625;
    output \data[9] ;
    input n29624;
    output \data[8] ;
    input n29617;
    output \data[7] ;
    input n29612;
    output \data[6] ;
    input n29608;
    output \data[5] ;
    input n29607;
    output \data[4] ;
    input n29606;
    output \data[3] ;
    input n29605;
    output \data[2] ;
    input n29604;
    output \data[1] ;
    input VCC_net;
    input n30506;
    output \data[0] ;
    input n30394;
    output \current[1] ;
    input n30393;
    output \current[2] ;
    input n30392;
    output \current[3] ;
    input n30391;
    output \current[4] ;
    input n30390;
    output \current[5] ;
    input n30389;
    output \current[6] ;
    input n30388;
    output \current[7] ;
    input n30387;
    output \current[8] ;
    input n30386;
    output \current[9] ;
    input n30385;
    output \current[10] ;
    input n30383;
    output \current[11] ;
    output \current[15] ;
    output CS_CLK_c;
    output n6_adj_9;
    output n5_adj_10;
    output n15;
    output n25532;
    output n25571;
    output n25523;
    output n25519;
    output n4;
    output n25527;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n27762, n65364, n22566;
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    
    wire n12180, n27989, n28887, clk_slow_N_4230, n29159;
    wire [2:0]n17;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire n50539, n50538;
    wire [11:0]n53;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire n50537, n50536, delay_counter_15__N_4312, clk_slow_N_4231, 
        n50535, n50534, n50533, n50532, n50531, n50530, n50529, 
        n50528, n50527;
    wire [7:0]n37;
    
    wire n22568, n22570, n22572, n50433, n50432, n50431, n50430, 
        n65363, n50429, n2, n65358, n50428, n65308, n50427;
    wire [1:0]n1859;
    
    wire n42838, n8, n12, n10, n6_adj_4449;
    
    SB_LUT4 i14023_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n27762));
    defparam i14023_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i8825_3_lut (.I0(\state[0] ), .I1(n65364), .I2(\state[1] ), 
            .I3(GND_net), .O(n22566));   // verilog/tli4970.v(55[24:39])
    defparam i8825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_333_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/tli4970.v(54[9:26])
    defparam equal_333_i6_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_324_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(54[9:26])
    defparam equal_324_i5_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_328_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_8));   // verilog/tli4970.v(54[9:26])
    defparam equal_328_i6_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i28872_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n42774));
    defparam i28872_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_7__I_0_77_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(state_7__N_4317));   // verilog/tli4970.v(53[7:17])
    defparam state_7__I_0_77_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i28877_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(GND_net), 
            .I3(GND_net), .O(n42779));
    defparam i28877_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i52684_3_lut (.I0(\data[15] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n27706));
    defparam i52684_3_lut.LUT_INIT = 16'h4040;
    SB_DFFNESR state_i1 (.Q(\state[1] ), .C(clk_slow), .E(n27989), .D(n12180), 
            .R(n28887));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFF clk_slow_63 (.Q(clk_slow), .C(clk16MHz), .D(clk_slow_N_4230));   // verilog/tli4970.v(13[10] 19[6])
    SB_LUT4 i15152_2_lut_2_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n29159));   // verilog/tli4970.v(55[24:39])
    defparam i15152_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 equal_264_i11_2_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(bit_counter[2]), .I3(bit_counter[3]), .O(n11));   // verilog/tli4970.v(56[12:26])
    defparam equal_264_i11_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFN clk_out_67 (.Q(clk_out), .C(clk_slow), .D(n9));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN slave_select_66 (.Q(CS_c), .C(clk_slow), .D(n29648));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i1 (.Q(\current[0] ), .C(clk_slow), .D(n29646));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n29643));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n29628));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n29627));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n29626));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n29625));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n29624));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n29617));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n29612));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n29608));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n29607));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n29606));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n29605));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n29604));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 counter_1948_1949_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n50539), .O(n17[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1948_1949_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFNE bit_counter_1940__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n27762), 
            .D(n22566));   // verilog/tli4970.v(55[24:39])
    SB_LUT4 counter_1948_1949_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n50538), .O(n17[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1948_1949_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1948_1949_add_4_3 (.CI(n50538), .I0(GND_net), .I1(counter[1]), 
            .CO(n50539));
    SB_LUT4 counter_1948_1949_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n17[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_1948_1949_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_1948_1949_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n50538));
    SB_LUT4 delay_counter_1946_1947_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n50537), .O(n53[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_1946_1947_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n50536), .O(n53[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_DFFNSR delay_counter_1946_1947__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n53[0]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_1948_1949__i1 (.Q(counter[0]), .C(clk16MHz), .D(n17[0]), 
            .R(clk_slow_N_4231));   // verilog/tli4970.v(14[16:27])
    SB_CARRY delay_counter_1946_1947_add_4_12 (.CI(n50536), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n50537));
    SB_LUT4 delay_counter_1946_1947_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n50535), .O(n53[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_11 (.CI(n50535), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n50536));
    SB_LUT4 delay_counter_1946_1947_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n50534), .O(n53[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_10 (.CI(n50534), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n50535));
    SB_LUT4 delay_counter_1946_1947_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n50533), .O(n53[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_9 (.CI(n50533), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n50534));
    SB_LUT4 delay_counter_1946_1947_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n50532), .O(n53[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_8 (.CI(n50532), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n50533));
    SB_LUT4 delay_counter_1946_1947_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n50531), .O(n53[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_7 (.CI(n50531), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n50532));
    SB_LUT4 delay_counter_1946_1947_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n50530), .O(n53[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_6 (.CI(n50530), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n50531));
    SB_LUT4 delay_counter_1946_1947_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n50529), .O(n53[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_5 (.CI(n50529), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n50530));
    SB_LUT4 delay_counter_1946_1947_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n50528), .O(n53[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_4 (.CI(n50528), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n50529));
    SB_LUT4 delay_counter_1946_1947_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n50527), .O(n53[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_3 (.CI(n50527), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n50528));
    SB_LUT4 delay_counter_1946_1947_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n53[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1946_1947_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1946_1947_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n50527));
    SB_DFFSR counter_1948_1949__i3 (.Q(counter[2]), .C(clk16MHz), .D(n17[2]), 
            .R(clk_slow_N_4231));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_1948_1949__i2 (.Q(counter[1]), .C(clk16MHz), .D(n17[1]), 
            .R(clk_slow_N_4231));   // verilog/tli4970.v(14[16:27])
    SB_DFFNSR delay_counter_1946_1947__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n53[11]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n53[10]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n53[9]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n53[8]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n53[7]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n53[6]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n53[5]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n53[4]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n53[3]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n53[2]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_1946_1947__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n53[1]), .R(delay_counter_15__N_4312));   // verilog/tli4970.v(40[24:39])
    SB_DFFNESR bit_counter_1940__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n27762), 
            .D(n37[4]), .R(n29159));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1940__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n27762), 
            .D(n37[5]), .R(n29159));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1940__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n27762), 
            .D(n37[6]), .R(n29159));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_1940__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n27762), 
            .D(n37[7]), .R(n29159));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_1940__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n27762), 
            .D(n22568));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_1940__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n27762), 
            .D(n22570));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_1940__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n27762), 
            .D(n22572));   // verilog/tli4970.v(55[24:39])
    SB_LUT4 bit_counter_1940_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n50433), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1940_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_1940_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n50432), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1940_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1940_add_4_8 (.CI(n50432), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n50433));
    SB_LUT4 bit_counter_1940_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n50431), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1940_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1940_add_4_7 (.CI(n50431), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n50432));
    SB_LUT4 bit_counter_1940_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n50430), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1940_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_1940_add_4_6 (.CI(n50430), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n50431));
    SB_LUT4 bit_counter_1940_add_4_5_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n50429), .O(n65363)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1940_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_1940_add_4_5 (.CI(n50429), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n50430));
    SB_LUT4 bit_counter_1940_add_4_4_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n50428), .O(n65358)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1940_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_1940_add_4_4 (.CI(n50428), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n50429));
    SB_LUT4 bit_counter_1940_add_4_3_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n50427), .O(n65308)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1940_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_1940_add_4_3 (.CI(n50427), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n50428));
    SB_LUT4 bit_counter_1940_add_4_2_lut (.I0(n2), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n65364)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_1940_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_1940_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n50427));
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n30506));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i2 (.Q(\current[1] ), .C(clk_slow), .D(n30394));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i3 (.Q(\current[2] ), .C(clk_slow), .D(n30393));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i4 (.Q(\current[3] ), .C(clk_slow), .D(n30392));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i5 (.Q(\current[4] ), .C(clk_slow), .D(n30391));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i6 (.Q(\current[5] ), .C(clk_slow), .D(n30390));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i7 (.Q(\current[6] ), .C(clk_slow), .D(n30389));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i8 (.Q(\current[7] ), .C(clk_slow), .D(n30388));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i9 (.Q(\current[8] ), .C(clk_slow), .D(n30387));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i10 (.Q(\current[9] ), .C(clk_slow), .D(n30386));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i11 (.Q(\current[10] ), .C(clk_slow), .D(n30385));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i12 (.Q(\current[11] ), .C(clk_slow), .D(n30383));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE current__i13 (.Q(\current[15] ), .C(clk_slow), .E(n27706), 
            .D(n1859[0]));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNESS state_i0 (.Q(\state[0] ), .C(clk_slow), .E(n27989), .D(n42838), 
            .S(n28887));   // verilog/tli4970.v(35[10] 68[6])
    SB_LUT4 i2121_1_lut (.I0(\data[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1859[0]));
    defparam i2121_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2065_3_lut (.I0(counter[0]), .I1(counter[2]), .I2(counter[1]), 
            .I3(GND_net), .O(clk_slow_N_4231));
    defparam i2065_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 clk_slow_I_0_72_2_lut (.I0(clk_slow), .I1(clk_slow_N_4231), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4230));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_72_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 equal_335_i6_2_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_9));   // verilog/tli4970.v(54[9:26])
    defparam equal_335_i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_326_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_10));   // verilog/tli4970.v(54[9:26])
    defparam equal_326_i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_3_lut (.I0(delay_counter[1]), .I1(delay_counter[2]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2066_4_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(n8), 
            .I3(delay_counter[0]), .O(n12));
    defparam i2066_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i4_4_lut (.I0(delay_counter[11]), .I1(delay_counter[7]), .I2(delay_counter[8]), 
            .I3(delay_counter[9]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut (.I0(delay_counter[10]), .I1(n10), .I2(n12), .I3(delay_counter[6]), 
            .O(delay_counter_15__N_4312));
    defparam i5_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 i1_2_lut (.I0(bit_counter[5]), .I1(bit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4449));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_964 (.I0(bit_counter[6]), .I1(bit_counter[7]), 
            .I2(n11), .I3(n6_adj_4449), .O(n15));   // verilog/tli4970.v(56[12:26])
    defparam i4_4_lut_adj_964.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_2033_i2_3_lut (.I0(n15), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n12180));
    defparam mux_2033_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut (.I0(n15), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(delay_counter_15__N_4312), .O(n27989));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hffdc;
    SB_LUT4 i14879_2_lut_4_lut (.I0(n15), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(delay_counter_15__N_4312), .O(n28887));
    defparam i14879_2_lut_4_lut.LUT_INIT = 16'h2300;
    SB_LUT4 i2397_1_lut (.I0(\state[0] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2));
    defparam i2397_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52702_2_lut (.I0(n15), .I1(\state[0] ), .I2(GND_net), .I3(GND_net), 
            .O(n42838));
    defparam i52702_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i8831_3_lut (.I0(\state[0] ), .I1(n65308), .I2(\state[1] ), 
            .I3(GND_net), .O(n22572));   // verilog/tli4970.v(55[24:39])
    defparam i8831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8829_3_lut (.I0(\state[0] ), .I1(n65358), .I2(\state[1] ), 
            .I3(GND_net), .O(n22570));   // verilog/tli4970.v(55[24:39])
    defparam i8829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8827_3_lut (.I0(\state[0] ), .I1(n65363), .I2(\state[1] ), 
            .I3(GND_net), .O(n22568));   // verilog/tli4970.v(55[24:39])
    defparam i8827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_965 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n25532));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_965.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_4_lut_adj_966 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[0]), 
            .I3(bit_counter[1]), .O(n25571));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_966.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_4_lut_adj_967 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n25523));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_967.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_3_lut_4_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n25519));   // verilog/tli4970.v(43[5] 67[12])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_4_lut_adj_968 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n4));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_968.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_4_lut_adj_969 (.I0(\state[0] ), .I1(\state[1] ), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n25527));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_4_lut_adj_969.LUT_INIT = 16'hfffb;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (\state[1] , \state[0] , n3, \state[2] , GND_net, enable_slow_N_4211, 
            ready_prev, n42699, n57012, n25516, data, ID, clk16MHz, 
            n5773, n25404, n27997, n29647, rw, n56425, data_ready, 
            n55999, n56203, baudrate, n30406, n30405, n30404, n30403, 
            n30402, n30401, n30400, n30399, \state_7__N_3916[0] , 
            \state[0]_adj_4 , n4, scl_enable, n6428, \state_7__N_4108[0] , 
            scl, sda_enable, sda_out, n29654, \saved_addr[0] , VCC_net, 
            n30492, n8, n30216, n30215, n30214, n30213, n30212, 
            n30211, n30210, n4_adj_5, n4_adj_6, n65481, n42804, 
            n10, n25540, n25535, \state_7__N_4124[3] , n10_adj_7) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \state[1] ;
    output \state[0] ;
    output n3;
    output \state[2] ;
    input GND_net;
    output enable_slow_N_4211;
    output ready_prev;
    output n42699;
    output n57012;
    output n25516;
    output [7:0]data;
    output [7:0]ID;
    input clk16MHz;
    output [0:0]n5773;
    output n25404;
    output n27997;
    input n29647;
    output rw;
    input n56425;
    output data_ready;
    input n55999;
    input n56203;
    output [31:0]baudrate;
    input n30406;
    input n30405;
    input n30404;
    input n30403;
    input n30402;
    input n30401;
    input n30400;
    input n30399;
    input \state_7__N_3916[0] ;
    output \state[0]_adj_4 ;
    output n4;
    output scl_enable;
    output n6428;
    output \state_7__N_4108[0] ;
    output scl;
    output sda_enable;
    output sda_out;
    input n29654;
    output \saved_addr[0] ;
    input VCC_net;
    input n30492;
    input n8;
    input n30216;
    input n30215;
    input n30214;
    input n30213;
    input n30212;
    input n30211;
    input n30210;
    output n4_adj_5;
    output n4_adj_6;
    output n65481;
    output n42804;
    output n10;
    output n25540;
    output n25535;
    input \state_7__N_4124[3] ;
    output n10_adj_7;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n47429;
    wire [15:0]delay_counter_15__N_3954;
    wire [15:0]delay_counter;   // verilog/eeprom.v(28[12:25])
    wire [15:0]n5113;
    
    wire n49420, n49421, n6681, n49419, n47410, n6, n50883;
    wire [2:0]byte_counter;   // verilog/eeprom.v(30[11:23])
    
    wire n15, n30432, n30433, n49418, enable, n30434, n30435, 
        n49417, n49416, n30436, n51818, n28, n26, n27, n30437, 
        n25, n30438, n29642, n27697;
    wire [2:0]n17;
    
    wire n27769, n29156, n30431, n30430, n30429, n30428, n30427, 
        n30426, n30425, n30424, n30423, n30422, n30421, n30419, 
        n56333, n56337, n56331, n56335, n30414, n30413, n30412, 
        n30411, n30410, n30409, n30408, n30407;
    wire [7:0]state_7__N_3883;
    
    wire n59887, n4_c, n62324;
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    wire n65490, n6687, n6686, n6685, n6684, n6683, n47407, n49430, 
        n49429, n49428, n49427, n49426, n49425, n49424, n49423, 
        n49422, n4_adj_4442, n47437;
    
    SB_LUT4 i1_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(n3), .I3(\state[2] ), 
            .O(n47429));
    defparam i1_4_lut.LUT_INIT = 16'h0144;
    SB_LUT4 add_1103_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n5113[11]), 
            .I3(n49420), .O(delay_counter_15__N_3954[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_7 (.CI(n49420), .I0(delay_counter[5]), .I1(n5113[11]), 
            .CO(n49421));
    SB_LUT4 add_1103_6_lut (.I0(n47410), .I1(delay_counter[4]), .I2(n5113[11]), 
            .I3(n49419), .O(n6681)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i28797_2_lut (.I0(enable_slow_N_4211), .I1(ready_prev), .I2(GND_net), 
            .I3(GND_net), .O(n42699));
    defparam i28797_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut (.I0(ready_prev), .I1(n57012), .I2(\state[2] ), .I3(n6), 
            .O(n50883));
    defparam i4_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_adj_954 (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n25516));   // verilog/eeprom.v(38[3] 80[10])
    defparam i1_2_lut_adj_954.LUT_INIT = 16'heeee;
    SB_LUT4 i16424_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[7]), 
            .I3(ID[7]), .O(n30432));
    defparam i16424_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16425_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[6]), 
            .I3(ID[6]), .O(n30433));
    defparam i16425_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_1103_6 (.CI(n49419), .I0(delay_counter[4]), .I1(n5113[11]), 
            .CO(n49420));
    SB_LUT4 add_1103_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n5113[11]), 
            .I3(n49418), .O(delay_counter_15__N_3954[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF ready_prev_59 (.Q(ready_prev), .C(clk16MHz), .D(enable_slow_N_4211));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFSR enable_58 (.Q(enable), .C(clk16MHz), .D(n5773[0]), .R(\state[2] ));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i16426_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[5]), 
            .I3(ID[5]), .O(n30434));
    defparam i16426_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_1103_5 (.CI(n49418), .I0(delay_counter[3]), .I1(n5113[11]), 
            .CO(n49419));
    SB_LUT4 i16427_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[4]), 
            .I3(ID[4]), .O(n30435));
    defparam i16427_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_1103_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n5113[11]), 
            .I3(n49417), .O(delay_counter_15__N_3954[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_4 (.CI(n49417), .I0(delay_counter[2]), .I1(n5113[11]), 
            .CO(n49418));
    SB_LUT4 add_1103_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n5113[11]), 
            .I3(n49416), .O(delay_counter_15__N_3954[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_3 (.CI(n49416), .I0(delay_counter[1]), .I1(n5113[11]), 
            .CO(n49417));
    SB_LUT4 add_1103_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n5113[11]), 
            .I3(GND_net), .O(delay_counter_15__N_3954[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n5113[11]), 
            .CO(n49416));
    SB_LUT4 i16428_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[3]), 
            .I3(ID[3]), .O(n30436));
    defparam i16428_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut (.I0(enable_slow_N_4211), .I1(ready_prev), .I2(byte_counter[0]), 
            .I3(GND_net), .O(n51818));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hd2d2;
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(55[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[2]), .I2(delay_counter[7]), 
            .I3(delay_counter[5]), .O(n26));   // verilog/eeprom.v(55[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n27));   // verilog/eeprom.v(55[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16429_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[2]), 
            .I3(ID[2]), .O(n30437));
    defparam i16429_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(55[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n25404));   // verilog/eeprom.v(55[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i52704_2_lut (.I0(n25404), .I1(enable_slow_N_4211), .I2(GND_net), 
            .I3(GND_net), .O(n5113[11]));   // verilog/eeprom.v(59[18] 61[12])
    defparam i52704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16430_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[1]), 
            .I3(ID[1]), .O(n30438));
    defparam i16430_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15634_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[0]), 
            .I3(ID[0]), .O(n29642));
    defparam i15634_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut (.I0(byte_counter[1]), .I1(n50883), .I2(byte_counter[2]), 
            .I3(byte_counter[0]), .O(n27997));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i25_4_lut_4_lut (.I0(\state[1] ), .I1(n3), .I2(\state[0] ), 
            .I3(\state[2] ), .O(n27697));
    defparam i25_4_lut_4_lut.LUT_INIT = 16'h015a;
    SB_LUT4 i1_2_lut_3_lut_adj_955 (.I0(byte_counter[1]), .I1(n50883), .I2(byte_counter[2]), 
            .I3(GND_net), .O(n15));
    defparam i1_2_lut_3_lut_adj_955.LUT_INIT = 16'hfbfb;
    SB_DFF rw_64 (.Q(rw), .C(clk16MHz), .D(n29647));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF data_ready_61 (.Q(data_ready), .C(clk16MHz), .D(n56425));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i1 (.Q(ID[0]), .C(clk16MHz), .D(n29642));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF state_i2 (.Q(\state[2] ), .C(clk16MHz), .D(n55999));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR byte_counter_1945__i1 (.Q(byte_counter[1]), .C(clk16MHz), 
            .E(n27769), .D(n17[1]), .R(n29156));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_1945__i2 (.Q(byte_counter[2]), .C(clk16MHz), 
            .E(n27769), .D(n17[2]), .R(n29156));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_1945__i0 (.Q(byte_counter[0]), .C(clk16MHz), 
            .E(n27769), .D(n51818), .R(n29156));   // verilog/eeprom.v(68[25:39])
    SB_DFF state_i0 (.Q(\state[0] ), .C(clk16MHz), .D(n56203));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i2 (.Q(ID[1]), .C(clk16MHz), .D(n30438));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i3 (.Q(ID[2]), .C(clk16MHz), .D(n30437));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i4 (.Q(ID[3]), .C(clk16MHz), .D(n30436));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i5 (.Q(ID[4]), .C(clk16MHz), .D(n30435));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i6 (.Q(ID[5]), .C(clk16MHz), .D(n30434));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i7 (.Q(ID[6]), .C(clk16MHz), .D(n30433));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i8 (.Q(ID[7]), .C(clk16MHz), .D(n30432));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i9 (.Q(baudrate[0]), .C(clk16MHz), .D(n30431));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i10 (.Q(baudrate[1]), .C(clk16MHz), .D(n30430));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i11 (.Q(baudrate[2]), .C(clk16MHz), .D(n30429));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i12 (.Q(baudrate[3]), .C(clk16MHz), .D(n30428));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i13 (.Q(baudrate[4]), .C(clk16MHz), .D(n30427));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i14 (.Q(baudrate[5]), .C(clk16MHz), .D(n30426));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i15 (.Q(baudrate[6]), .C(clk16MHz), .D(n30425));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i16 (.Q(baudrate[7]), .C(clk16MHz), .D(n30424));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i17 (.Q(baudrate[8]), .C(clk16MHz), .D(n30423));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i18 (.Q(baudrate[9]), .C(clk16MHz), .D(n30422));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i19 (.Q(baudrate[10]), .C(clk16MHz), .D(n30421));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i20 (.Q(baudrate[11]), .C(clk16MHz), .D(n30419));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i21 (.Q(baudrate[12]), .C(clk16MHz), .D(n56333));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i22 (.Q(baudrate[13]), .C(clk16MHz), .D(n56337));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i23 (.Q(baudrate[14]), .C(clk16MHz), .D(n56331));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i24 (.Q(baudrate[15]), .C(clk16MHz), .D(n56335));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i25 (.Q(baudrate[16]), .C(clk16MHz), .D(n30414));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i26 (.Q(baudrate[17]), .C(clk16MHz), .D(n30413));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i27 (.Q(baudrate[18]), .C(clk16MHz), .D(n30412));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i28 (.Q(baudrate[19]), .C(clk16MHz), .D(n30411));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i29 (.Q(baudrate[20]), .C(clk16MHz), .D(n30410));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i30 (.Q(baudrate[21]), .C(clk16MHz), .D(n30409));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i31 (.Q(baudrate[22]), .C(clk16MHz), .D(n30408));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i32 (.Q(baudrate[23]), .C(clk16MHz), .D(n30407));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i33 (.Q(baudrate[24]), .C(clk16MHz), .D(n30406));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i34 (.Q(baudrate[25]), .C(clk16MHz), .D(n30405));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i35 (.Q(baudrate[26]), .C(clk16MHz), .D(n30404));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i36 (.Q(baudrate[27]), .C(clk16MHz), .D(n30403));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i37 (.Q(baudrate[28]), .C(clk16MHz), .D(n30402));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i38 (.Q(baudrate[29]), .C(clk16MHz), .D(n30401));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i39 (.Q(baudrate[30]), .C(clk16MHz), .D(n30400));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i40 (.Q(baudrate[31]), .C(clk16MHz), .D(n30399));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk16MHz), .E(n59887), .D(state_7__N_3883[1]));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i1_4_lut_adj_956 (.I0(\state[2] ), .I1(\state[1] ), .I2(\state_7__N_3916[0] ), 
            .I3(\state[0] ), .O(n4_c));
    defparam i1_4_lut_adj_956.LUT_INIT = 16'hbbba;
    SB_LUT4 i50674_4_lut (.I0(n62324), .I1(n25404), .I2(\state[1] ), .I3(state[3]), 
            .O(n65490));
    defparam i50674_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i2_4_lut (.I0(n65490), .I1(n4_c), .I2(n42699), .I3(\state[0] ), 
            .O(n59887));
    defparam i2_4_lut.LUT_INIT = 16'hcfee;
    SB_LUT4 i1_4_lut_adj_957 (.I0(n3), .I1(\state[0] ), .I2(\state[2] ), 
            .I3(\state[1] ), .O(state_7__N_3883[1]));
    defparam i1_4_lut_adj_957.LUT_INIT = 16'hf31c;
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(clk16MHz), 
            .E(n27697), .D(delay_counter_15__N_3954[15]), .R(n47429));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(clk16MHz), 
            .E(n27697), .D(delay_counter_15__N_3954[14]), .R(n47429));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(clk16MHz), 
            .E(n27697), .D(delay_counter_15__N_3954[13]), .R(n47429));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(clk16MHz), 
            .E(n27697), .D(delay_counter_15__N_3954[12]), .R(n47429));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(clk16MHz), 
            .E(n27697), .D(delay_counter_15__N_3954[11]), .R(n47429));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(clk16MHz), 
            .E(n27697), .D(n6687), .S(n47429));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n27697), 
            .D(n6686), .S(n47429));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n27697), 
            .D(n6685), .S(n47429));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n27697), 
            .D(n6684), .S(n47429));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n27697), 
            .D(n6683), .S(n47429));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n27697), 
            .D(delay_counter_15__N_3954[5]), .R(n47429));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n27697), 
            .D(n6681), .S(n47407));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n27697), 
            .D(delay_counter_15__N_3954[3]), .R(n47429));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n27697), 
            .D(delay_counter_15__N_3954[2]), .R(n47429));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n27697), 
            .D(delay_counter_15__N_3954[1]), .R(n47429));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n27697), 
            .D(delay_counter_15__N_3954[0]), .R(n47429));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 add_1103_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n5113[11]), 
            .I3(n49430), .O(delay_counter_15__N_3954[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1103_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n5113[11]), 
            .I3(n49429), .O(delay_counter_15__N_3954[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_16 (.CI(n49429), .I0(delay_counter[14]), .I1(n5113[11]), 
            .CO(n49430));
    SB_LUT4 add_1103_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n5113[11]), 
            .I3(n49428), .O(delay_counter_15__N_3954[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_15 (.CI(n49428), .I0(delay_counter[13]), .I1(n5113[11]), 
            .CO(n49429));
    SB_LUT4 add_1103_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n5113[11]), 
            .I3(n49427), .O(delay_counter_15__N_3954[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_14 (.CI(n49427), .I0(delay_counter[12]), .I1(n5113[11]), 
            .CO(n49428));
    SB_LUT4 add_1103_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n5113[11]), 
            .I3(n49426), .O(delay_counter_15__N_3954[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1103_13 (.CI(n49426), .I0(delay_counter[11]), .I1(n5113[11]), 
            .CO(n49427));
    SB_LUT4 add_1103_12_lut (.I0(n47410), .I1(delay_counter[10]), .I2(n5113[11]), 
            .I3(n49425), .O(n6687)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1103_12 (.CI(n49425), .I0(delay_counter[10]), .I1(n5113[11]), 
            .CO(n49426));
    SB_LUT4 add_1103_11_lut (.I0(n47410), .I1(delay_counter[9]), .I2(n5113[11]), 
            .I3(n49424), .O(n6686)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1103_11 (.CI(n49424), .I0(delay_counter[9]), .I1(n5113[11]), 
            .CO(n49425));
    SB_LUT4 add_1103_10_lut (.I0(n47410), .I1(delay_counter[8]), .I2(n5113[11]), 
            .I3(n49423), .O(n6685)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1103_10 (.CI(n49423), .I0(delay_counter[8]), .I1(n5113[11]), 
            .CO(n49424));
    SB_LUT4 add_1103_9_lut (.I0(n47410), .I1(delay_counter[7]), .I2(n5113[11]), 
            .I3(n49422), .O(n6684)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1103_9 (.CI(n49422), .I0(delay_counter[7]), .I1(n5113[11]), 
            .CO(n49423));
    SB_LUT4 add_1103_8_lut (.I0(n47410), .I1(delay_counter[6]), .I2(n5113[11]), 
            .I3(n49421), .O(n6683)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1103_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1103_8 (.CI(n49421), .I0(delay_counter[6]), .I1(n5113[11]), 
            .CO(n49422));
    SB_LUT4 i46653_2_lut_3_lut (.I0(state[1]), .I1(state[2]), .I2(\state[0]_adj_4 ), 
            .I3(GND_net), .O(n62324));   // verilog/eeprom.v(55[12:28])
    defparam i46653_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(state[1]), .I1(state[2]), .I2(state[3]), 
            .I3(\state[0]_adj_4 ), .O(n4));   // verilog/eeprom.v(55[12:28])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_4_lut (.I0(state[1]), .I1(state[2]), .I2(\state[0]_adj_4 ), 
            .I3(state[3]), .O(n4_adj_4442));   // verilog/eeprom.v(55[12:28])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hffc1;
    SB_LUT4 i2_3_lut_4_lut_adj_958 (.I0(\state[1] ), .I1(\state_7__N_3916[0] ), 
            .I2(\state[0] ), .I3(\state[2] ), .O(n29156));   // verilog/eeprom.v(68[25:39])
    defparam i2_3_lut_4_lut_adj_958.LUT_INIT = 16'h0004;
    SB_LUT4 i1_4_lut_4_lut_adj_959 (.I0(\state[1] ), .I1(\state_7__N_3916[0] ), 
            .I2(\state[0] ), .I3(\state[2] ), .O(n27769));   // verilog/eeprom.v(68[25:39])
    defparam i1_4_lut_4_lut_adj_959.LUT_INIT = 16'h00a4;
    SB_LUT4 i35150_3_lut_4_lut (.I0(n42699), .I1(byte_counter[0]), .I2(byte_counter[1]), 
            .I3(byte_counter[2]), .O(n17[2]));   // verilog/eeprom.v(68[25:39])
    defparam i35150_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 i35143_2_lut_3_lut_4_lut (.I0(enable_slow_N_4211), .I1(ready_prev), 
            .I2(byte_counter[0]), .I3(byte_counter[1]), .O(n17[1]));   // verilog/eeprom.v(68[25:39])
    defparam i35143_2_lut_3_lut_4_lut.LUT_INIT = 16'hdf20;
    SB_LUT4 mux_1450_Mux_0_i3_4_lut (.I0(\state[0] ), .I1(enable_slow_N_4211), 
            .I2(\state[1] ), .I3(n25404), .O(n5773[0]));   // verilog/eeprom.v(38[3] 80[10])
    defparam mux_1450_Mux_0_i3_4_lut.LUT_INIT = 16'h0a4a;
    SB_LUT4 i2_3_lut (.I0(byte_counter[2]), .I1(n50883), .I2(byte_counter[1]), 
            .I3(GND_net), .O(n47437));
    defparam i2_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1_3_lut (.I0(byte_counter[0]), .I1(byte_counter[2]), .I2(byte_counter[1]), 
            .I3(GND_net), .O(n3));   // verilog/eeprom.v(30[11:23])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13_2_lut (.I0(\state[2] ), .I1(n3), .I2(GND_net), .I3(GND_net), 
            .O(n47410));
    defparam i13_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i16423_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[0]), 
            .I3(baudrate[0]), .O(n30431));   // verilog/eeprom.v(68[25:39])
    defparam i16423_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16416_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[7]), 
            .I3(baudrate[7]), .O(n30424));   // verilog/eeprom.v(68[25:39])
    defparam i16416_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16417_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[6]), 
            .I3(baudrate[6]), .O(n30425));   // verilog/eeprom.v(68[25:39])
    defparam i16417_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16418_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[5]), 
            .I3(baudrate[5]), .O(n30426));   // verilog/eeprom.v(68[25:39])
    defparam i16418_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16419_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[4]), 
            .I3(baudrate[4]), .O(n30427));   // verilog/eeprom.v(68[25:39])
    defparam i16419_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16420_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[3]), 
            .I3(baudrate[3]), .O(n30428));   // verilog/eeprom.v(68[25:39])
    defparam i16420_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16421_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[2]), 
            .I3(baudrate[2]), .O(n30429));   // verilog/eeprom.v(68[25:39])
    defparam i16421_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16422_3_lut_4_lut (.I0(byte_counter[0]), .I1(n15), .I2(data[1]), 
            .I3(baudrate[1]), .O(n30430));   // verilog/eeprom.v(68[25:39])
    defparam i16422_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16411_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47437), .I2(data[3]), 
            .I3(baudrate[11]), .O(n30419));   // verilog/eeprom.v(68[25:39])
    defparam i16411_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i11_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47437), .I2(data[7]), 
            .I3(baudrate[15]), .O(n56335));   // verilog/eeprom.v(68[25:39])
    defparam i11_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i11_3_lut_4_lut_adj_960 (.I0(byte_counter[0]), .I1(n47437), 
            .I2(data[6]), .I3(baudrate[14]), .O(n56331));   // verilog/eeprom.v(68[25:39])
    defparam i11_3_lut_4_lut_adj_960.LUT_INIT = 16'hfb40;
    SB_LUT4 i11_3_lut_4_lut_adj_961 (.I0(byte_counter[0]), .I1(n47437), 
            .I2(data[4]), .I3(baudrate[12]), .O(n56333));   // verilog/eeprom.v(68[25:39])
    defparam i11_3_lut_4_lut_adj_961.LUT_INIT = 16'hfb40;
    SB_LUT4 i16414_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47437), .I2(data[1]), 
            .I3(baudrate[9]), .O(n30422));   // verilog/eeprom.v(68[25:39])
    defparam i16414_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16413_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47437), .I2(data[2]), 
            .I3(baudrate[10]), .O(n30421));   // verilog/eeprom.v(68[25:39])
    defparam i16413_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16415_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47437), .I2(data[0]), 
            .I3(baudrate[8]), .O(n30423));   // verilog/eeprom.v(68[25:39])
    defparam i16415_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i11_3_lut_4_lut_adj_962 (.I0(byte_counter[0]), .I1(n47437), 
            .I2(data[5]), .I3(baudrate[13]), .O(n56337));   // verilog/eeprom.v(68[25:39])
    defparam i11_3_lut_4_lut_adj_962.LUT_INIT = 16'hfb40;
    SB_LUT4 i16406_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47437), .I2(data[0]), 
            .I3(baudrate[16]), .O(n30414));   // verilog/eeprom.v(68[25:39])
    defparam i16406_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16399_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47437), .I2(data[7]), 
            .I3(baudrate[23]), .O(n30407));   // verilog/eeprom.v(68[25:39])
    defparam i16399_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16400_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47437), .I2(data[6]), 
            .I3(baudrate[22]), .O(n30408));   // verilog/eeprom.v(68[25:39])
    defparam i16400_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16401_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47437), .I2(data[5]), 
            .I3(baudrate[21]), .O(n30409));   // verilog/eeprom.v(68[25:39])
    defparam i16401_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16402_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47437), .I2(data[4]), 
            .I3(baudrate[20]), .O(n30410));   // verilog/eeprom.v(68[25:39])
    defparam i16402_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_4_lut_adj_963 (.I0(\state[0]_adj_4 ), .I1(state[3]), 
            .I2(state[2]), .I3(state[1]), .O(n57012));   // verilog/eeprom.v(55[12:28])
    defparam i2_3_lut_4_lut_adj_963.LUT_INIT = 16'hfffe;
    SB_LUT4 i16403_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47437), .I2(data[3]), 
            .I3(baudrate[19]), .O(n30411));   // verilog/eeprom.v(68[25:39])
    defparam i16403_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16404_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47437), .I2(data[2]), 
            .I3(baudrate[18]), .O(n30412));   // verilog/eeprom.v(68[25:39])
    defparam i16404_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16405_3_lut_4_lut (.I0(byte_counter[0]), .I1(n47437), .I2(data[1]), 
            .I3(baudrate[17]), .O(n30413));   // verilog/eeprom.v(68[25:39])
    defparam i16405_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i33521_4_lut_4_lut (.I0(\state[1] ), .I1(n3), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n47407));
    defparam i33521_4_lut_4_lut.LUT_INIT = 16'h0510;
    i2c_controller i2c (.\state[0] (\state[0]_adj_4 ), .\state[1] (state[1]), 
            .\state[2] (state[2]), .\state[3] (state[3]), .clk16MHz(clk16MHz), 
            .scl_enable(scl_enable), .GND_net(GND_net), .n6428(n6428), 
            .\state_7__N_4108[0] (\state_7__N_4108[0] ), .enable_slow_N_4211(enable_slow_N_4211), 
            .scl(scl), .sda_enable(sda_enable), .sda_out(sda_out), .n29654(n29654), 
            .\saved_addr[0] (\saved_addr[0] ), .VCC_net(VCC_net), .n30492(n30492), 
            .data({data}), .n8(n8), .n30216(n30216), .n30215(n30215), 
            .n30214(n30214), .n30213(n30213), .n30212(n30212), .n30211(n30211), 
            .n30210(n30210), .n4(n4_adj_5), .n4_adj_1(n4_adj_6), .n65481(n65481), 
            .n42804(n42804), .n10(n10), .n25540(n25540), .n25535(n25535), 
            .enable(enable), .\state_7__N_4124[3] (\state_7__N_4124[3] ), 
            .n10_adj_2(n10_adj_7), .n4_adj_3(n4_adj_4442)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(83[16] 97[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (\state[0] , \state[1] , \state[2] , \state[3] , 
            clk16MHz, scl_enable, GND_net, n6428, \state_7__N_4108[0] , 
            enable_slow_N_4211, scl, sda_enable, sda_out, n29654, 
            \saved_addr[0] , VCC_net, n30492, data, n8, n30216, 
            n30215, n30214, n30213, n30212, n30211, n30210, n4, 
            n4_adj_1, n65481, n42804, n10, n25540, n25535, enable, 
            \state_7__N_4124[3] , n10_adj_2, n4_adj_3) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output \state[0] ;
    output \state[1] ;
    output \state[2] ;
    output \state[3] ;
    input clk16MHz;
    output scl_enable;
    input GND_net;
    output n6428;
    output \state_7__N_4108[0] ;
    output enable_slow_N_4211;
    output scl;
    output sda_enable;
    output sda_out;
    input n29654;
    output \saved_addr[0] ;
    input VCC_net;
    input n30492;
    output [7:0]data;
    input n8;
    input n30216;
    input n30215;
    input n30214;
    input n30213;
    input n30212;
    input n30211;
    input n30210;
    output n4;
    output n4_adj_1;
    output n65481;
    output n42804;
    output n10;
    output n25540;
    output n25535;
    input enable;
    input \state_7__N_4124[3] ;
    output n10_adj_2;
    input n4_adj_3;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n15, i2c_clk_N_4197, scl_enable_N_4198, n27952, n28897, n42750, 
        n58968, n58866, enable_slow_N_4210, n27757, sda_out_adj_4428;
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n50559, n50558, n50557, n50556, n50555, n29139;
    wire [7:0]n119;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n5, n43435, n42949, n43239, n60107, n27752, n56275, n59097, 
        n27750, n49437, n49436, n49435, n49434, n49433, n49432, 
        n49431, n10_c, n11, n11_adj_4430, n11_adj_4431, n27619, 
        n4_adj_4432, n9, n11_adj_4434;
    wire [1:0]n6491;
    
    wire n6758, n28, n68345, n57925, n6421, n11_adj_4435, n12, 
        n65492;
    
    SB_LUT4 equal_272_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n15));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_272_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_DFF i2c_clk_122 (.Q(i2c_clk), .C(clk16MHz), .D(i2c_clk_N_4197));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_124 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4198));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_LUT4 i14889_2_lut_4_lut (.I0(n27952), .I1(\state[3] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n28897));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14889_2_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i29439_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n42750));
    defparam i29439_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i53263_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[1] ), 
            .I3(n6428), .O(n58968));
    defparam i53263_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n58866));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h1110;
    SB_DFFE enable_slow_121 (.Q(\state_7__N_4108[0] ), .C(clk16MHz), .E(n27757), 
            .D(enable_slow_N_4210));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_LUT4 i52697_2_lut (.I0(\state_7__N_4108[0] ), .I1(enable_slow_N_4211), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4210));   // verilog/i2c_controller.v(62[6:32])
    defparam i52697_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i28817_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i28817_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2431_2_lut (.I0(sda_out_adj_4428), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2431_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter2_1954_1955_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n50559), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1954_1955_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_1954_1955_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n50558), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1954_1955_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1954_1955_add_4_6 (.CI(n50558), .I0(GND_net), .I1(counter2[4]), 
            .CO(n50559));
    SB_LUT4 counter2_1954_1955_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n50557), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1954_1955_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1954_1955_add_4_5 (.CI(n50557), .I0(GND_net), .I1(counter2[3]), 
            .CO(n50558));
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n29654));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 counter2_1954_1955_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n50556), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1954_1955_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1954_1955_add_4_4 (.CI(n50556), .I0(GND_net), .I1(counter2[2]), 
            .CO(n50557));
    SB_LUT4 counter2_1954_1955_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n50555), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1954_1955_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1954_1955_add_4_3 (.CI(n50555), .I0(GND_net), .I1(counter2[1]), 
            .CO(n50556));
    SB_LUT4 counter2_1954_1955_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1954_1955_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1954_1955_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n50555));
    SB_DFFSR counter2_1954_1955__i6 (.Q(counter2[5]), .C(clk16MHz), .D(n29[5]), 
            .R(n29139));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1954_1955__i5 (.Q(counter2[4]), .C(clk16MHz), .D(n29[4]), 
            .R(n29139));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1954_1955__i4 (.Q(counter2[3]), .C(clk16MHz), .D(n29[3]), 
            .R(n29139));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1954_1955__i3 (.Q(counter2[2]), .C(clk16MHz), .D(n29[2]), 
            .R(n29139));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1954_1955__i2 (.Q(counter2[1]), .C(clk16MHz), .D(n29[1]), 
            .R(n29139));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n27952), .D(n119[1]), 
            .S(n28897));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n27952), .D(n119[2]), 
            .S(n28897));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n27952), .D(n119[3]), 
            .R(n28897));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n27952), .D(n119[4]), 
            .R(n28897));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n27952), .D(n119[5]), 
            .R(n28897));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n27952), .D(n119[6]), 
            .R(n28897));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n27952), .D(n119[7]), 
            .R(n28897));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n6428), .D(n5), 
            .S(n43435));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n6428), .D(n42949), 
            .S(n43239));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n6428), .D(n60107), 
            .S(n58968));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_1954_1955__i1 (.Q(counter2[0]), .C(clk16MHz), .D(n29[0]), 
            .R(n29139));   // verilog/i2c_controller.v(69[20:35])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n30492));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n30216));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n30215));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n30214));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n30213));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n30212));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n30211));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n30210));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFNESS write_enable_132 (.Q(sda_enable), .C(i2c_clk), .E(n27752), 
            .D(n58866), .S(n56275));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFNESS sda_out_133 (.Q(sda_out_adj_4428), .C(i2c_clk), .E(n27750), 
            .D(n59097), .S(n56275));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n27952), .D(n119[0]), 
            .S(n28897));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n49437), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n49436), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n49436), .I0(counter[6]), .I1(VCC_net), 
            .CO(n49437));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n49435), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n49435), .I0(counter[5]), .I1(VCC_net), 
            .CO(n49436));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n49434), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n49434), .I0(counter[4]), .I1(VCC_net), 
            .CO(n49435));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n49433), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n49433), .I0(counter[3]), .I1(VCC_net), 
            .CO(n49434));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n49432), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n49432), .I0(counter[2]), .I1(VCC_net), 
            .CO(n49433));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n49431), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n49431), .I0(counter[1]), .I1(VCC_net), 
            .CO(n49432));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n49431));
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_c));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_c), .I2(counter2[0]), 
            .I3(GND_net), .O(n29139));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut (.I0(i2c_clk), .I1(n29139), .I2(GND_net), .I3(GND_net), 
            .O(i2c_clk_N_4197));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[3] ), .I1(\state[2] ), 
            .I2(\state[0] ), .I3(\state[1] ), .O(n11));
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 equal_351_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_351_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_349_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_1));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_349_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i50365_3_lut_4_lut (.I0(n11), .I1(n11_adj_4430), .I2(enable_slow_N_4211), 
            .I3(\state_7__N_4108[0] ), .O(n65481));
    defparam i50365_3_lut_4_lut.LUT_INIT = 16'h0888;
    SB_LUT4 i53273_3_lut_4_lut (.I0(n11), .I1(n11_adj_4430), .I2(n15), 
            .I3(n6428), .O(n43435));
    defparam i53273_3_lut_4_lut.LUT_INIT = 16'h7f00;
    SB_LUT4 i28902_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n42804));
    defparam i28902_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_7__I_0_140_i11_2_lut_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4431));
    defparam state_7__I_0_140_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n27619));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 state_7__I_0_142_i11_2_lut_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(\state[1] ), .I3(\state[0] ), .O(n11_adj_4430));   // verilog/i2c_controller.v(77[47:62])
    defparam state_7__I_0_142_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_3_lut_4_lut_adj_945 (.I0(\state[2] ), .I1(\state[3] ), .I2(n4_adj_4432), 
            .I3(n9), .O(n60107));   // verilog/i2c_controller.v(77[47:62])
    defparam i2_3_lut_4_lut_adj_945.LUT_INIT = 16'hf0f4;
    SB_LUT4 i1_2_lut_3_lut (.I0(n9), .I1(n10), .I2(counter[0]), .I3(GND_net), 
            .O(n25540));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_946 (.I0(n9), .I1(n10), .I2(counter[0]), 
            .I3(GND_net), .O(n25535));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_946.LUT_INIT = 16'hefef;
    SB_LUT4 i53271_3_lut_4_lut (.I0(n9), .I1(n10), .I2(n11_adj_4430), 
            .I3(n6428), .O(n43239));   // verilog/i2c_controller.v(151[5:14])
    defparam i53271_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_LUT4 i28860_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(n15), .O(scl_enable_N_4198));   // verilog/i2c_controller.v(44[32:47])
    defparam i28860_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i52711_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(enable_slow_N_4211));   // verilog/i2c_controller.v(44[32:47])
    defparam i52711_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 equal_1517_i11_2_lut_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4434));
    defparam equal_1517_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i2_3_lut_4_lut_adj_947 (.I0(\state[3] ), .I1(\state[2] ), .I2(n6491[1]), 
            .I3(\state[1] ), .O(n59097));
    defparam i2_3_lut_4_lut_adj_947.LUT_INIT = 16'h1000;
    SB_LUT4 i1_2_lut_3_lut_adj_948 (.I0(\state[3] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n6758));
    defparam i1_2_lut_3_lut_adj_948.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_949 (.I0(enable), .I1(\state_7__N_4108[0] ), 
            .I2(enable_slow_N_4211), .I3(GND_net), .O(n27757));
    defparam i1_2_lut_3_lut_adj_949.LUT_INIT = 16'haeae;
    SB_LUT4 i1_4_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\state[2] ), .O(n28));
    defparam i1_4_lut.LUT_INIT = 16'h5110;
    SB_LUT4 i52659_2_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n68345));
    defparam i52659_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_950 (.I0(n11_adj_4434), .I1(n68345), .I2(n28), 
            .I3(n57925), .O(n27750));
    defparam i1_4_lut_adj_950.LUT_INIT = 16'ha0a8;
    SB_LUT4 mux_1730_Mux_1_i7_4_lut (.I0(counter[1]), .I1(counter[0]), .I2(counter[2]), 
            .I3(\saved_addr[0] ), .O(n6491[1]));   // verilog/i2c_controller.v(201[28:35])
    defparam mux_1730_Mux_1_i7_4_lut.LUT_INIT = 16'hc1c0;
    SB_LUT4 i29525_2_lut (.I0(\state[2] ), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n57925));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i29525_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(n11_adj_4434), .I1(n57925), .I2(\state[3] ), 
            .I3(\state[1] ), .O(n56275));
    defparam i3_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i1_4_lut_adj_951 (.I0(n11_adj_4434), .I1(\state[1] ), .I2(\state[3] ), 
            .I3(n57925), .O(n27752));
    defparam i1_4_lut_adj_951.LUT_INIT = 16'h0a22;
    SB_LUT4 i1_4_lut_adj_952 (.I0(\state_7__N_4124[3] ), .I1(n11_adj_4431), 
            .I2(n11_adj_4434), .I3(enable), .O(n4_adj_4432));
    defparam i1_4_lut_adj_952.LUT_INIT = 16'h2a2f;
    SB_LUT4 i53177_2_lut (.I0(\state_7__N_4124[3] ), .I1(n11_adj_4431), 
            .I2(GND_net), .I3(GND_net), .O(n42949));
    defparam i53177_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 state_7__I_0_141_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(130[5:15])
    defparam state_7__I_0_141_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 state_7__I_0_144_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_144_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i52682_4_lut (.I0(n27619), .I1(n6421), .I2(n11), .I3(n42750), 
            .O(n6428));
    defparam i52682_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i1_4_lut_adj_953 (.I0(n11_adj_4435), .I1(n11_adj_4431), .I2(\state_7__N_4124[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_953.LUT_INIT = 16'h5755;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_2));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10_adj_2), 
            .O(n6421));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 state_7__I_0_145_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4435));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_145_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i50739_2_lut (.I0(n15), .I1(\state_7__N_4124[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n65492));
    defparam i50739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14_4_lut (.I0(n6421), .I1(n65492), .I2(n6758), .I3(n4_adj_3), 
            .O(n27952));
    defparam i14_4_lut.LUT_INIT = 16'h303a;
    
endmodule
