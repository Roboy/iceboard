-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Feb 17 2020 11:47:55

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    TX : out std_logic;
    SDA : in std_logic;
    SCL : in std_logic;
    RX : in std_logic;
    NEOPXL : out std_logic;
    LED : out std_logic;
    INLC : out std_logic;
    INLB : out std_logic;
    INLA : out std_logic;
    INHC : out std_logic;
    INHB : out std_logic;
    INHA : out std_logic;
    HALL3 : in std_logic;
    HALL2 : in std_logic;
    HALL1 : in std_logic;
    FAULT_N : in std_logic;
    ENCODER1_B : in std_logic;
    ENCODER1_A : in std_logic;
    ENCODER0_B : in std_logic;
    ENCODER0_A : in std_logic;
    DE : out std_logic;
    CS_MISO : in std_logic;
    CS_CLK : out std_logic;
    CS : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__56752\ : std_logic;
signal \N__56751\ : std_logic;
signal \N__56750\ : std_logic;
signal \N__56743\ : std_logic;
signal \N__56742\ : std_logic;
signal \N__56741\ : std_logic;
signal \N__56734\ : std_logic;
signal \N__56733\ : std_logic;
signal \N__56732\ : std_logic;
signal \N__56725\ : std_logic;
signal \N__56724\ : std_logic;
signal \N__56723\ : std_logic;
signal \N__56716\ : std_logic;
signal \N__56715\ : std_logic;
signal \N__56714\ : std_logic;
signal \N__56707\ : std_logic;
signal \N__56706\ : std_logic;
signal \N__56705\ : std_logic;
signal \N__56698\ : std_logic;
signal \N__56697\ : std_logic;
signal \N__56696\ : std_logic;
signal \N__56689\ : std_logic;
signal \N__56688\ : std_logic;
signal \N__56687\ : std_logic;
signal \N__56680\ : std_logic;
signal \N__56679\ : std_logic;
signal \N__56678\ : std_logic;
signal \N__56671\ : std_logic;
signal \N__56670\ : std_logic;
signal \N__56669\ : std_logic;
signal \N__56662\ : std_logic;
signal \N__56661\ : std_logic;
signal \N__56660\ : std_logic;
signal \N__56653\ : std_logic;
signal \N__56652\ : std_logic;
signal \N__56651\ : std_logic;
signal \N__56644\ : std_logic;
signal \N__56643\ : std_logic;
signal \N__56642\ : std_logic;
signal \N__56635\ : std_logic;
signal \N__56634\ : std_logic;
signal \N__56633\ : std_logic;
signal \N__56626\ : std_logic;
signal \N__56625\ : std_logic;
signal \N__56624\ : std_logic;
signal \N__56617\ : std_logic;
signal \N__56616\ : std_logic;
signal \N__56615\ : std_logic;
signal \N__56608\ : std_logic;
signal \N__56607\ : std_logic;
signal \N__56606\ : std_logic;
signal \N__56599\ : std_logic;
signal \N__56598\ : std_logic;
signal \N__56597\ : std_logic;
signal \N__56590\ : std_logic;
signal \N__56589\ : std_logic;
signal \N__56588\ : std_logic;
signal \N__56571\ : std_logic;
signal \N__56568\ : std_logic;
signal \N__56565\ : std_logic;
signal \N__56562\ : std_logic;
signal \N__56559\ : std_logic;
signal \N__56556\ : std_logic;
signal \N__56553\ : std_logic;
signal \N__56550\ : std_logic;
signal \N__56547\ : std_logic;
signal \N__56544\ : std_logic;
signal \N__56541\ : std_logic;
signal \N__56538\ : std_logic;
signal \N__56535\ : std_logic;
signal \N__56532\ : std_logic;
signal \N__56529\ : std_logic;
signal \N__56526\ : std_logic;
signal \N__56523\ : std_logic;
signal \N__56522\ : std_logic;
signal \N__56521\ : std_logic;
signal \N__56520\ : std_logic;
signal \N__56519\ : std_logic;
signal \N__56518\ : std_logic;
signal \N__56517\ : std_logic;
signal \N__56516\ : std_logic;
signal \N__56515\ : std_logic;
signal \N__56514\ : std_logic;
signal \N__56513\ : std_logic;
signal \N__56512\ : std_logic;
signal \N__56511\ : std_logic;
signal \N__56510\ : std_logic;
signal \N__56509\ : std_logic;
signal \N__56508\ : std_logic;
signal \N__56497\ : std_logic;
signal \N__56494\ : std_logic;
signal \N__56491\ : std_logic;
signal \N__56488\ : std_logic;
signal \N__56485\ : std_logic;
signal \N__56476\ : std_logic;
signal \N__56469\ : std_logic;
signal \N__56466\ : std_logic;
signal \N__56461\ : std_logic;
signal \N__56450\ : std_logic;
signal \N__56447\ : std_logic;
signal \N__56442\ : std_logic;
signal \N__56441\ : std_logic;
signal \N__56440\ : std_logic;
signal \N__56439\ : std_logic;
signal \N__56436\ : std_logic;
signal \N__56433\ : std_logic;
signal \N__56432\ : std_logic;
signal \N__56431\ : std_logic;
signal \N__56428\ : std_logic;
signal \N__56425\ : std_logic;
signal \N__56416\ : std_logic;
signal \N__56413\ : std_logic;
signal \N__56410\ : std_logic;
signal \N__56407\ : std_logic;
signal \N__56406\ : std_logic;
signal \N__56405\ : std_logic;
signal \N__56404\ : std_logic;
signal \N__56403\ : std_logic;
signal \N__56398\ : std_logic;
signal \N__56395\ : std_logic;
signal \N__56392\ : std_logic;
signal \N__56389\ : std_logic;
signal \N__56384\ : std_logic;
signal \N__56381\ : std_logic;
signal \N__56378\ : std_logic;
signal \N__56373\ : std_logic;
signal \N__56364\ : std_logic;
signal \N__56363\ : std_logic;
signal \N__56360\ : std_logic;
signal \N__56359\ : std_logic;
signal \N__56356\ : std_logic;
signal \N__56355\ : std_logic;
signal \N__56354\ : std_logic;
signal \N__56353\ : std_logic;
signal \N__56344\ : std_logic;
signal \N__56341\ : std_logic;
signal \N__56338\ : std_logic;
signal \N__56333\ : std_logic;
signal \N__56328\ : std_logic;
signal \N__56327\ : std_logic;
signal \N__56326\ : std_logic;
signal \N__56325\ : std_logic;
signal \N__56324\ : std_logic;
signal \N__56323\ : std_logic;
signal \N__56322\ : std_logic;
signal \N__56321\ : std_logic;
signal \N__56320\ : std_logic;
signal \N__56319\ : std_logic;
signal \N__56316\ : std_logic;
signal \N__56307\ : std_logic;
signal \N__56304\ : std_logic;
signal \N__56297\ : std_logic;
signal \N__56294\ : std_logic;
signal \N__56287\ : std_logic;
signal \N__56284\ : std_logic;
signal \N__56277\ : std_logic;
signal \N__56274\ : std_logic;
signal \N__56271\ : std_logic;
signal \N__56268\ : std_logic;
signal \N__56265\ : std_logic;
signal \N__56262\ : std_logic;
signal \N__56261\ : std_logic;
signal \N__56260\ : std_logic;
signal \N__56259\ : std_logic;
signal \N__56258\ : std_logic;
signal \N__56257\ : std_logic;
signal \N__56256\ : std_logic;
signal \N__56255\ : std_logic;
signal \N__56254\ : std_logic;
signal \N__56253\ : std_logic;
signal \N__56252\ : std_logic;
signal \N__56251\ : std_logic;
signal \N__56250\ : std_logic;
signal \N__56249\ : std_logic;
signal \N__56248\ : std_logic;
signal \N__56247\ : std_logic;
signal \N__56246\ : std_logic;
signal \N__56245\ : std_logic;
signal \N__56244\ : std_logic;
signal \N__56243\ : std_logic;
signal \N__56242\ : std_logic;
signal \N__56241\ : std_logic;
signal \N__56240\ : std_logic;
signal \N__56239\ : std_logic;
signal \N__56238\ : std_logic;
signal \N__56237\ : std_logic;
signal \N__56236\ : std_logic;
signal \N__56235\ : std_logic;
signal \N__56234\ : std_logic;
signal \N__56233\ : std_logic;
signal \N__56232\ : std_logic;
signal \N__56231\ : std_logic;
signal \N__56230\ : std_logic;
signal \N__56229\ : std_logic;
signal \N__56228\ : std_logic;
signal \N__56227\ : std_logic;
signal \N__56226\ : std_logic;
signal \N__56225\ : std_logic;
signal \N__56224\ : std_logic;
signal \N__56223\ : std_logic;
signal \N__56222\ : std_logic;
signal \N__56221\ : std_logic;
signal \N__56220\ : std_logic;
signal \N__56219\ : std_logic;
signal \N__56218\ : std_logic;
signal \N__56217\ : std_logic;
signal \N__56216\ : std_logic;
signal \N__56215\ : std_logic;
signal \N__56214\ : std_logic;
signal \N__56213\ : std_logic;
signal \N__56212\ : std_logic;
signal \N__56211\ : std_logic;
signal \N__56210\ : std_logic;
signal \N__56209\ : std_logic;
signal \N__56208\ : std_logic;
signal \N__56207\ : std_logic;
signal \N__56206\ : std_logic;
signal \N__56205\ : std_logic;
signal \N__56204\ : std_logic;
signal \N__56203\ : std_logic;
signal \N__56202\ : std_logic;
signal \N__56201\ : std_logic;
signal \N__56200\ : std_logic;
signal \N__56199\ : std_logic;
signal \N__56070\ : std_logic;
signal \N__56067\ : std_logic;
signal \N__56064\ : std_logic;
signal \N__56063\ : std_logic;
signal \N__56060\ : std_logic;
signal \N__56057\ : std_logic;
signal \N__56056\ : std_logic;
signal \N__56053\ : std_logic;
signal \N__56050\ : std_logic;
signal \N__56047\ : std_logic;
signal \N__56040\ : std_logic;
signal \N__56037\ : std_logic;
signal \N__56034\ : std_logic;
signal \N__56031\ : std_logic;
signal \N__56030\ : std_logic;
signal \N__56029\ : std_logic;
signal \N__56026\ : std_logic;
signal \N__56023\ : std_logic;
signal \N__56020\ : std_logic;
signal \N__56015\ : std_logic;
signal \N__56012\ : std_logic;
signal \N__56009\ : std_logic;
signal \N__56006\ : std_logic;
signal \N__56001\ : std_logic;
signal \N__55998\ : std_logic;
signal \N__55995\ : std_logic;
signal \N__55994\ : std_logic;
signal \N__55993\ : std_logic;
signal \N__55990\ : std_logic;
signal \N__55985\ : std_logic;
signal \N__55980\ : std_logic;
signal \N__55977\ : std_logic;
signal \N__55974\ : std_logic;
signal \N__55971\ : std_logic;
signal \N__55968\ : std_logic;
signal \N__55965\ : std_logic;
signal \N__55962\ : std_logic;
signal \N__55959\ : std_logic;
signal \N__55956\ : std_logic;
signal \N__55955\ : std_logic;
signal \N__55952\ : std_logic;
signal \N__55949\ : std_logic;
signal \N__55946\ : std_logic;
signal \N__55941\ : std_logic;
signal \N__55938\ : std_logic;
signal \N__55937\ : std_logic;
signal \N__55934\ : std_logic;
signal \N__55931\ : std_logic;
signal \N__55928\ : std_logic;
signal \N__55923\ : std_logic;
signal \N__55920\ : std_logic;
signal \N__55917\ : std_logic;
signal \N__55916\ : std_logic;
signal \N__55913\ : std_logic;
signal \N__55912\ : std_logic;
signal \N__55911\ : std_logic;
signal \N__55908\ : std_logic;
signal \N__55905\ : std_logic;
signal \N__55902\ : std_logic;
signal \N__55899\ : std_logic;
signal \N__55898\ : std_logic;
signal \N__55897\ : std_logic;
signal \N__55894\ : std_logic;
signal \N__55891\ : std_logic;
signal \N__55888\ : std_logic;
signal \N__55885\ : std_logic;
signal \N__55882\ : std_logic;
signal \N__55881\ : std_logic;
signal \N__55878\ : std_logic;
signal \N__55875\ : std_logic;
signal \N__55872\ : std_logic;
signal \N__55869\ : std_logic;
signal \N__55866\ : std_logic;
signal \N__55863\ : std_logic;
signal \N__55860\ : std_logic;
signal \N__55857\ : std_logic;
signal \N__55850\ : std_logic;
signal \N__55841\ : std_logic;
signal \N__55836\ : std_logic;
signal \N__55835\ : std_logic;
signal \N__55832\ : std_logic;
signal \N__55829\ : std_logic;
signal \N__55826\ : std_logic;
signal \N__55821\ : std_logic;
signal \N__55820\ : std_logic;
signal \N__55817\ : std_logic;
signal \N__55814\ : std_logic;
signal \N__55811\ : std_logic;
signal \N__55806\ : std_logic;
signal \N__55805\ : std_logic;
signal \N__55802\ : std_logic;
signal \N__55799\ : std_logic;
signal \N__55796\ : std_logic;
signal \N__55791\ : std_logic;
signal \N__55790\ : std_logic;
signal \N__55787\ : std_logic;
signal \N__55784\ : std_logic;
signal \N__55779\ : std_logic;
signal \N__55776\ : std_logic;
signal \N__55775\ : std_logic;
signal \N__55772\ : std_logic;
signal \N__55769\ : std_logic;
signal \N__55766\ : std_logic;
signal \N__55761\ : std_logic;
signal \N__55760\ : std_logic;
signal \N__55757\ : std_logic;
signal \N__55754\ : std_logic;
signal \N__55751\ : std_logic;
signal \N__55748\ : std_logic;
signal \N__55745\ : std_logic;
signal \N__55742\ : std_logic;
signal \N__55739\ : std_logic;
signal \N__55734\ : std_logic;
signal \N__55731\ : std_logic;
signal \N__55728\ : std_logic;
signal \N__55725\ : std_logic;
signal \N__55722\ : std_logic;
signal \N__55719\ : std_logic;
signal \N__55716\ : std_logic;
signal \N__55715\ : std_logic;
signal \N__55712\ : std_logic;
signal \N__55709\ : std_logic;
signal \N__55706\ : std_logic;
signal \N__55701\ : std_logic;
signal \N__55698\ : std_logic;
signal \N__55695\ : std_logic;
signal \N__55694\ : std_logic;
signal \N__55691\ : std_logic;
signal \N__55688\ : std_logic;
signal \N__55685\ : std_logic;
signal \N__55680\ : std_logic;
signal \N__55677\ : std_logic;
signal \N__55674\ : std_logic;
signal \N__55671\ : std_logic;
signal \N__55668\ : std_logic;
signal \N__55667\ : std_logic;
signal \N__55664\ : std_logic;
signal \N__55661\ : std_logic;
signal \N__55658\ : std_logic;
signal \N__55653\ : std_logic;
signal \N__55650\ : std_logic;
signal \N__55647\ : std_logic;
signal \N__55646\ : std_logic;
signal \N__55643\ : std_logic;
signal \N__55640\ : std_logic;
signal \N__55637\ : std_logic;
signal \N__55632\ : std_logic;
signal \N__55629\ : std_logic;
signal \N__55626\ : std_logic;
signal \N__55625\ : std_logic;
signal \N__55622\ : std_logic;
signal \N__55619\ : std_logic;
signal \N__55616\ : std_logic;
signal \N__55611\ : std_logic;
signal \N__55608\ : std_logic;
signal \N__55605\ : std_logic;
signal \N__55602\ : std_logic;
signal \N__55599\ : std_logic;
signal \N__55596\ : std_logic;
signal \N__55593\ : std_logic;
signal \N__55592\ : std_logic;
signal \N__55591\ : std_logic;
signal \N__55588\ : std_logic;
signal \N__55583\ : std_logic;
signal \N__55580\ : std_logic;
signal \N__55575\ : std_logic;
signal \N__55572\ : std_logic;
signal \N__55569\ : std_logic;
signal \N__55566\ : std_logic;
signal \N__55563\ : std_logic;
signal \N__55562\ : std_logic;
signal \N__55559\ : std_logic;
signal \N__55558\ : std_logic;
signal \N__55557\ : std_logic;
signal \N__55556\ : std_logic;
signal \N__55555\ : std_logic;
signal \N__55554\ : std_logic;
signal \N__55553\ : std_logic;
signal \N__55552\ : std_logic;
signal \N__55551\ : std_logic;
signal \N__55550\ : std_logic;
signal \N__55549\ : std_logic;
signal \N__55548\ : std_logic;
signal \N__55547\ : std_logic;
signal \N__55546\ : std_logic;
signal \N__55545\ : std_logic;
signal \N__55544\ : std_logic;
signal \N__55543\ : std_logic;
signal \N__55542\ : std_logic;
signal \N__55541\ : std_logic;
signal \N__55540\ : std_logic;
signal \N__55539\ : std_logic;
signal \N__55538\ : std_logic;
signal \N__55537\ : std_logic;
signal \N__55536\ : std_logic;
signal \N__55535\ : std_logic;
signal \N__55534\ : std_logic;
signal \N__55533\ : std_logic;
signal \N__55532\ : std_logic;
signal \N__55531\ : std_logic;
signal \N__55530\ : std_logic;
signal \N__55529\ : std_logic;
signal \N__55528\ : std_logic;
signal \N__55527\ : std_logic;
signal \N__55526\ : std_logic;
signal \N__55521\ : std_logic;
signal \N__55518\ : std_logic;
signal \N__55515\ : std_logic;
signal \N__55512\ : std_logic;
signal \N__55509\ : std_logic;
signal \N__55506\ : std_logic;
signal \N__55503\ : std_logic;
signal \N__55500\ : std_logic;
signal \N__55497\ : std_logic;
signal \N__55496\ : std_logic;
signal \N__55495\ : std_logic;
signal \N__55494\ : std_logic;
signal \N__55493\ : std_logic;
signal \N__55492\ : std_logic;
signal \N__55491\ : std_logic;
signal \N__55490\ : std_logic;
signal \N__55487\ : std_logic;
signal \N__55486\ : std_logic;
signal \N__55485\ : std_logic;
signal \N__55482\ : std_logic;
signal \N__55479\ : std_logic;
signal \N__55478\ : std_logic;
signal \N__55477\ : std_logic;
signal \N__55476\ : std_logic;
signal \N__55473\ : std_logic;
signal \N__55470\ : std_logic;
signal \N__55463\ : std_logic;
signal \N__55456\ : std_logic;
signal \N__55455\ : std_logic;
signal \N__55454\ : std_logic;
signal \N__55453\ : std_logic;
signal \N__55450\ : std_logic;
signal \N__55447\ : std_logic;
signal \N__55446\ : std_logic;
signal \N__55445\ : std_logic;
signal \N__55444\ : std_logic;
signal \N__55441\ : std_logic;
signal \N__55438\ : std_logic;
signal \N__55437\ : std_logic;
signal \N__55436\ : std_logic;
signal \N__55435\ : std_logic;
signal \N__55434\ : std_logic;
signal \N__55433\ : std_logic;
signal \N__55432\ : std_logic;
signal \N__55431\ : std_logic;
signal \N__55428\ : std_logic;
signal \N__55427\ : std_logic;
signal \N__55426\ : std_logic;
signal \N__55425\ : std_logic;
signal \N__55422\ : std_logic;
signal \N__55421\ : std_logic;
signal \N__55420\ : std_logic;
signal \N__55419\ : std_logic;
signal \N__55418\ : std_logic;
signal \N__55415\ : std_logic;
signal \N__55412\ : std_logic;
signal \N__55409\ : std_logic;
signal \N__55406\ : std_logic;
signal \N__55403\ : std_logic;
signal \N__55400\ : std_logic;
signal \N__55397\ : std_logic;
signal \N__55394\ : std_logic;
signal \N__55393\ : std_logic;
signal \N__55392\ : std_logic;
signal \N__55389\ : std_logic;
signal \N__55380\ : std_logic;
signal \N__55371\ : std_logic;
signal \N__55368\ : std_logic;
signal \N__55361\ : std_logic;
signal \N__55358\ : std_logic;
signal \N__55357\ : std_logic;
signal \N__55356\ : std_logic;
signal \N__55355\ : std_logic;
signal \N__55352\ : std_logic;
signal \N__55351\ : std_logic;
signal \N__55350\ : std_logic;
signal \N__55349\ : std_logic;
signal \N__55348\ : std_logic;
signal \N__55347\ : std_logic;
signal \N__55346\ : std_logic;
signal \N__55345\ : std_logic;
signal \N__55344\ : std_logic;
signal \N__55341\ : std_logic;
signal \N__55340\ : std_logic;
signal \N__55333\ : std_logic;
signal \N__55322\ : std_logic;
signal \N__55319\ : std_logic;
signal \N__55312\ : std_logic;
signal \N__55305\ : std_logic;
signal \N__55294\ : std_logic;
signal \N__55289\ : std_logic;
signal \N__55288\ : std_logic;
signal \N__55287\ : std_logic;
signal \N__55286\ : std_logic;
signal \N__55285\ : std_logic;
signal \N__55284\ : std_logic;
signal \N__55283\ : std_logic;
signal \N__55282\ : std_logic;
signal \N__55281\ : std_logic;
signal \N__55280\ : std_logic;
signal \N__55279\ : std_logic;
signal \N__55278\ : std_logic;
signal \N__55277\ : std_logic;
signal \N__55276\ : std_logic;
signal \N__55275\ : std_logic;
signal \N__55270\ : std_logic;
signal \N__55263\ : std_logic;
signal \N__55252\ : std_logic;
signal \N__55241\ : std_logic;
signal \N__55240\ : std_logic;
signal \N__55237\ : std_logic;
signal \N__55228\ : std_logic;
signal \N__55219\ : std_logic;
signal \N__55218\ : std_logic;
signal \N__55215\ : std_logic;
signal \N__55214\ : std_logic;
signal \N__55213\ : std_logic;
signal \N__55212\ : std_logic;
signal \N__55211\ : std_logic;
signal \N__55210\ : std_logic;
signal \N__55209\ : std_logic;
signal \N__55206\ : std_logic;
signal \N__55205\ : std_logic;
signal \N__55204\ : std_logic;
signal \N__55203\ : std_logic;
signal \N__55192\ : std_logic;
signal \N__55183\ : std_logic;
signal \N__55174\ : std_logic;
signal \N__55167\ : std_logic;
signal \N__55166\ : std_logic;
signal \N__55165\ : std_logic;
signal \N__55164\ : std_logic;
signal \N__55161\ : std_logic;
signal \N__55160\ : std_logic;
signal \N__55159\ : std_logic;
signal \N__55158\ : std_logic;
signal \N__55157\ : std_logic;
signal \N__55152\ : std_logic;
signal \N__55151\ : std_logic;
signal \N__55148\ : std_logic;
signal \N__55141\ : std_logic;
signal \N__55132\ : std_logic;
signal \N__55131\ : std_logic;
signal \N__55130\ : std_logic;
signal \N__55129\ : std_logic;
signal \N__55128\ : std_logic;
signal \N__55127\ : std_logic;
signal \N__55126\ : std_logic;
signal \N__55125\ : std_logic;
signal \N__55122\ : std_logic;
signal \N__55121\ : std_logic;
signal \N__55120\ : std_logic;
signal \N__55119\ : std_logic;
signal \N__55118\ : std_logic;
signal \N__55117\ : std_logic;
signal \N__55110\ : std_logic;
signal \N__55101\ : std_logic;
signal \N__55098\ : std_logic;
signal \N__55097\ : std_logic;
signal \N__55096\ : std_logic;
signal \N__55093\ : std_logic;
signal \N__55092\ : std_logic;
signal \N__55091\ : std_logic;
signal \N__55088\ : std_logic;
signal \N__55087\ : std_logic;
signal \N__55086\ : std_logic;
signal \N__55085\ : std_logic;
signal \N__55084\ : std_logic;
signal \N__55083\ : std_logic;
signal \N__55082\ : std_logic;
signal \N__55081\ : std_logic;
signal \N__55080\ : std_logic;
signal \N__55079\ : std_logic;
signal \N__55078\ : std_logic;
signal \N__55077\ : std_logic;
signal \N__55076\ : std_logic;
signal \N__55073\ : std_logic;
signal \N__55070\ : std_logic;
signal \N__55067\ : std_logic;
signal \N__55066\ : std_logic;
signal \N__55065\ : std_logic;
signal \N__55064\ : std_logic;
signal \N__55063\ : std_logic;
signal \N__55062\ : std_logic;
signal \N__55061\ : std_logic;
signal \N__55060\ : std_logic;
signal \N__55059\ : std_logic;
signal \N__55058\ : std_logic;
signal \N__55057\ : std_logic;
signal \N__55056\ : std_logic;
signal \N__55055\ : std_logic;
signal \N__55046\ : std_logic;
signal \N__55045\ : std_logic;
signal \N__55042\ : std_logic;
signal \N__55041\ : std_logic;
signal \N__55040\ : std_logic;
signal \N__55039\ : std_logic;
signal \N__55038\ : std_logic;
signal \N__55037\ : std_logic;
signal \N__55036\ : std_logic;
signal \N__55035\ : std_logic;
signal \N__55034\ : std_logic;
signal \N__55033\ : std_logic;
signal \N__55032\ : std_logic;
signal \N__55031\ : std_logic;
signal \N__55030\ : std_logic;
signal \N__55023\ : std_logic;
signal \N__55020\ : std_logic;
signal \N__55011\ : std_logic;
signal \N__55004\ : std_logic;
signal \N__54995\ : std_logic;
signal \N__54988\ : std_logic;
signal \N__54985\ : std_logic;
signal \N__54974\ : std_logic;
signal \N__54967\ : std_logic;
signal \N__54964\ : std_logic;
signal \N__54959\ : std_logic;
signal \N__54958\ : std_logic;
signal \N__54957\ : std_logic;
signal \N__54956\ : std_logic;
signal \N__54955\ : std_logic;
signal \N__54954\ : std_logic;
signal \N__54953\ : std_logic;
signal \N__54952\ : std_logic;
signal \N__54947\ : std_logic;
signal \N__54944\ : std_logic;
signal \N__54937\ : std_logic;
signal \N__54932\ : std_logic;
signal \N__54925\ : std_logic;
signal \N__54922\ : std_logic;
signal \N__54915\ : std_logic;
signal \N__54908\ : std_logic;
signal \N__54903\ : std_logic;
signal \N__54894\ : std_logic;
signal \N__54893\ : std_logic;
signal \N__54892\ : std_logic;
signal \N__54891\ : std_logic;
signal \N__54890\ : std_logic;
signal \N__54887\ : std_logic;
signal \N__54884\ : std_logic;
signal \N__54883\ : std_logic;
signal \N__54882\ : std_logic;
signal \N__54881\ : std_logic;
signal \N__54880\ : std_logic;
signal \N__54879\ : std_logic;
signal \N__54878\ : std_logic;
signal \N__54877\ : std_logic;
signal \N__54876\ : std_logic;
signal \N__54875\ : std_logic;
signal \N__54874\ : std_logic;
signal \N__54873\ : std_logic;
signal \N__54872\ : std_logic;
signal \N__54871\ : std_logic;
signal \N__54870\ : std_logic;
signal \N__54869\ : std_logic;
signal \N__54868\ : std_logic;
signal \N__54867\ : std_logic;
signal \N__54866\ : std_logic;
signal \N__54865\ : std_logic;
signal \N__54864\ : std_logic;
signal \N__54863\ : std_logic;
signal \N__54862\ : std_logic;
signal \N__54861\ : std_logic;
signal \N__54860\ : std_logic;
signal \N__54857\ : std_logic;
signal \N__54854\ : std_logic;
signal \N__54851\ : std_logic;
signal \N__54848\ : std_logic;
signal \N__54845\ : std_logic;
signal \N__54842\ : std_logic;
signal \N__54839\ : std_logic;
signal \N__54836\ : std_logic;
signal \N__54833\ : std_logic;
signal \N__54830\ : std_logic;
signal \N__54823\ : std_logic;
signal \N__54820\ : std_logic;
signal \N__54817\ : std_logic;
signal \N__54814\ : std_logic;
signal \N__54813\ : std_logic;
signal \N__54810\ : std_logic;
signal \N__54807\ : std_logic;
signal \N__54804\ : std_logic;
signal \N__54801\ : std_logic;
signal \N__54798\ : std_logic;
signal \N__54795\ : std_logic;
signal \N__54794\ : std_logic;
signal \N__54793\ : std_logic;
signal \N__54792\ : std_logic;
signal \N__54789\ : std_logic;
signal \N__54788\ : std_logic;
signal \N__54787\ : std_logic;
signal \N__54786\ : std_logic;
signal \N__54785\ : std_logic;
signal \N__54784\ : std_logic;
signal \N__54783\ : std_logic;
signal \N__54780\ : std_logic;
signal \N__54777\ : std_logic;
signal \N__54776\ : std_logic;
signal \N__54773\ : std_logic;
signal \N__54770\ : std_logic;
signal \N__54767\ : std_logic;
signal \N__54764\ : std_logic;
signal \N__54763\ : std_logic;
signal \N__54762\ : std_logic;
signal \N__54759\ : std_logic;
signal \N__54758\ : std_logic;
signal \N__54757\ : std_logic;
signal \N__54756\ : std_logic;
signal \N__54753\ : std_logic;
signal \N__54750\ : std_logic;
signal \N__54747\ : std_logic;
signal \N__54746\ : std_logic;
signal \N__54745\ : std_logic;
signal \N__54744\ : std_logic;
signal \N__54743\ : std_logic;
signal \N__54740\ : std_logic;
signal \N__54737\ : std_logic;
signal \N__54736\ : std_logic;
signal \N__54733\ : std_logic;
signal \N__54732\ : std_logic;
signal \N__54731\ : std_logic;
signal \N__54730\ : std_logic;
signal \N__54729\ : std_logic;
signal \N__54728\ : std_logic;
signal \N__54727\ : std_logic;
signal \N__54726\ : std_logic;
signal \N__54725\ : std_logic;
signal \N__54724\ : std_logic;
signal \N__54723\ : std_logic;
signal \N__54722\ : std_logic;
signal \N__54721\ : std_logic;
signal \N__54714\ : std_logic;
signal \N__54713\ : std_logic;
signal \N__54710\ : std_logic;
signal \N__54709\ : std_logic;
signal \N__54708\ : std_logic;
signal \N__54707\ : std_logic;
signal \N__54706\ : std_logic;
signal \N__54705\ : std_logic;
signal \N__54702\ : std_logic;
signal \N__54701\ : std_logic;
signal \N__54700\ : std_logic;
signal \N__54695\ : std_logic;
signal \N__54690\ : std_logic;
signal \N__54677\ : std_logic;
signal \N__54668\ : std_logic;
signal \N__54663\ : std_logic;
signal \N__54662\ : std_logic;
signal \N__54661\ : std_logic;
signal \N__54658\ : std_logic;
signal \N__54657\ : std_logic;
signal \N__54656\ : std_logic;
signal \N__54655\ : std_logic;
signal \N__54654\ : std_logic;
signal \N__54653\ : std_logic;
signal \N__54652\ : std_logic;
signal \N__54651\ : std_logic;
signal \N__54650\ : std_logic;
signal \N__54649\ : std_logic;
signal \N__54648\ : std_logic;
signal \N__54647\ : std_logic;
signal \N__54646\ : std_logic;
signal \N__54645\ : std_logic;
signal \N__54644\ : std_logic;
signal \N__54643\ : std_logic;
signal \N__54640\ : std_logic;
signal \N__54627\ : std_logic;
signal \N__54624\ : std_logic;
signal \N__54621\ : std_logic;
signal \N__54618\ : std_logic;
signal \N__54615\ : std_logic;
signal \N__54608\ : std_logic;
signal \N__54603\ : std_logic;
signal \N__54596\ : std_logic;
signal \N__54593\ : std_logic;
signal \N__54592\ : std_logic;
signal \N__54591\ : std_logic;
signal \N__54590\ : std_logic;
signal \N__54589\ : std_logic;
signal \N__54588\ : std_logic;
signal \N__54587\ : std_logic;
signal \N__54586\ : std_logic;
signal \N__54583\ : std_logic;
signal \N__54582\ : std_logic;
signal \N__54581\ : std_logic;
signal \N__54580\ : std_logic;
signal \N__54579\ : std_logic;
signal \N__54578\ : std_logic;
signal \N__54577\ : std_logic;
signal \N__54576\ : std_logic;
signal \N__54575\ : std_logic;
signal \N__54574\ : std_logic;
signal \N__54573\ : std_logic;
signal \N__54572\ : std_logic;
signal \N__54569\ : std_logic;
signal \N__54566\ : std_logic;
signal \N__54565\ : std_logic;
signal \N__54564\ : std_logic;
signal \N__54561\ : std_logic;
signal \N__54558\ : std_logic;
signal \N__54557\ : std_logic;
signal \N__54556\ : std_logic;
signal \N__54553\ : std_logic;
signal \N__54550\ : std_logic;
signal \N__54547\ : std_logic;
signal \N__54544\ : std_logic;
signal \N__54541\ : std_logic;
signal \N__54538\ : std_logic;
signal \N__54535\ : std_logic;
signal \N__54534\ : std_logic;
signal \N__54531\ : std_logic;
signal \N__54528\ : std_logic;
signal \N__54525\ : std_logic;
signal \N__54522\ : std_logic;
signal \N__54519\ : std_logic;
signal \N__54516\ : std_logic;
signal \N__54515\ : std_logic;
signal \N__54512\ : std_logic;
signal \N__54509\ : std_logic;
signal \N__54508\ : std_logic;
signal \N__54507\ : std_logic;
signal \N__54506\ : std_logic;
signal \N__54499\ : std_logic;
signal \N__54492\ : std_logic;
signal \N__54483\ : std_logic;
signal \N__54480\ : std_logic;
signal \N__54477\ : std_logic;
signal \N__54466\ : std_logic;
signal \N__54457\ : std_logic;
signal \N__54452\ : std_logic;
signal \N__54447\ : std_logic;
signal \N__54446\ : std_logic;
signal \N__54445\ : std_logic;
signal \N__54444\ : std_logic;
signal \N__54443\ : std_logic;
signal \N__54438\ : std_logic;
signal \N__54431\ : std_logic;
signal \N__54424\ : std_logic;
signal \N__54423\ : std_logic;
signal \N__54422\ : std_logic;
signal \N__54421\ : std_logic;
signal \N__54418\ : std_logic;
signal \N__54417\ : std_logic;
signal \N__54416\ : std_logic;
signal \N__54415\ : std_logic;
signal \N__54414\ : std_logic;
signal \N__54407\ : std_logic;
signal \N__54402\ : std_logic;
signal \N__54391\ : std_logic;
signal \N__54382\ : std_logic;
signal \N__54381\ : std_logic;
signal \N__54380\ : std_logic;
signal \N__54379\ : std_logic;
signal \N__54376\ : std_logic;
signal \N__54375\ : std_logic;
signal \N__54374\ : std_logic;
signal \N__54373\ : std_logic;
signal \N__54370\ : std_logic;
signal \N__54369\ : std_logic;
signal \N__54368\ : std_logic;
signal \N__54367\ : std_logic;
signal \N__54364\ : std_logic;
signal \N__54357\ : std_logic;
signal \N__54352\ : std_logic;
signal \N__54351\ : std_logic;
signal \N__54348\ : std_logic;
signal \N__54347\ : std_logic;
signal \N__54346\ : std_logic;
signal \N__54345\ : std_logic;
signal \N__54342\ : std_logic;
signal \N__54339\ : std_logic;
signal \N__54336\ : std_logic;
signal \N__54333\ : std_logic;
signal \N__54330\ : std_logic;
signal \N__54329\ : std_logic;
signal \N__54328\ : std_logic;
signal \N__54327\ : std_logic;
signal \N__54326\ : std_logic;
signal \N__54325\ : std_logic;
signal \N__54324\ : std_logic;
signal \N__54321\ : std_logic;
signal \N__54318\ : std_logic;
signal \N__54315\ : std_logic;
signal \N__54312\ : std_logic;
signal \N__54309\ : std_logic;
signal \N__54306\ : std_logic;
signal \N__54297\ : std_logic;
signal \N__54294\ : std_logic;
signal \N__54293\ : std_logic;
signal \N__54292\ : std_logic;
signal \N__54289\ : std_logic;
signal \N__54288\ : std_logic;
signal \N__54287\ : std_logic;
signal \N__54284\ : std_logic;
signal \N__54283\ : std_logic;
signal \N__54280\ : std_logic;
signal \N__54275\ : std_logic;
signal \N__54270\ : std_logic;
signal \N__54263\ : std_logic;
signal \N__54258\ : std_logic;
signal \N__54253\ : std_logic;
signal \N__54252\ : std_logic;
signal \N__54249\ : std_logic;
signal \N__54248\ : std_logic;
signal \N__54247\ : std_logic;
signal \N__54246\ : std_logic;
signal \N__54245\ : std_logic;
signal \N__54244\ : std_logic;
signal \N__54243\ : std_logic;
signal \N__54242\ : std_logic;
signal \N__54241\ : std_logic;
signal \N__54240\ : std_logic;
signal \N__54237\ : std_logic;
signal \N__54236\ : std_logic;
signal \N__54233\ : std_logic;
signal \N__54230\ : std_logic;
signal \N__54223\ : std_logic;
signal \N__54218\ : std_logic;
signal \N__54215\ : std_logic;
signal \N__54212\ : std_logic;
signal \N__54205\ : std_logic;
signal \N__54186\ : std_logic;
signal \N__54177\ : std_logic;
signal \N__54168\ : std_logic;
signal \N__54163\ : std_logic;
signal \N__54154\ : std_logic;
signal \N__54145\ : std_logic;
signal \N__54140\ : std_logic;
signal \N__54131\ : std_logic;
signal \N__54122\ : std_logic;
signal \N__54113\ : std_logic;
signal \N__54106\ : std_logic;
signal \N__54095\ : std_logic;
signal \N__54090\ : std_logic;
signal \N__54083\ : std_logic;
signal \N__54076\ : std_logic;
signal \N__54075\ : std_logic;
signal \N__54074\ : std_logic;
signal \N__54067\ : std_logic;
signal \N__54058\ : std_logic;
signal \N__54053\ : std_logic;
signal \N__54050\ : std_logic;
signal \N__54043\ : std_logic;
signal \N__54036\ : std_logic;
signal \N__54025\ : std_logic;
signal \N__54024\ : std_logic;
signal \N__54023\ : std_logic;
signal \N__54022\ : std_logic;
signal \N__54021\ : std_logic;
signal \N__54020\ : std_logic;
signal \N__54017\ : std_logic;
signal \N__54014\ : std_logic;
signal \N__54011\ : std_logic;
signal \N__54010\ : std_logic;
signal \N__54001\ : std_logic;
signal \N__53994\ : std_logic;
signal \N__53983\ : std_logic;
signal \N__53982\ : std_logic;
signal \N__53979\ : std_logic;
signal \N__53978\ : std_logic;
signal \N__53977\ : std_logic;
signal \N__53976\ : std_logic;
signal \N__53975\ : std_logic;
signal \N__53972\ : std_logic;
signal \N__53969\ : std_logic;
signal \N__53968\ : std_logic;
signal \N__53967\ : std_logic;
signal \N__53960\ : std_logic;
signal \N__53957\ : std_logic;
signal \N__53950\ : std_logic;
signal \N__53945\ : std_logic;
signal \N__53936\ : std_logic;
signal \N__53935\ : std_logic;
signal \N__53932\ : std_logic;
signal \N__53929\ : std_logic;
signal \N__53926\ : std_logic;
signal \N__53923\ : std_logic;
signal \N__53920\ : std_logic;
signal \N__53919\ : std_logic;
signal \N__53918\ : std_logic;
signal \N__53917\ : std_logic;
signal \N__53910\ : std_logic;
signal \N__53903\ : std_logic;
signal \N__53898\ : std_logic;
signal \N__53891\ : std_logic;
signal \N__53880\ : std_logic;
signal \N__53875\ : std_logic;
signal \N__53868\ : std_logic;
signal \N__53865\ : std_logic;
signal \N__53856\ : std_logic;
signal \N__53855\ : std_logic;
signal \N__53852\ : std_logic;
signal \N__53851\ : std_logic;
signal \N__53850\ : std_logic;
signal \N__53847\ : std_logic;
signal \N__53846\ : std_logic;
signal \N__53843\ : std_logic;
signal \N__53842\ : std_logic;
signal \N__53841\ : std_logic;
signal \N__53838\ : std_logic;
signal \N__53835\ : std_logic;
signal \N__53834\ : std_logic;
signal \N__53831\ : std_logic;
signal \N__53828\ : std_logic;
signal \N__53825\ : std_logic;
signal \N__53820\ : std_logic;
signal \N__53819\ : std_logic;
signal \N__53818\ : std_logic;
signal \N__53817\ : std_logic;
signal \N__53816\ : std_logic;
signal \N__53815\ : std_logic;
signal \N__53814\ : std_logic;
signal \N__53813\ : std_logic;
signal \N__53810\ : std_logic;
signal \N__53799\ : std_logic;
signal \N__53792\ : std_logic;
signal \N__53791\ : std_logic;
signal \N__53790\ : std_logic;
signal \N__53789\ : std_logic;
signal \N__53788\ : std_logic;
signal \N__53787\ : std_logic;
signal \N__53786\ : std_logic;
signal \N__53785\ : std_logic;
signal \N__53778\ : std_logic;
signal \N__53761\ : std_logic;
signal \N__53758\ : std_logic;
signal \N__53753\ : std_logic;
signal \N__53742\ : std_logic;
signal \N__53737\ : std_logic;
signal \N__53728\ : std_logic;
signal \N__53717\ : std_logic;
signal \N__53710\ : std_logic;
signal \N__53705\ : std_logic;
signal \N__53696\ : std_logic;
signal \N__53689\ : std_logic;
signal \N__53686\ : std_logic;
signal \N__53677\ : std_logic;
signal \N__53674\ : std_logic;
signal \N__53667\ : std_logic;
signal \N__53660\ : std_logic;
signal \N__53659\ : std_logic;
signal \N__53656\ : std_logic;
signal \N__53653\ : std_logic;
signal \N__53650\ : std_logic;
signal \N__53649\ : std_logic;
signal \N__53648\ : std_logic;
signal \N__53647\ : std_logic;
signal \N__53646\ : std_logic;
signal \N__53635\ : std_logic;
signal \N__53630\ : std_logic;
signal \N__53625\ : std_logic;
signal \N__53616\ : std_logic;
signal \N__53605\ : std_logic;
signal \N__53594\ : std_logic;
signal \N__53589\ : std_logic;
signal \N__53586\ : std_logic;
signal \N__53579\ : std_logic;
signal \N__53572\ : std_logic;
signal \N__53565\ : std_logic;
signal \N__53562\ : std_logic;
signal \N__53557\ : std_logic;
signal \N__53552\ : std_logic;
signal \N__53547\ : std_logic;
signal \N__53542\ : std_logic;
signal \N__53537\ : std_logic;
signal \N__53528\ : std_logic;
signal \N__53519\ : std_logic;
signal \N__53516\ : std_logic;
signal \N__53513\ : std_logic;
signal \N__53506\ : std_logic;
signal \N__53497\ : std_logic;
signal \N__53494\ : std_logic;
signal \N__53491\ : std_logic;
signal \N__53488\ : std_logic;
signal \N__53485\ : std_logic;
signal \N__53482\ : std_logic;
signal \N__53477\ : std_logic;
signal \N__53472\ : std_logic;
signal \N__53461\ : std_logic;
signal \N__53450\ : std_logic;
signal \N__53445\ : std_logic;
signal \N__53440\ : std_logic;
signal \N__53435\ : std_logic;
signal \N__53430\ : std_logic;
signal \N__53421\ : std_logic;
signal \N__53418\ : std_logic;
signal \N__53415\ : std_logic;
signal \N__53408\ : std_logic;
signal \N__53403\ : std_logic;
signal \N__53396\ : std_logic;
signal \N__53385\ : std_logic;
signal \N__53384\ : std_logic;
signal \N__53381\ : std_logic;
signal \N__53378\ : std_logic;
signal \N__53377\ : std_logic;
signal \N__53374\ : std_logic;
signal \N__53371\ : std_logic;
signal \N__53368\ : std_logic;
signal \N__53365\ : std_logic;
signal \N__53358\ : std_logic;
signal \N__53355\ : std_logic;
signal \N__53352\ : std_logic;
signal \N__53349\ : std_logic;
signal \N__53346\ : std_logic;
signal \N__53345\ : std_logic;
signal \N__53342\ : std_logic;
signal \N__53339\ : std_logic;
signal \N__53336\ : std_logic;
signal \N__53331\ : std_logic;
signal \N__53328\ : std_logic;
signal \N__53327\ : std_logic;
signal \N__53324\ : std_logic;
signal \N__53321\ : std_logic;
signal \N__53318\ : std_logic;
signal \N__53313\ : std_logic;
signal \N__53310\ : std_logic;
signal \N__53309\ : std_logic;
signal \N__53306\ : std_logic;
signal \N__53303\ : std_logic;
signal \N__53300\ : std_logic;
signal \N__53295\ : std_logic;
signal \N__53292\ : std_logic;
signal \N__53289\ : std_logic;
signal \N__53286\ : std_logic;
signal \N__53285\ : std_logic;
signal \N__53282\ : std_logic;
signal \N__53279\ : std_logic;
signal \N__53276\ : std_logic;
signal \N__53271\ : std_logic;
signal \N__53268\ : std_logic;
signal \N__53265\ : std_logic;
signal \N__53264\ : std_logic;
signal \N__53261\ : std_logic;
signal \N__53258\ : std_logic;
signal \N__53255\ : std_logic;
signal \N__53250\ : std_logic;
signal \N__53247\ : std_logic;
signal \N__53246\ : std_logic;
signal \N__53243\ : std_logic;
signal \N__53240\ : std_logic;
signal \N__53237\ : std_logic;
signal \N__53232\ : std_logic;
signal \N__53229\ : std_logic;
signal \N__53226\ : std_logic;
signal \N__53223\ : std_logic;
signal \N__53222\ : std_logic;
signal \N__53221\ : std_logic;
signal \N__53218\ : std_logic;
signal \N__53215\ : std_logic;
signal \N__53212\ : std_logic;
signal \N__53209\ : std_logic;
signal \N__53206\ : std_logic;
signal \N__53203\ : std_logic;
signal \N__53200\ : std_logic;
signal \N__53193\ : std_logic;
signal \N__53190\ : std_logic;
signal \N__53187\ : std_logic;
signal \N__53184\ : std_logic;
signal \N__53181\ : std_logic;
signal \N__53180\ : std_logic;
signal \N__53179\ : std_logic;
signal \N__53176\ : std_logic;
signal \N__53175\ : std_logic;
signal \N__53174\ : std_logic;
signal \N__53173\ : std_logic;
signal \N__53172\ : std_logic;
signal \N__53171\ : std_logic;
signal \N__53168\ : std_logic;
signal \N__53167\ : std_logic;
signal \N__53166\ : std_logic;
signal \N__53163\ : std_logic;
signal \N__53162\ : std_logic;
signal \N__53159\ : std_logic;
signal \N__53156\ : std_logic;
signal \N__53153\ : std_logic;
signal \N__53150\ : std_logic;
signal \N__53145\ : std_logic;
signal \N__53134\ : std_logic;
signal \N__53121\ : std_logic;
signal \N__53118\ : std_logic;
signal \N__53115\ : std_logic;
signal \N__53114\ : std_logic;
signal \N__53113\ : std_logic;
signal \N__53110\ : std_logic;
signal \N__53107\ : std_logic;
signal \N__53104\ : std_logic;
signal \N__53101\ : std_logic;
signal \N__53096\ : std_logic;
signal \N__53091\ : std_logic;
signal \N__53088\ : std_logic;
signal \N__53085\ : std_logic;
signal \N__53084\ : std_logic;
signal \N__53083\ : std_logic;
signal \N__53080\ : std_logic;
signal \N__53075\ : std_logic;
signal \N__53070\ : std_logic;
signal \N__53067\ : std_logic;
signal \N__53064\ : std_logic;
signal \N__53061\ : std_logic;
signal \N__53058\ : std_logic;
signal \N__53055\ : std_logic;
signal \N__53052\ : std_logic;
signal \N__53051\ : std_logic;
signal \N__53050\ : std_logic;
signal \N__53047\ : std_logic;
signal \N__53042\ : std_logic;
signal \N__53039\ : std_logic;
signal \N__53034\ : std_logic;
signal \N__53031\ : std_logic;
signal \N__53028\ : std_logic;
signal \N__53025\ : std_logic;
signal \N__53022\ : std_logic;
signal \N__53021\ : std_logic;
signal \N__53018\ : std_logic;
signal \N__53017\ : std_logic;
signal \N__53014\ : std_logic;
signal \N__53011\ : std_logic;
signal \N__53008\ : std_logic;
signal \N__53005\ : std_logic;
signal \N__53002\ : std_logic;
signal \N__52995\ : std_logic;
signal \N__52992\ : std_logic;
signal \N__52989\ : std_logic;
signal \N__52986\ : std_logic;
signal \N__52983\ : std_logic;
signal \N__52980\ : std_logic;
signal \N__52979\ : std_logic;
signal \N__52976\ : std_logic;
signal \N__52973\ : std_logic;
signal \N__52972\ : std_logic;
signal \N__52969\ : std_logic;
signal \N__52966\ : std_logic;
signal \N__52963\ : std_logic;
signal \N__52960\ : std_logic;
signal \N__52953\ : std_logic;
signal \N__52950\ : std_logic;
signal \N__52947\ : std_logic;
signal \N__52944\ : std_logic;
signal \N__52941\ : std_logic;
signal \N__52938\ : std_logic;
signal \N__52937\ : std_logic;
signal \N__52934\ : std_logic;
signal \N__52931\ : std_logic;
signal \N__52930\ : std_logic;
signal \N__52927\ : std_logic;
signal \N__52924\ : std_logic;
signal \N__52921\ : std_logic;
signal \N__52918\ : std_logic;
signal \N__52911\ : std_logic;
signal \N__52908\ : std_logic;
signal \N__52905\ : std_logic;
signal \N__52902\ : std_logic;
signal \N__52899\ : std_logic;
signal \N__52896\ : std_logic;
signal \N__52895\ : std_logic;
signal \N__52892\ : std_logic;
signal \N__52889\ : std_logic;
signal \N__52886\ : std_logic;
signal \N__52885\ : std_logic;
signal \N__52880\ : std_logic;
signal \N__52877\ : std_logic;
signal \N__52874\ : std_logic;
signal \N__52869\ : std_logic;
signal \N__52866\ : std_logic;
signal \N__52863\ : std_logic;
signal \N__52860\ : std_logic;
signal \N__52859\ : std_logic;
signal \N__52856\ : std_logic;
signal \N__52853\ : std_logic;
signal \N__52852\ : std_logic;
signal \N__52849\ : std_logic;
signal \N__52846\ : std_logic;
signal \N__52843\ : std_logic;
signal \N__52840\ : std_logic;
signal \N__52833\ : std_logic;
signal \N__52830\ : std_logic;
signal \N__52827\ : std_logic;
signal \N__52824\ : std_logic;
signal \N__52821\ : std_logic;
signal \N__52820\ : std_logic;
signal \N__52817\ : std_logic;
signal \N__52814\ : std_logic;
signal \N__52813\ : std_logic;
signal \N__52810\ : std_logic;
signal \N__52807\ : std_logic;
signal \N__52804\ : std_logic;
signal \N__52799\ : std_logic;
signal \N__52794\ : std_logic;
signal \N__52791\ : std_logic;
signal \N__52788\ : std_logic;
signal \N__52785\ : std_logic;
signal \N__52782\ : std_logic;
signal \N__52781\ : std_logic;
signal \N__52778\ : std_logic;
signal \N__52775\ : std_logic;
signal \N__52774\ : std_logic;
signal \N__52771\ : std_logic;
signal \N__52768\ : std_logic;
signal \N__52765\ : std_logic;
signal \N__52762\ : std_logic;
signal \N__52755\ : std_logic;
signal \N__52752\ : std_logic;
signal \N__52749\ : std_logic;
signal \N__52746\ : std_logic;
signal \N__52745\ : std_logic;
signal \N__52742\ : std_logic;
signal \N__52739\ : std_logic;
signal \N__52736\ : std_logic;
signal \N__52733\ : std_logic;
signal \N__52732\ : std_logic;
signal \N__52727\ : std_logic;
signal \N__52724\ : std_logic;
signal \N__52719\ : std_logic;
signal \N__52716\ : std_logic;
signal \N__52713\ : std_logic;
signal \N__52710\ : std_logic;
signal \N__52709\ : std_logic;
signal \N__52706\ : std_logic;
signal \N__52703\ : std_logic;
signal \N__52700\ : std_logic;
signal \N__52697\ : std_logic;
signal \N__52692\ : std_logic;
signal \N__52689\ : std_logic;
signal \N__52686\ : std_logic;
signal \N__52683\ : std_logic;
signal \N__52680\ : std_logic;
signal \N__52679\ : std_logic;
signal \N__52678\ : std_logic;
signal \N__52675\ : std_logic;
signal \N__52670\ : std_logic;
signal \N__52665\ : std_logic;
signal \N__52662\ : std_logic;
signal \N__52659\ : std_logic;
signal \N__52656\ : std_logic;
signal \N__52653\ : std_logic;
signal \N__52652\ : std_logic;
signal \N__52649\ : std_logic;
signal \N__52646\ : std_logic;
signal \N__52641\ : std_logic;
signal \N__52638\ : std_logic;
signal \N__52635\ : std_logic;
signal \N__52632\ : std_logic;
signal \N__52629\ : std_logic;
signal \N__52626\ : std_logic;
signal \N__52623\ : std_logic;
signal \N__52620\ : std_logic;
signal \N__52619\ : std_logic;
signal \N__52616\ : std_logic;
signal \N__52613\ : std_logic;
signal \N__52608\ : std_logic;
signal \N__52605\ : std_logic;
signal \N__52602\ : std_logic;
signal \N__52601\ : std_logic;
signal \N__52598\ : std_logic;
signal \N__52595\ : std_logic;
signal \N__52592\ : std_logic;
signal \N__52589\ : std_logic;
signal \N__52584\ : std_logic;
signal \N__52581\ : std_logic;
signal \N__52578\ : std_logic;
signal \N__52577\ : std_logic;
signal \N__52574\ : std_logic;
signal \N__52571\ : std_logic;
signal \N__52568\ : std_logic;
signal \N__52565\ : std_logic;
signal \N__52562\ : std_logic;
signal \N__52559\ : std_logic;
signal \N__52554\ : std_logic;
signal \N__52551\ : std_logic;
signal \N__52548\ : std_logic;
signal \N__52545\ : std_logic;
signal \N__52542\ : std_logic;
signal \N__52539\ : std_logic;
signal \N__52536\ : std_logic;
signal \N__52533\ : std_logic;
signal \N__52532\ : std_logic;
signal \N__52529\ : std_logic;
signal \N__52526\ : std_logic;
signal \N__52525\ : std_logic;
signal \N__52522\ : std_logic;
signal \N__52519\ : std_logic;
signal \N__52516\ : std_logic;
signal \N__52509\ : std_logic;
signal \N__52506\ : std_logic;
signal \N__52503\ : std_logic;
signal \N__52500\ : std_logic;
signal \N__52497\ : std_logic;
signal \N__52496\ : std_logic;
signal \N__52493\ : std_logic;
signal \N__52490\ : std_logic;
signal \N__52487\ : std_logic;
signal \N__52484\ : std_logic;
signal \N__52479\ : std_logic;
signal \N__52476\ : std_logic;
signal \N__52475\ : std_logic;
signal \N__52472\ : std_logic;
signal \N__52469\ : std_logic;
signal \N__52466\ : std_logic;
signal \N__52463\ : std_logic;
signal \N__52460\ : std_logic;
signal \N__52457\ : std_logic;
signal \N__52454\ : std_logic;
signal \N__52451\ : std_logic;
signal \N__52446\ : std_logic;
signal \N__52443\ : std_logic;
signal \N__52440\ : std_logic;
signal \N__52439\ : std_logic;
signal \N__52436\ : std_logic;
signal \N__52433\ : std_logic;
signal \N__52430\ : std_logic;
signal \N__52427\ : std_logic;
signal \N__52424\ : std_logic;
signal \N__52421\ : std_logic;
signal \N__52416\ : std_logic;
signal \N__52413\ : std_logic;
signal \N__52410\ : std_logic;
signal \N__52409\ : std_logic;
signal \N__52408\ : std_logic;
signal \N__52405\ : std_logic;
signal \N__52402\ : std_logic;
signal \N__52399\ : std_logic;
signal \N__52394\ : std_logic;
signal \N__52389\ : std_logic;
signal \N__52386\ : std_logic;
signal \N__52383\ : std_logic;
signal \N__52380\ : std_logic;
signal \N__52377\ : std_logic;
signal \N__52374\ : std_logic;
signal \N__52371\ : std_logic;
signal \N__52368\ : std_logic;
signal \N__52365\ : std_logic;
signal \N__52362\ : std_logic;
signal \N__52359\ : std_logic;
signal \N__52356\ : std_logic;
signal \N__52353\ : std_logic;
signal \N__52350\ : std_logic;
signal \N__52349\ : std_logic;
signal \N__52348\ : std_logic;
signal \N__52347\ : std_logic;
signal \N__52344\ : std_logic;
signal \N__52343\ : std_logic;
signal \N__52342\ : std_logic;
signal \N__52339\ : std_logic;
signal \N__52338\ : std_logic;
signal \N__52337\ : std_logic;
signal \N__52336\ : std_logic;
signal \N__52333\ : std_logic;
signal \N__52332\ : std_logic;
signal \N__52331\ : std_logic;
signal \N__52328\ : std_logic;
signal \N__52327\ : std_logic;
signal \N__52324\ : std_logic;
signal \N__52319\ : std_logic;
signal \N__52314\ : std_logic;
signal \N__52311\ : std_logic;
signal \N__52304\ : std_logic;
signal \N__52301\ : std_logic;
signal \N__52296\ : std_logic;
signal \N__52281\ : std_logic;
signal \N__52280\ : std_logic;
signal \N__52277\ : std_logic;
signal \N__52276\ : std_logic;
signal \N__52273\ : std_logic;
signal \N__52270\ : std_logic;
signal \N__52267\ : std_logic;
signal \N__52264\ : std_logic;
signal \N__52261\ : std_logic;
signal \N__52258\ : std_logic;
signal \N__52255\ : std_logic;
signal \N__52248\ : std_logic;
signal \N__52247\ : std_logic;
signal \N__52246\ : std_logic;
signal \N__52243\ : std_logic;
signal \N__52240\ : std_logic;
signal \N__52237\ : std_logic;
signal \N__52230\ : std_logic;
signal \N__52227\ : std_logic;
signal \N__52224\ : std_logic;
signal \N__52221\ : std_logic;
signal \N__52218\ : std_logic;
signal \N__52215\ : std_logic;
signal \N__52214\ : std_logic;
signal \N__52211\ : std_logic;
signal \N__52208\ : std_logic;
signal \N__52205\ : std_logic;
signal \N__52202\ : std_logic;
signal \N__52199\ : std_logic;
signal \N__52194\ : std_logic;
signal \N__52191\ : std_logic;
signal \N__52188\ : std_logic;
signal \N__52185\ : std_logic;
signal \N__52182\ : std_logic;
signal \N__52179\ : std_logic;
signal \N__52178\ : std_logic;
signal \N__52177\ : std_logic;
signal \N__52174\ : std_logic;
signal \N__52171\ : std_logic;
signal \N__52168\ : std_logic;
signal \N__52165\ : std_logic;
signal \N__52158\ : std_logic;
signal \N__52155\ : std_logic;
signal \N__52152\ : std_logic;
signal \N__52149\ : std_logic;
signal \N__52148\ : std_logic;
signal \N__52145\ : std_logic;
signal \N__52142\ : std_logic;
signal \N__52141\ : std_logic;
signal \N__52138\ : std_logic;
signal \N__52135\ : std_logic;
signal \N__52132\ : std_logic;
signal \N__52125\ : std_logic;
signal \N__52122\ : std_logic;
signal \N__52119\ : std_logic;
signal \N__52116\ : std_logic;
signal \N__52113\ : std_logic;
signal \N__52110\ : std_logic;
signal \N__52109\ : std_logic;
signal \N__52106\ : std_logic;
signal \N__52105\ : std_logic;
signal \N__52102\ : std_logic;
signal \N__52099\ : std_logic;
signal \N__52096\ : std_logic;
signal \N__52089\ : std_logic;
signal \N__52086\ : std_logic;
signal \N__52083\ : std_logic;
signal \N__52080\ : std_logic;
signal \N__52077\ : std_logic;
signal \N__52076\ : std_logic;
signal \N__52075\ : std_logic;
signal \N__52072\ : std_logic;
signal \N__52069\ : std_logic;
signal \N__52066\ : std_logic;
signal \N__52063\ : std_logic;
signal \N__52060\ : std_logic;
signal \N__52057\ : std_logic;
signal \N__52050\ : std_logic;
signal \N__52047\ : std_logic;
signal \N__52044\ : std_logic;
signal \N__52041\ : std_logic;
signal \N__52038\ : std_logic;
signal \N__52035\ : std_logic;
signal \N__52034\ : std_logic;
signal \N__52031\ : std_logic;
signal \N__52028\ : std_logic;
signal \N__52027\ : std_logic;
signal \N__52024\ : std_logic;
signal \N__52021\ : std_logic;
signal \N__52018\ : std_logic;
signal \N__52011\ : std_logic;
signal \N__52008\ : std_logic;
signal \N__52005\ : std_logic;
signal \N__52002\ : std_logic;
signal \N__51999\ : std_logic;
signal \N__51996\ : std_logic;
signal \N__51993\ : std_logic;
signal \N__51992\ : std_logic;
signal \N__51989\ : std_logic;
signal \N__51986\ : std_logic;
signal \N__51985\ : std_logic;
signal \N__51982\ : std_logic;
signal \N__51979\ : std_logic;
signal \N__51976\ : std_logic;
signal \N__51969\ : std_logic;
signal \N__51966\ : std_logic;
signal \N__51963\ : std_logic;
signal \N__51960\ : std_logic;
signal \N__51957\ : std_logic;
signal \N__51954\ : std_logic;
signal \N__51953\ : std_logic;
signal \N__51950\ : std_logic;
signal \N__51947\ : std_logic;
signal \N__51944\ : std_logic;
signal \N__51943\ : std_logic;
signal \N__51940\ : std_logic;
signal \N__51937\ : std_logic;
signal \N__51934\ : std_logic;
signal \N__51927\ : std_logic;
signal \N__51924\ : std_logic;
signal \N__51921\ : std_logic;
signal \N__51918\ : std_logic;
signal \N__51915\ : std_logic;
signal \N__51912\ : std_logic;
signal \N__51909\ : std_logic;
signal \N__51906\ : std_logic;
signal \N__51905\ : std_logic;
signal \N__51904\ : std_logic;
signal \N__51901\ : std_logic;
signal \N__51896\ : std_logic;
signal \N__51891\ : std_logic;
signal \N__51888\ : std_logic;
signal \N__51885\ : std_logic;
signal \N__51882\ : std_logic;
signal \N__51879\ : std_logic;
signal \N__51876\ : std_logic;
signal \N__51873\ : std_logic;
signal \N__51870\ : std_logic;
signal \N__51867\ : std_logic;
signal \N__51866\ : std_logic;
signal \N__51863\ : std_logic;
signal \N__51860\ : std_logic;
signal \N__51855\ : std_logic;
signal \N__51854\ : std_logic;
signal \N__51851\ : std_logic;
signal \N__51848\ : std_logic;
signal \N__51843\ : std_logic;
signal \N__51840\ : std_logic;
signal \N__51837\ : std_logic;
signal \N__51834\ : std_logic;
signal \N__51833\ : std_logic;
signal \N__51830\ : std_logic;
signal \N__51827\ : std_logic;
signal \N__51824\ : std_logic;
signal \N__51821\ : std_logic;
signal \N__51816\ : std_logic;
signal \N__51815\ : std_logic;
signal \N__51812\ : std_logic;
signal \N__51809\ : std_logic;
signal \N__51804\ : std_logic;
signal \N__51801\ : std_logic;
signal \N__51798\ : std_logic;
signal \N__51795\ : std_logic;
signal \N__51792\ : std_logic;
signal \N__51791\ : std_logic;
signal \N__51788\ : std_logic;
signal \N__51785\ : std_logic;
signal \N__51782\ : std_logic;
signal \N__51781\ : std_logic;
signal \N__51778\ : std_logic;
signal \N__51775\ : std_logic;
signal \N__51772\ : std_logic;
signal \N__51765\ : std_logic;
signal \N__51762\ : std_logic;
signal \N__51759\ : std_logic;
signal \N__51756\ : std_logic;
signal \N__51753\ : std_logic;
signal \N__51750\ : std_logic;
signal \N__51747\ : std_logic;
signal \N__51746\ : std_logic;
signal \N__51743\ : std_logic;
signal \N__51740\ : std_logic;
signal \N__51735\ : std_logic;
signal \N__51732\ : std_logic;
signal \N__51729\ : std_logic;
signal \N__51728\ : std_logic;
signal \N__51725\ : std_logic;
signal \N__51722\ : std_logic;
signal \N__51717\ : std_logic;
signal \N__51714\ : std_logic;
signal \N__51711\ : std_logic;
signal \N__51710\ : std_logic;
signal \N__51707\ : std_logic;
signal \N__51706\ : std_logic;
signal \N__51703\ : std_logic;
signal \N__51700\ : std_logic;
signal \N__51697\ : std_logic;
signal \N__51694\ : std_logic;
signal \N__51689\ : std_logic;
signal \N__51686\ : std_logic;
signal \N__51683\ : std_logic;
signal \N__51678\ : std_logic;
signal \N__51675\ : std_logic;
signal \N__51672\ : std_logic;
signal \N__51669\ : std_logic;
signal \N__51666\ : std_logic;
signal \N__51663\ : std_logic;
signal \N__51662\ : std_logic;
signal \N__51659\ : std_logic;
signal \N__51658\ : std_logic;
signal \N__51655\ : std_logic;
signal \N__51652\ : std_logic;
signal \N__51649\ : std_logic;
signal \N__51642\ : std_logic;
signal \N__51639\ : std_logic;
signal \N__51636\ : std_logic;
signal \N__51633\ : std_logic;
signal \N__51630\ : std_logic;
signal \N__51627\ : std_logic;
signal \N__51626\ : std_logic;
signal \N__51623\ : std_logic;
signal \N__51622\ : std_logic;
signal \N__51619\ : std_logic;
signal \N__51616\ : std_logic;
signal \N__51613\ : std_logic;
signal \N__51606\ : std_logic;
signal \N__51603\ : std_logic;
signal \N__51600\ : std_logic;
signal \N__51597\ : std_logic;
signal \N__51594\ : std_logic;
signal \N__51591\ : std_logic;
signal \N__51590\ : std_logic;
signal \N__51587\ : std_logic;
signal \N__51584\ : std_logic;
signal \N__51581\ : std_logic;
signal \N__51578\ : std_logic;
signal \N__51573\ : std_logic;
signal \N__51570\ : std_logic;
signal \N__51567\ : std_logic;
signal \N__51564\ : std_logic;
signal \N__51561\ : std_logic;
signal \N__51558\ : std_logic;
signal \N__51557\ : std_logic;
signal \N__51554\ : std_logic;
signal \N__51551\ : std_logic;
signal \N__51548\ : std_logic;
signal \N__51545\ : std_logic;
signal \N__51542\ : std_logic;
signal \N__51539\ : std_logic;
signal \N__51538\ : std_logic;
signal \N__51535\ : std_logic;
signal \N__51532\ : std_logic;
signal \N__51529\ : std_logic;
signal \N__51526\ : std_logic;
signal \N__51519\ : std_logic;
signal \N__51516\ : std_logic;
signal \N__51513\ : std_logic;
signal \N__51510\ : std_logic;
signal \N__51507\ : std_logic;
signal \N__51504\ : std_logic;
signal \N__51503\ : std_logic;
signal \N__51500\ : std_logic;
signal \N__51497\ : std_logic;
signal \N__51494\ : std_logic;
signal \N__51489\ : std_logic;
signal \N__51486\ : std_logic;
signal \N__51483\ : std_logic;
signal \N__51480\ : std_logic;
signal \N__51477\ : std_logic;
signal \N__51476\ : std_logic;
signal \N__51473\ : std_logic;
signal \N__51470\ : std_logic;
signal \N__51467\ : std_logic;
signal \N__51466\ : std_logic;
signal \N__51461\ : std_logic;
signal \N__51458\ : std_logic;
signal \N__51455\ : std_logic;
signal \N__51450\ : std_logic;
signal \N__51447\ : std_logic;
signal \N__51444\ : std_logic;
signal \N__51441\ : std_logic;
signal \N__51440\ : std_logic;
signal \N__51437\ : std_logic;
signal \N__51434\ : std_logic;
signal \N__51431\ : std_logic;
signal \N__51428\ : std_logic;
signal \N__51425\ : std_logic;
signal \N__51420\ : std_logic;
signal \N__51417\ : std_logic;
signal \N__51414\ : std_logic;
signal \N__51411\ : std_logic;
signal \N__51408\ : std_logic;
signal \N__51405\ : std_logic;
signal \N__51402\ : std_logic;
signal \N__51399\ : std_logic;
signal \N__51396\ : std_logic;
signal \N__51393\ : std_logic;
signal \N__51392\ : std_logic;
signal \N__51389\ : std_logic;
signal \N__51388\ : std_logic;
signal \N__51385\ : std_logic;
signal \N__51382\ : std_logic;
signal \N__51379\ : std_logic;
signal \N__51372\ : std_logic;
signal \N__51369\ : std_logic;
signal \N__51366\ : std_logic;
signal \N__51363\ : std_logic;
signal \N__51360\ : std_logic;
signal \N__51357\ : std_logic;
signal \N__51356\ : std_logic;
signal \N__51353\ : std_logic;
signal \N__51350\ : std_logic;
signal \N__51347\ : std_logic;
signal \N__51342\ : std_logic;
signal \N__51339\ : std_logic;
signal \N__51336\ : std_logic;
signal \N__51333\ : std_logic;
signal \N__51332\ : std_logic;
signal \N__51329\ : std_logic;
signal \N__51326\ : std_logic;
signal \N__51325\ : std_logic;
signal \N__51322\ : std_logic;
signal \N__51319\ : std_logic;
signal \N__51316\ : std_logic;
signal \N__51309\ : std_logic;
signal \N__51306\ : std_logic;
signal \N__51303\ : std_logic;
signal \N__51300\ : std_logic;
signal \N__51297\ : std_logic;
signal \N__51296\ : std_logic;
signal \N__51293\ : std_logic;
signal \N__51292\ : std_logic;
signal \N__51291\ : std_logic;
signal \N__51288\ : std_logic;
signal \N__51285\ : std_logic;
signal \N__51280\ : std_logic;
signal \N__51273\ : std_logic;
signal \N__51270\ : std_logic;
signal \N__51267\ : std_logic;
signal \N__51266\ : std_logic;
signal \N__51265\ : std_logic;
signal \N__51264\ : std_logic;
signal \N__51261\ : std_logic;
signal \N__51256\ : std_logic;
signal \N__51253\ : std_logic;
signal \N__51250\ : std_logic;
signal \N__51247\ : std_logic;
signal \N__51244\ : std_logic;
signal \N__51241\ : std_logic;
signal \N__51238\ : std_logic;
signal \N__51231\ : std_logic;
signal \N__51228\ : std_logic;
signal \N__51227\ : std_logic;
signal \N__51224\ : std_logic;
signal \N__51221\ : std_logic;
signal \N__51220\ : std_logic;
signal \N__51217\ : std_logic;
signal \N__51216\ : std_logic;
signal \N__51213\ : std_logic;
signal \N__51210\ : std_logic;
signal \N__51207\ : std_logic;
signal \N__51204\ : std_logic;
signal \N__51201\ : std_logic;
signal \N__51192\ : std_logic;
signal \N__51189\ : std_logic;
signal \N__51188\ : std_logic;
signal \N__51187\ : std_logic;
signal \N__51186\ : std_logic;
signal \N__51185\ : std_logic;
signal \N__51182\ : std_logic;
signal \N__51181\ : std_logic;
signal \N__51178\ : std_logic;
signal \N__51177\ : std_logic;
signal \N__51174\ : std_logic;
signal \N__51173\ : std_logic;
signal \N__51170\ : std_logic;
signal \N__51169\ : std_logic;
signal \N__51168\ : std_logic;
signal \N__51167\ : std_logic;
signal \N__51166\ : std_logic;
signal \N__51165\ : std_logic;
signal \N__51164\ : std_logic;
signal \N__51161\ : std_logic;
signal \N__51144\ : std_logic;
signal \N__51143\ : std_logic;
signal \N__51140\ : std_logic;
signal \N__51139\ : std_logic;
signal \N__51136\ : std_logic;
signal \N__51135\ : std_logic;
signal \N__51132\ : std_logic;
signal \N__51131\ : std_logic;
signal \N__51128\ : std_logic;
signal \N__51127\ : std_logic;
signal \N__51126\ : std_logic;
signal \N__51125\ : std_logic;
signal \N__51122\ : std_logic;
signal \N__51121\ : std_logic;
signal \N__51120\ : std_logic;
signal \N__51119\ : std_logic;
signal \N__51118\ : std_logic;
signal \N__51117\ : std_logic;
signal \N__51116\ : std_logic;
signal \N__51115\ : std_logic;
signal \N__51110\ : std_logic;
signal \N__51093\ : std_logic;
signal \N__51084\ : std_logic;
signal \N__51075\ : std_logic;
signal \N__51068\ : std_logic;
signal \N__51057\ : std_logic;
signal \N__51054\ : std_logic;
signal \N__51051\ : std_logic;
signal \N__51050\ : std_logic;
signal \N__51049\ : std_logic;
signal \N__51046\ : std_logic;
signal \N__51043\ : std_logic;
signal \N__51040\ : std_logic;
signal \N__51039\ : std_logic;
signal \N__51038\ : std_logic;
signal \N__51037\ : std_logic;
signal \N__51034\ : std_logic;
signal \N__51031\ : std_logic;
signal \N__51028\ : std_logic;
signal \N__51025\ : std_logic;
signal \N__51022\ : std_logic;
signal \N__51019\ : std_logic;
signal \N__51016\ : std_logic;
signal \N__51013\ : std_logic;
signal \N__51006\ : std_logic;
signal \N__50997\ : std_logic;
signal \N__50994\ : std_logic;
signal \N__50991\ : std_logic;
signal \N__50988\ : std_logic;
signal \N__50985\ : std_logic;
signal \N__50982\ : std_logic;
signal \N__50981\ : std_logic;
signal \N__50980\ : std_logic;
signal \N__50977\ : std_logic;
signal \N__50974\ : std_logic;
signal \N__50971\ : std_logic;
signal \N__50964\ : std_logic;
signal \N__50961\ : std_logic;
signal \N__50958\ : std_logic;
signal \N__50955\ : std_logic;
signal \N__50952\ : std_logic;
signal \N__50951\ : std_logic;
signal \N__50950\ : std_logic;
signal \N__50947\ : std_logic;
signal \N__50944\ : std_logic;
signal \N__50941\ : std_logic;
signal \N__50934\ : std_logic;
signal \N__50933\ : std_logic;
signal \N__50930\ : std_logic;
signal \N__50927\ : std_logic;
signal \N__50924\ : std_logic;
signal \N__50919\ : std_logic;
signal \N__50916\ : std_logic;
signal \N__50913\ : std_logic;
signal \N__50910\ : std_logic;
signal \N__50909\ : std_logic;
signal \N__50908\ : std_logic;
signal \N__50907\ : std_logic;
signal \N__50906\ : std_logic;
signal \N__50905\ : std_logic;
signal \N__50902\ : std_logic;
signal \N__50901\ : std_logic;
signal \N__50900\ : std_logic;
signal \N__50899\ : std_logic;
signal \N__50896\ : std_logic;
signal \N__50895\ : std_logic;
signal \N__50894\ : std_logic;
signal \N__50893\ : std_logic;
signal \N__50892\ : std_logic;
signal \N__50885\ : std_logic;
signal \N__50882\ : std_logic;
signal \N__50879\ : std_logic;
signal \N__50874\ : std_logic;
signal \N__50873\ : std_logic;
signal \N__50870\ : std_logic;
signal \N__50869\ : std_logic;
signal \N__50868\ : std_logic;
signal \N__50867\ : std_logic;
signal \N__50864\ : std_logic;
signal \N__50863\ : std_logic;
signal \N__50858\ : std_logic;
signal \N__50853\ : std_logic;
signal \N__50850\ : std_logic;
signal \N__50847\ : std_logic;
signal \N__50842\ : std_logic;
signal \N__50839\ : std_logic;
signal \N__50838\ : std_logic;
signal \N__50837\ : std_logic;
signal \N__50836\ : std_logic;
signal \N__50835\ : std_logic;
signal \N__50834\ : std_logic;
signal \N__50833\ : std_logic;
signal \N__50832\ : std_logic;
signal \N__50829\ : std_logic;
signal \N__50822\ : std_logic;
signal \N__50819\ : std_logic;
signal \N__50816\ : std_logic;
signal \N__50811\ : std_logic;
signal \N__50806\ : std_logic;
signal \N__50801\ : std_logic;
signal \N__50798\ : std_logic;
signal \N__50795\ : std_logic;
signal \N__50792\ : std_logic;
signal \N__50789\ : std_logic;
signal \N__50782\ : std_logic;
signal \N__50773\ : std_logic;
signal \N__50754\ : std_logic;
signal \N__50751\ : std_logic;
signal \N__50750\ : std_logic;
signal \N__50747\ : std_logic;
signal \N__50744\ : std_logic;
signal \N__50743\ : std_logic;
signal \N__50740\ : std_logic;
signal \N__50737\ : std_logic;
signal \N__50734\ : std_logic;
signal \N__50731\ : std_logic;
signal \N__50728\ : std_logic;
signal \N__50725\ : std_logic;
signal \N__50718\ : std_logic;
signal \N__50715\ : std_logic;
signal \N__50712\ : std_logic;
signal \N__50709\ : std_logic;
signal \N__50706\ : std_logic;
signal \N__50705\ : std_logic;
signal \N__50704\ : std_logic;
signal \N__50701\ : std_logic;
signal \N__50700\ : std_logic;
signal \N__50697\ : std_logic;
signal \N__50694\ : std_logic;
signal \N__50691\ : std_logic;
signal \N__50686\ : std_logic;
signal \N__50679\ : std_logic;
signal \N__50676\ : std_logic;
signal \N__50675\ : std_logic;
signal \N__50674\ : std_logic;
signal \N__50671\ : std_logic;
signal \N__50670\ : std_logic;
signal \N__50667\ : std_logic;
signal \N__50664\ : std_logic;
signal \N__50661\ : std_logic;
signal \N__50658\ : std_logic;
signal \N__50655\ : std_logic;
signal \N__50652\ : std_logic;
signal \N__50647\ : std_logic;
signal \N__50640\ : std_logic;
signal \N__50637\ : std_logic;
signal \N__50634\ : std_logic;
signal \N__50631\ : std_logic;
signal \N__50630\ : std_logic;
signal \N__50629\ : std_logic;
signal \N__50626\ : std_logic;
signal \N__50625\ : std_logic;
signal \N__50622\ : std_logic;
signal \N__50619\ : std_logic;
signal \N__50616\ : std_logic;
signal \N__50613\ : std_logic;
signal \N__50610\ : std_logic;
signal \N__50601\ : std_logic;
signal \N__50598\ : std_logic;
signal \N__50597\ : std_logic;
signal \N__50594\ : std_logic;
signal \N__50591\ : std_logic;
signal \N__50588\ : std_logic;
signal \N__50587\ : std_logic;
signal \N__50586\ : std_logic;
signal \N__50583\ : std_logic;
signal \N__50580\ : std_logic;
signal \N__50575\ : std_logic;
signal \N__50568\ : std_logic;
signal \N__50565\ : std_logic;
signal \N__50562\ : std_logic;
signal \N__50559\ : std_logic;
signal \N__50558\ : std_logic;
signal \N__50557\ : std_logic;
signal \N__50554\ : std_logic;
signal \N__50551\ : std_logic;
signal \N__50548\ : std_logic;
signal \N__50545\ : std_logic;
signal \N__50544\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50535\ : std_logic;
signal \N__50532\ : std_logic;
signal \N__50527\ : std_logic;
signal \N__50520\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50514\ : std_logic;
signal \N__50511\ : std_logic;
signal \N__50510\ : std_logic;
signal \N__50509\ : std_logic;
signal \N__50506\ : std_logic;
signal \N__50505\ : std_logic;
signal \N__50502\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50496\ : std_logic;
signal \N__50491\ : std_logic;
signal \N__50484\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50478\ : std_logic;
signal \N__50477\ : std_logic;
signal \N__50476\ : std_logic;
signal \N__50473\ : std_logic;
signal \N__50470\ : std_logic;
signal \N__50467\ : std_logic;
signal \N__50464\ : std_logic;
signal \N__50463\ : std_logic;
signal \N__50460\ : std_logic;
signal \N__50457\ : std_logic;
signal \N__50454\ : std_logic;
signal \N__50451\ : std_logic;
signal \N__50446\ : std_logic;
signal \N__50439\ : std_logic;
signal \N__50436\ : std_logic;
signal \N__50433\ : std_logic;
signal \N__50430\ : std_logic;
signal \N__50429\ : std_logic;
signal \N__50426\ : std_logic;
signal \N__50423\ : std_logic;
signal \N__50420\ : std_logic;
signal \N__50419\ : std_logic;
signal \N__50418\ : std_logic;
signal \N__50413\ : std_logic;
signal \N__50410\ : std_logic;
signal \N__50407\ : std_logic;
signal \N__50400\ : std_logic;
signal \N__50397\ : std_logic;
signal \N__50396\ : std_logic;
signal \N__50393\ : std_logic;
signal \N__50392\ : std_logic;
signal \N__50391\ : std_logic;
signal \N__50388\ : std_logic;
signal \N__50385\ : std_logic;
signal \N__50382\ : std_logic;
signal \N__50379\ : std_logic;
signal \N__50376\ : std_logic;
signal \N__50371\ : std_logic;
signal \N__50368\ : std_logic;
signal \N__50365\ : std_logic;
signal \N__50362\ : std_logic;
signal \N__50355\ : std_logic;
signal \N__50352\ : std_logic;
signal \N__50351\ : std_logic;
signal \N__50348\ : std_logic;
signal \N__50347\ : std_logic;
signal \N__50344\ : std_logic;
signal \N__50341\ : std_logic;
signal \N__50338\ : std_logic;
signal \N__50335\ : std_logic;
signal \N__50332\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50322\ : std_logic;
signal \N__50319\ : std_logic;
signal \N__50318\ : std_logic;
signal \N__50317\ : std_logic;
signal \N__50314\ : std_logic;
signal \N__50311\ : std_logic;
signal \N__50310\ : std_logic;
signal \N__50307\ : std_logic;
signal \N__50304\ : std_logic;
signal \N__50301\ : std_logic;
signal \N__50298\ : std_logic;
signal \N__50295\ : std_logic;
signal \N__50292\ : std_logic;
signal \N__50289\ : std_logic;
signal \N__50286\ : std_logic;
signal \N__50277\ : std_logic;
signal \N__50274\ : std_logic;
signal \N__50271\ : std_logic;
signal \N__50270\ : std_logic;
signal \N__50267\ : std_logic;
signal \N__50266\ : std_logic;
signal \N__50265\ : std_logic;
signal \N__50262\ : std_logic;
signal \N__50259\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50246\ : std_logic;
signal \N__50241\ : std_logic;
signal \N__50238\ : std_logic;
signal \N__50237\ : std_logic;
signal \N__50234\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50232\ : std_logic;
signal \N__50229\ : std_logic;
signal \N__50226\ : std_logic;
signal \N__50221\ : std_logic;
signal \N__50218\ : std_logic;
signal \N__50215\ : std_logic;
signal \N__50212\ : std_logic;
signal \N__50205\ : std_logic;
signal \N__50202\ : std_logic;
signal \N__50199\ : std_logic;
signal \N__50198\ : std_logic;
signal \N__50195\ : std_logic;
signal \N__50192\ : std_logic;
signal \N__50191\ : std_logic;
signal \N__50188\ : std_logic;
signal \N__50185\ : std_logic;
signal \N__50182\ : std_logic;
signal \N__50181\ : std_logic;
signal \N__50178\ : std_logic;
signal \N__50173\ : std_logic;
signal \N__50170\ : std_logic;
signal \N__50165\ : std_logic;
signal \N__50160\ : std_logic;
signal \N__50157\ : std_logic;
signal \N__50154\ : std_logic;
signal \N__50153\ : std_logic;
signal \N__50152\ : std_logic;
signal \N__50151\ : std_logic;
signal \N__50148\ : std_logic;
signal \N__50145\ : std_logic;
signal \N__50142\ : std_logic;
signal \N__50139\ : std_logic;
signal \N__50134\ : std_logic;
signal \N__50131\ : std_logic;
signal \N__50126\ : std_logic;
signal \N__50121\ : std_logic;
signal \N__50118\ : std_logic;
signal \N__50117\ : std_logic;
signal \N__50114\ : std_logic;
signal \N__50111\ : std_logic;
signal \N__50108\ : std_logic;
signal \N__50107\ : std_logic;
signal \N__50106\ : std_logic;
signal \N__50103\ : std_logic;
signal \N__50100\ : std_logic;
signal \N__50097\ : std_logic;
signal \N__50094\ : std_logic;
signal \N__50091\ : std_logic;
signal \N__50086\ : std_logic;
signal \N__50079\ : std_logic;
signal \N__50076\ : std_logic;
signal \N__50073\ : std_logic;
signal \N__50072\ : std_logic;
signal \N__50071\ : std_logic;
signal \N__50070\ : std_logic;
signal \N__50067\ : std_logic;
signal \N__50062\ : std_logic;
signal \N__50059\ : std_logic;
signal \N__50056\ : std_logic;
signal \N__50053\ : std_logic;
signal \N__50050\ : std_logic;
signal \N__50047\ : std_logic;
signal \N__50044\ : std_logic;
signal \N__50037\ : std_logic;
signal \N__50034\ : std_logic;
signal \N__50033\ : std_logic;
signal \N__50030\ : std_logic;
signal \N__50027\ : std_logic;
signal \N__50026\ : std_logic;
signal \N__50023\ : std_logic;
signal \N__50020\ : std_logic;
signal \N__50017\ : std_logic;
signal \N__50010\ : std_logic;
signal \N__50007\ : std_logic;
signal \N__50004\ : std_logic;
signal \N__50001\ : std_logic;
signal \N__50000\ : std_logic;
signal \N__49999\ : std_logic;
signal \N__49996\ : std_logic;
signal \N__49991\ : std_logic;
signal \N__49986\ : std_logic;
signal \N__49983\ : std_logic;
signal \N__49980\ : std_logic;
signal \N__49979\ : std_logic;
signal \N__49976\ : std_logic;
signal \N__49973\ : std_logic;
signal \N__49970\ : std_logic;
signal \N__49967\ : std_logic;
signal \N__49962\ : std_logic;
signal \N__49959\ : std_logic;
signal \N__49956\ : std_logic;
signal \N__49953\ : std_logic;
signal \N__49950\ : std_logic;
signal \N__49947\ : std_logic;
signal \N__49944\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49942\ : std_logic;
signal \N__49941\ : std_logic;
signal \N__49938\ : std_logic;
signal \N__49935\ : std_logic;
signal \N__49934\ : std_logic;
signal \N__49931\ : std_logic;
signal \N__49930\ : std_logic;
signal \N__49929\ : std_logic;
signal \N__49928\ : std_logic;
signal \N__49925\ : std_logic;
signal \N__49924\ : std_logic;
signal \N__49923\ : std_logic;
signal \N__49922\ : std_logic;
signal \N__49919\ : std_logic;
signal \N__49916\ : std_logic;
signal \N__49913\ : std_logic;
signal \N__49904\ : std_logic;
signal \N__49901\ : std_logic;
signal \N__49894\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49878\ : std_logic;
signal \N__49877\ : std_logic;
signal \N__49876\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49872\ : std_logic;
signal \N__49869\ : std_logic;
signal \N__49868\ : std_logic;
signal \N__49867\ : std_logic;
signal \N__49864\ : std_logic;
signal \N__49861\ : std_logic;
signal \N__49860\ : std_logic;
signal \N__49855\ : std_logic;
signal \N__49854\ : std_logic;
signal \N__49851\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49843\ : std_logic;
signal \N__49842\ : std_logic;
signal \N__49841\ : std_logic;
signal \N__49838\ : std_logic;
signal \N__49835\ : std_logic;
signal \N__49832\ : std_logic;
signal \N__49827\ : std_logic;
signal \N__49824\ : std_logic;
signal \N__49817\ : std_logic;
signal \N__49806\ : std_logic;
signal \N__49805\ : std_logic;
signal \N__49802\ : std_logic;
signal \N__49801\ : std_logic;
signal \N__49798\ : std_logic;
signal \N__49795\ : std_logic;
signal \N__49792\ : std_logic;
signal \N__49789\ : std_logic;
signal \N__49782\ : std_logic;
signal \N__49779\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49770\ : std_logic;
signal \N__49767\ : std_logic;
signal \N__49764\ : std_logic;
signal \N__49763\ : std_logic;
signal \N__49762\ : std_logic;
signal \N__49759\ : std_logic;
signal \N__49756\ : std_logic;
signal \N__49753\ : std_logic;
signal \N__49748\ : std_logic;
signal \N__49743\ : std_logic;
signal \N__49740\ : std_logic;
signal \N__49737\ : std_logic;
signal \N__49736\ : std_logic;
signal \N__49735\ : std_logic;
signal \N__49732\ : std_logic;
signal \N__49729\ : std_logic;
signal \N__49726\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49720\ : std_logic;
signal \N__49717\ : std_logic;
signal \N__49712\ : std_logic;
signal \N__49707\ : std_logic;
signal \N__49704\ : std_logic;
signal \N__49703\ : std_logic;
signal \N__49700\ : std_logic;
signal \N__49699\ : std_logic;
signal \N__49696\ : std_logic;
signal \N__49693\ : std_logic;
signal \N__49690\ : std_logic;
signal \N__49687\ : std_logic;
signal \N__49684\ : std_logic;
signal \N__49681\ : std_logic;
signal \N__49674\ : std_logic;
signal \N__49671\ : std_logic;
signal \N__49668\ : std_logic;
signal \N__49665\ : std_logic;
signal \N__49664\ : std_logic;
signal \N__49661\ : std_logic;
signal \N__49658\ : std_logic;
signal \N__49657\ : std_logic;
signal \N__49654\ : std_logic;
signal \N__49651\ : std_logic;
signal \N__49648\ : std_logic;
signal \N__49641\ : std_logic;
signal \N__49638\ : std_logic;
signal \N__49635\ : std_logic;
signal \N__49632\ : std_logic;
signal \N__49629\ : std_logic;
signal \N__49626\ : std_logic;
signal \N__49625\ : std_logic;
signal \N__49624\ : std_logic;
signal \N__49623\ : std_logic;
signal \N__49622\ : std_logic;
signal \N__49621\ : std_logic;
signal \N__49612\ : std_logic;
signal \N__49611\ : std_logic;
signal \N__49610\ : std_logic;
signal \N__49607\ : std_logic;
signal \N__49606\ : std_logic;
signal \N__49605\ : std_logic;
signal \N__49604\ : std_logic;
signal \N__49603\ : std_logic;
signal \N__49602\ : std_logic;
signal \N__49601\ : std_logic;
signal \N__49600\ : std_logic;
signal \N__49599\ : std_logic;
signal \N__49598\ : std_logic;
signal \N__49597\ : std_logic;
signal \N__49594\ : std_logic;
signal \N__49593\ : std_logic;
signal \N__49592\ : std_logic;
signal \N__49591\ : std_logic;
signal \N__49590\ : std_logic;
signal \N__49589\ : std_logic;
signal \N__49586\ : std_logic;
signal \N__49581\ : std_logic;
signal \N__49580\ : std_logic;
signal \N__49577\ : std_logic;
signal \N__49574\ : std_logic;
signal \N__49569\ : std_logic;
signal \N__49566\ : std_logic;
signal \N__49561\ : std_logic;
signal \N__49560\ : std_logic;
signal \N__49557\ : std_logic;
signal \N__49554\ : std_logic;
signal \N__49553\ : std_logic;
signal \N__49552\ : std_logic;
signal \N__49549\ : std_logic;
signal \N__49548\ : std_logic;
signal \N__49547\ : std_logic;
signal \N__49546\ : std_logic;
signal \N__49543\ : std_logic;
signal \N__49542\ : std_logic;
signal \N__49541\ : std_logic;
signal \N__49540\ : std_logic;
signal \N__49539\ : std_logic;
signal \N__49538\ : std_logic;
signal \N__49535\ : std_logic;
signal \N__49528\ : std_logic;
signal \N__49523\ : std_logic;
signal \N__49518\ : std_logic;
signal \N__49517\ : std_logic;
signal \N__49514\ : std_logic;
signal \N__49513\ : std_logic;
signal \N__49508\ : std_logic;
signal \N__49505\ : std_logic;
signal \N__49500\ : std_logic;
signal \N__49497\ : std_logic;
signal \N__49496\ : std_logic;
signal \N__49495\ : std_logic;
signal \N__49494\ : std_logic;
signal \N__49493\ : std_logic;
signal \N__49488\ : std_logic;
signal \N__49485\ : std_logic;
signal \N__49482\ : std_logic;
signal \N__49469\ : std_logic;
signal \N__49466\ : std_logic;
signal \N__49463\ : std_logic;
signal \N__49460\ : std_logic;
signal \N__49457\ : std_logic;
signal \N__49452\ : std_logic;
signal \N__49447\ : std_logic;
signal \N__49440\ : std_logic;
signal \N__49437\ : std_logic;
signal \N__49430\ : std_logic;
signal \N__49427\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49412\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49380\ : std_logic;
signal \N__49377\ : std_logic;
signal \N__49376\ : std_logic;
signal \N__49373\ : std_logic;
signal \N__49370\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49366\ : std_logic;
signal \N__49363\ : std_logic;
signal \N__49360\ : std_logic;
signal \N__49353\ : std_logic;
signal \N__49350\ : std_logic;
signal \N__49347\ : std_logic;
signal \N__49344\ : std_logic;
signal \N__49341\ : std_logic;
signal \N__49338\ : std_logic;
signal \N__49335\ : std_logic;
signal \N__49332\ : std_logic;
signal \N__49329\ : std_logic;
signal \N__49328\ : std_logic;
signal \N__49325\ : std_logic;
signal \N__49322\ : std_logic;
signal \N__49319\ : std_logic;
signal \N__49316\ : std_logic;
signal \N__49311\ : std_logic;
signal \N__49308\ : std_logic;
signal \N__49307\ : std_logic;
signal \N__49304\ : std_logic;
signal \N__49301\ : std_logic;
signal \N__49296\ : std_logic;
signal \N__49293\ : std_logic;
signal \N__49290\ : std_logic;
signal \N__49287\ : std_logic;
signal \N__49286\ : std_logic;
signal \N__49283\ : std_logic;
signal \N__49280\ : std_logic;
signal \N__49277\ : std_logic;
signal \N__49274\ : std_logic;
signal \N__49269\ : std_logic;
signal \N__49266\ : std_logic;
signal \N__49263\ : std_logic;
signal \N__49260\ : std_logic;
signal \N__49257\ : std_logic;
signal \N__49256\ : std_logic;
signal \N__49253\ : std_logic;
signal \N__49250\ : std_logic;
signal \N__49249\ : std_logic;
signal \N__49246\ : std_logic;
signal \N__49243\ : std_logic;
signal \N__49240\ : std_logic;
signal \N__49233\ : std_logic;
signal \N__49232\ : std_logic;
signal \N__49229\ : std_logic;
signal \N__49226\ : std_logic;
signal \N__49225\ : std_logic;
signal \N__49222\ : std_logic;
signal \N__49217\ : std_logic;
signal \N__49212\ : std_logic;
signal \N__49209\ : std_logic;
signal \N__49208\ : std_logic;
signal \N__49205\ : std_logic;
signal \N__49202\ : std_logic;
signal \N__49197\ : std_logic;
signal \N__49194\ : std_logic;
signal \N__49191\ : std_logic;
signal \N__49188\ : std_logic;
signal \N__49185\ : std_logic;
signal \N__49184\ : std_logic;
signal \N__49181\ : std_logic;
signal \N__49178\ : std_logic;
signal \N__49177\ : std_logic;
signal \N__49174\ : std_logic;
signal \N__49171\ : std_logic;
signal \N__49168\ : std_logic;
signal \N__49161\ : std_logic;
signal \N__49158\ : std_logic;
signal \N__49155\ : std_logic;
signal \N__49152\ : std_logic;
signal \N__49149\ : std_logic;
signal \N__49146\ : std_logic;
signal \N__49143\ : std_logic;
signal \N__49140\ : std_logic;
signal \N__49139\ : std_logic;
signal \N__49138\ : std_logic;
signal \N__49135\ : std_logic;
signal \N__49132\ : std_logic;
signal \N__49129\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49121\ : std_logic;
signal \N__49118\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49104\ : std_logic;
signal \N__49101\ : std_logic;
signal \N__49098\ : std_logic;
signal \N__49095\ : std_logic;
signal \N__49092\ : std_logic;
signal \N__49089\ : std_logic;
signal \N__49086\ : std_logic;
signal \N__49083\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49079\ : std_logic;
signal \N__49076\ : std_logic;
signal \N__49075\ : std_logic;
signal \N__49072\ : std_logic;
signal \N__49069\ : std_logic;
signal \N__49064\ : std_logic;
signal \N__49059\ : std_logic;
signal \N__49056\ : std_logic;
signal \N__49053\ : std_logic;
signal \N__49050\ : std_logic;
signal \N__49047\ : std_logic;
signal \N__49044\ : std_logic;
signal \N__49041\ : std_logic;
signal \N__49038\ : std_logic;
signal \N__49035\ : std_logic;
signal \N__49032\ : std_logic;
signal \N__49029\ : std_logic;
signal \N__49026\ : std_logic;
signal \N__49023\ : std_logic;
signal \N__49020\ : std_logic;
signal \N__49017\ : std_logic;
signal \N__49014\ : std_logic;
signal \N__49011\ : std_logic;
signal \N__49008\ : std_logic;
signal \N__49007\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__49001\ : std_logic;
signal \N__49000\ : std_logic;
signal \N__48999\ : std_logic;
signal \N__48998\ : std_logic;
signal \N__48997\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48993\ : std_logic;
signal \N__48992\ : std_logic;
signal \N__48991\ : std_logic;
signal \N__48988\ : std_logic;
signal \N__48987\ : std_logic;
signal \N__48984\ : std_logic;
signal \N__48981\ : std_logic;
signal \N__48980\ : std_logic;
signal \N__48977\ : std_logic;
signal \N__48976\ : std_logic;
signal \N__48973\ : std_logic;
signal \N__48972\ : std_logic;
signal \N__48969\ : std_logic;
signal \N__48966\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48958\ : std_logic;
signal \N__48941\ : std_logic;
signal \N__48930\ : std_logic;
signal \N__48927\ : std_logic;
signal \N__48926\ : std_logic;
signal \N__48923\ : std_logic;
signal \N__48920\ : std_logic;
signal \N__48917\ : std_logic;
signal \N__48914\ : std_logic;
signal \N__48913\ : std_logic;
signal \N__48908\ : std_logic;
signal \N__48905\ : std_logic;
signal \N__48900\ : std_logic;
signal \N__48897\ : std_logic;
signal \N__48894\ : std_logic;
signal \N__48893\ : std_logic;
signal \N__48890\ : std_logic;
signal \N__48887\ : std_logic;
signal \N__48886\ : std_logic;
signal \N__48885\ : std_logic;
signal \N__48884\ : std_logic;
signal \N__48881\ : std_logic;
signal \N__48878\ : std_logic;
signal \N__48877\ : std_logic;
signal \N__48876\ : std_logic;
signal \N__48875\ : std_logic;
signal \N__48874\ : std_logic;
signal \N__48871\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48866\ : std_logic;
signal \N__48863\ : std_logic;
signal \N__48862\ : std_logic;
signal \N__48861\ : std_logic;
signal \N__48860\ : std_logic;
signal \N__48857\ : std_logic;
signal \N__48854\ : std_logic;
signal \N__48851\ : std_logic;
signal \N__48844\ : std_logic;
signal \N__48839\ : std_logic;
signal \N__48834\ : std_logic;
signal \N__48825\ : std_logic;
signal \N__48810\ : std_logic;
signal \N__48809\ : std_logic;
signal \N__48806\ : std_logic;
signal \N__48803\ : std_logic;
signal \N__48800\ : std_logic;
signal \N__48797\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48789\ : std_logic;
signal \N__48788\ : std_logic;
signal \N__48787\ : std_logic;
signal \N__48784\ : std_logic;
signal \N__48781\ : std_logic;
signal \N__48778\ : std_logic;
signal \N__48775\ : std_logic;
signal \N__48770\ : std_logic;
signal \N__48767\ : std_logic;
signal \N__48764\ : std_logic;
signal \N__48759\ : std_logic;
signal \N__48756\ : std_logic;
signal \N__48753\ : std_logic;
signal \N__48750\ : std_logic;
signal \N__48749\ : std_logic;
signal \N__48746\ : std_logic;
signal \N__48743\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48733\ : std_logic;
signal \N__48726\ : std_logic;
signal \N__48723\ : std_logic;
signal \N__48720\ : std_logic;
signal \N__48717\ : std_logic;
signal \N__48714\ : std_logic;
signal \N__48711\ : std_logic;
signal \N__48708\ : std_logic;
signal \N__48705\ : std_logic;
signal \N__48702\ : std_logic;
signal \N__48699\ : std_logic;
signal \N__48696\ : std_logic;
signal \N__48695\ : std_logic;
signal \N__48694\ : std_logic;
signal \N__48693\ : std_logic;
signal \N__48690\ : std_logic;
signal \N__48687\ : std_logic;
signal \N__48684\ : std_logic;
signal \N__48681\ : std_logic;
signal \N__48672\ : std_logic;
signal \N__48671\ : std_logic;
signal \N__48668\ : std_logic;
signal \N__48665\ : std_logic;
signal \N__48660\ : std_logic;
signal \N__48659\ : std_logic;
signal \N__48656\ : std_logic;
signal \N__48653\ : std_logic;
signal \N__48648\ : std_logic;
signal \N__48647\ : std_logic;
signal \N__48644\ : std_logic;
signal \N__48641\ : std_logic;
signal \N__48638\ : std_logic;
signal \N__48633\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48629\ : std_logic;
signal \N__48626\ : std_logic;
signal \N__48621\ : std_logic;
signal \N__48620\ : std_logic;
signal \N__48617\ : std_logic;
signal \N__48614\ : std_logic;
signal \N__48609\ : std_logic;
signal \N__48608\ : std_logic;
signal \N__48605\ : std_logic;
signal \N__48602\ : std_logic;
signal \N__48597\ : std_logic;
signal \N__48594\ : std_logic;
signal \N__48593\ : std_logic;
signal \N__48590\ : std_logic;
signal \N__48587\ : std_logic;
signal \N__48582\ : std_logic;
signal \N__48579\ : std_logic;
signal \N__48578\ : std_logic;
signal \N__48577\ : std_logic;
signal \N__48574\ : std_logic;
signal \N__48571\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48565\ : std_logic;
signal \N__48558\ : std_logic;
signal \N__48555\ : std_logic;
signal \N__48554\ : std_logic;
signal \N__48551\ : std_logic;
signal \N__48550\ : std_logic;
signal \N__48547\ : std_logic;
signal \N__48544\ : std_logic;
signal \N__48541\ : std_logic;
signal \N__48536\ : std_logic;
signal \N__48531\ : std_logic;
signal \N__48528\ : std_logic;
signal \N__48527\ : std_logic;
signal \N__48526\ : std_logic;
signal \N__48523\ : std_logic;
signal \N__48520\ : std_logic;
signal \N__48517\ : std_logic;
signal \N__48514\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48501\ : std_logic;
signal \N__48500\ : std_logic;
signal \N__48499\ : std_logic;
signal \N__48496\ : std_logic;
signal \N__48493\ : std_logic;
signal \N__48490\ : std_logic;
signal \N__48487\ : std_logic;
signal \N__48480\ : std_logic;
signal \N__48477\ : std_logic;
signal \N__48476\ : std_logic;
signal \N__48475\ : std_logic;
signal \N__48472\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48464\ : std_logic;
signal \N__48463\ : std_logic;
signal \N__48462\ : std_logic;
signal \N__48459\ : std_logic;
signal \N__48456\ : std_logic;
signal \N__48453\ : std_logic;
signal \N__48450\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48444\ : std_logic;
signal \N__48435\ : std_logic;
signal \N__48432\ : std_logic;
signal \N__48429\ : std_logic;
signal \N__48428\ : std_logic;
signal \N__48427\ : std_logic;
signal \N__48424\ : std_logic;
signal \N__48421\ : std_logic;
signal \N__48418\ : std_logic;
signal \N__48415\ : std_logic;
signal \N__48408\ : std_logic;
signal \N__48405\ : std_logic;
signal \N__48402\ : std_logic;
signal \N__48399\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48395\ : std_logic;
signal \N__48394\ : std_logic;
signal \N__48393\ : std_logic;
signal \N__48388\ : std_logic;
signal \N__48385\ : std_logic;
signal \N__48382\ : std_logic;
signal \N__48379\ : std_logic;
signal \N__48372\ : std_logic;
signal \N__48369\ : std_logic;
signal \N__48368\ : std_logic;
signal \N__48367\ : std_logic;
signal \N__48364\ : std_logic;
signal \N__48361\ : std_logic;
signal \N__48358\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48348\ : std_logic;
signal \N__48345\ : std_logic;
signal \N__48344\ : std_logic;
signal \N__48341\ : std_logic;
signal \N__48340\ : std_logic;
signal \N__48337\ : std_logic;
signal \N__48334\ : std_logic;
signal \N__48331\ : std_logic;
signal \N__48328\ : std_logic;
signal \N__48321\ : std_logic;
signal \N__48318\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48313\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48307\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48301\ : std_logic;
signal \N__48294\ : std_logic;
signal \N__48291\ : std_logic;
signal \N__48290\ : std_logic;
signal \N__48289\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48280\ : std_logic;
signal \N__48273\ : std_logic;
signal \N__48270\ : std_logic;
signal \N__48267\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48265\ : std_logic;
signal \N__48262\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48256\ : std_logic;
signal \N__48251\ : std_logic;
signal \N__48246\ : std_logic;
signal \N__48243\ : std_logic;
signal \N__48242\ : std_logic;
signal \N__48239\ : std_logic;
signal \N__48236\ : std_logic;
signal \N__48235\ : std_logic;
signal \N__48232\ : std_logic;
signal \N__48229\ : std_logic;
signal \N__48226\ : std_logic;
signal \N__48221\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48212\ : std_logic;
signal \N__48211\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48203\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48199\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48193\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48187\ : std_logic;
signal \N__48180\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48174\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48170\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48164\ : std_logic;
signal \N__48159\ : std_logic;
signal \N__48156\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48152\ : std_logic;
signal \N__48149\ : std_logic;
signal \N__48146\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48138\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48128\ : std_logic;
signal \N__48123\ : std_logic;
signal \N__48120\ : std_logic;
signal \N__48119\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48115\ : std_logic;
signal \N__48110\ : std_logic;
signal \N__48105\ : std_logic;
signal \N__48102\ : std_logic;
signal \N__48099\ : std_logic;
signal \N__48098\ : std_logic;
signal \N__48095\ : std_logic;
signal \N__48092\ : std_logic;
signal \N__48089\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48080\ : std_logic;
signal \N__48079\ : std_logic;
signal \N__48076\ : std_logic;
signal \N__48073\ : std_logic;
signal \N__48070\ : std_logic;
signal \N__48067\ : std_logic;
signal \N__48060\ : std_logic;
signal \N__48057\ : std_logic;
signal \N__48056\ : std_logic;
signal \N__48053\ : std_logic;
signal \N__48050\ : std_logic;
signal \N__48049\ : std_logic;
signal \N__48048\ : std_logic;
signal \N__48045\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48039\ : std_logic;
signal \N__48036\ : std_logic;
signal \N__48033\ : std_logic;
signal \N__48030\ : std_logic;
signal \N__48021\ : std_logic;
signal \N__48018\ : std_logic;
signal \N__48017\ : std_logic;
signal \N__48014\ : std_logic;
signal \N__48011\ : std_logic;
signal \N__48010\ : std_logic;
signal \N__48009\ : std_logic;
signal \N__48006\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__48000\ : std_logic;
signal \N__47997\ : std_logic;
signal \N__47994\ : std_logic;
signal \N__47991\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47979\ : std_logic;
signal \N__47978\ : std_logic;
signal \N__47977\ : std_logic;
signal \N__47974\ : std_logic;
signal \N__47971\ : std_logic;
signal \N__47968\ : std_logic;
signal \N__47967\ : std_logic;
signal \N__47964\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47958\ : std_logic;
signal \N__47955\ : std_logic;
signal \N__47950\ : std_logic;
signal \N__47943\ : std_logic;
signal \N__47940\ : std_logic;
signal \N__47937\ : std_logic;
signal \N__47934\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47928\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47919\ : std_logic;
signal \N__47916\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47910\ : std_logic;
signal \N__47907\ : std_logic;
signal \N__47904\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47892\ : std_logic;
signal \N__47889\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47883\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47877\ : std_logic;
signal \N__47874\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47864\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47858\ : std_logic;
signal \N__47855\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47838\ : std_logic;
signal \N__47837\ : std_logic;
signal \N__47832\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47826\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47820\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47808\ : std_logic;
signal \N__47805\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47793\ : std_logic;
signal \N__47790\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47786\ : std_logic;
signal \N__47783\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47766\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47760\ : std_logic;
signal \N__47757\ : std_logic;
signal \N__47754\ : std_logic;
signal \N__47751\ : std_logic;
signal \N__47748\ : std_logic;
signal \N__47745\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47739\ : std_logic;
signal \N__47738\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47727\ : std_logic;
signal \N__47724\ : std_logic;
signal \N__47721\ : std_logic;
signal \N__47718\ : std_logic;
signal \N__47715\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47711\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47707\ : std_logic;
signal \N__47704\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47698\ : std_logic;
signal \N__47695\ : std_logic;
signal \N__47692\ : std_logic;
signal \N__47689\ : std_logic;
signal \N__47682\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47675\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47658\ : std_logic;
signal \N__47655\ : std_logic;
signal \N__47652\ : std_logic;
signal \N__47649\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47647\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47638\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47628\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47619\ : std_logic;
signal \N__47616\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47595\ : std_logic;
signal \N__47592\ : std_logic;
signal \N__47589\ : std_logic;
signal \N__47586\ : std_logic;
signal \N__47583\ : std_logic;
signal \N__47580\ : std_logic;
signal \N__47579\ : std_logic;
signal \N__47576\ : std_logic;
signal \N__47573\ : std_logic;
signal \N__47572\ : std_logic;
signal \N__47569\ : std_logic;
signal \N__47566\ : std_logic;
signal \N__47563\ : std_logic;
signal \N__47556\ : std_logic;
signal \N__47553\ : std_logic;
signal \N__47550\ : std_logic;
signal \N__47547\ : std_logic;
signal \N__47544\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47536\ : std_logic;
signal \N__47533\ : std_logic;
signal \N__47530\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47514\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47505\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47486\ : std_logic;
signal \N__47483\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47475\ : std_logic;
signal \N__47472\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47466\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47454\ : std_logic;
signal \N__47451\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47445\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47433\ : std_logic;
signal \N__47430\ : std_logic;
signal \N__47427\ : std_logic;
signal \N__47424\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47415\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47409\ : std_logic;
signal \N__47406\ : std_logic;
signal \N__47405\ : std_logic;
signal \N__47402\ : std_logic;
signal \N__47401\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47392\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47382\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47373\ : std_logic;
signal \N__47370\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47362\ : std_logic;
signal \N__47359\ : std_logic;
signal \N__47356\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47335\ : std_logic;
signal \N__47332\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47321\ : std_logic;
signal \N__47318\ : std_logic;
signal \N__47315\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47309\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47283\ : std_logic;
signal \N__47280\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47276\ : std_logic;
signal \N__47273\ : std_logic;
signal \N__47270\ : std_logic;
signal \N__47267\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47259\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47245\ : std_logic;
signal \N__47242\ : std_logic;
signal \N__47239\ : std_logic;
signal \N__47236\ : std_logic;
signal \N__47229\ : std_logic;
signal \N__47226\ : std_logic;
signal \N__47223\ : std_logic;
signal \N__47220\ : std_logic;
signal \N__47217\ : std_logic;
signal \N__47214\ : std_logic;
signal \N__47211\ : std_logic;
signal \N__47208\ : std_logic;
signal \N__47207\ : std_logic;
signal \N__47204\ : std_logic;
signal \N__47201\ : std_logic;
signal \N__47200\ : std_logic;
signal \N__47197\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47184\ : std_logic;
signal \N__47181\ : std_logic;
signal \N__47180\ : std_logic;
signal \N__47177\ : std_logic;
signal \N__47174\ : std_logic;
signal \N__47173\ : std_logic;
signal \N__47170\ : std_logic;
signal \N__47167\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47157\ : std_logic;
signal \N__47154\ : std_logic;
signal \N__47151\ : std_logic;
signal \N__47148\ : std_logic;
signal \N__47145\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47141\ : std_logic;
signal \N__47138\ : std_logic;
signal \N__47135\ : std_logic;
signal \N__47132\ : std_logic;
signal \N__47129\ : std_logic;
signal \N__47126\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47118\ : std_logic;
signal \N__47117\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47109\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47103\ : std_logic;
signal \N__47100\ : std_logic;
signal \N__47097\ : std_logic;
signal \N__47094\ : std_logic;
signal \N__47091\ : std_logic;
signal \N__47088\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47082\ : std_logic;
signal \N__47081\ : std_logic;
signal \N__47078\ : std_logic;
signal \N__47075\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47064\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47060\ : std_logic;
signal \N__47057\ : std_logic;
signal \N__47056\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47050\ : std_logic;
signal \N__47047\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47031\ : std_logic;
signal \N__47028\ : std_logic;
signal \N__47025\ : std_logic;
signal \N__47022\ : std_logic;
signal \N__47019\ : std_logic;
signal \N__47016\ : std_logic;
signal \N__47013\ : std_logic;
signal \N__47010\ : std_logic;
signal \N__47007\ : std_logic;
signal \N__47006\ : std_logic;
signal \N__47005\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__47001\ : std_logic;
signal \N__47000\ : std_logic;
signal \N__46997\ : std_logic;
signal \N__46992\ : std_logic;
signal \N__46989\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46980\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46968\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46958\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46955\ : std_logic;
signal \N__46952\ : std_logic;
signal \N__46949\ : std_logic;
signal \N__46944\ : std_logic;
signal \N__46941\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46921\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46912\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46903\ : std_logic;
signal \N__46900\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46887\ : std_logic;
signal \N__46884\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46870\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46866\ : std_logic;
signal \N__46863\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46839\ : std_logic;
signal \N__46836\ : std_logic;
signal \N__46833\ : std_logic;
signal \N__46830\ : std_logic;
signal \N__46829\ : std_logic;
signal \N__46826\ : std_logic;
signal \N__46823\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46815\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46809\ : std_logic;
signal \N__46806\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46793\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46785\ : std_logic;
signal \N__46784\ : std_logic;
signal \N__46781\ : std_logic;
signal \N__46778\ : std_logic;
signal \N__46775\ : std_logic;
signal \N__46770\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46765\ : std_logic;
signal \N__46760\ : std_logic;
signal \N__46757\ : std_logic;
signal \N__46752\ : std_logic;
signal \N__46749\ : std_logic;
signal \N__46748\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46737\ : std_logic;
signal \N__46734\ : std_logic;
signal \N__46731\ : std_logic;
signal \N__46728\ : std_logic;
signal \N__46725\ : std_logic;
signal \N__46722\ : std_logic;
signal \N__46721\ : std_logic;
signal \N__46720\ : std_logic;
signal \N__46719\ : std_logic;
signal \N__46718\ : std_logic;
signal \N__46715\ : std_logic;
signal \N__46712\ : std_logic;
signal \N__46711\ : std_logic;
signal \N__46710\ : std_logic;
signal \N__46699\ : std_logic;
signal \N__46694\ : std_logic;
signal \N__46693\ : std_logic;
signal \N__46692\ : std_logic;
signal \N__46687\ : std_logic;
signal \N__46682\ : std_logic;
signal \N__46677\ : std_logic;
signal \N__46674\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46668\ : std_logic;
signal \N__46665\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46661\ : std_logic;
signal \N__46660\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46652\ : std_logic;
signal \N__46649\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46633\ : std_logic;
signal \N__46630\ : std_logic;
signal \N__46623\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46616\ : std_logic;
signal \N__46615\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46602\ : std_logic;
signal \N__46601\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46591\ : std_logic;
signal \N__46588\ : std_logic;
signal \N__46583\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46575\ : std_logic;
signal \N__46572\ : std_logic;
signal \N__46571\ : std_logic;
signal \N__46568\ : std_logic;
signal \N__46565\ : std_logic;
signal \N__46562\ : std_logic;
signal \N__46559\ : std_logic;
signal \N__46556\ : std_logic;
signal \N__46553\ : std_logic;
signal \N__46548\ : std_logic;
signal \N__46547\ : std_logic;
signal \N__46544\ : std_logic;
signal \N__46541\ : std_logic;
signal \N__46540\ : std_logic;
signal \N__46535\ : std_logic;
signal \N__46532\ : std_logic;
signal \N__46527\ : std_logic;
signal \N__46526\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46506\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46499\ : std_logic;
signal \N__46496\ : std_logic;
signal \N__46493\ : std_logic;
signal \N__46490\ : std_logic;
signal \N__46485\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46479\ : std_logic;
signal \N__46476\ : std_logic;
signal \N__46475\ : std_logic;
signal \N__46470\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46464\ : std_logic;
signal \N__46461\ : std_logic;
signal \N__46458\ : std_logic;
signal \N__46457\ : std_logic;
signal \N__46456\ : std_logic;
signal \N__46453\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46442\ : std_logic;
signal \N__46439\ : std_logic;
signal \N__46434\ : std_logic;
signal \N__46431\ : std_logic;
signal \N__46428\ : std_logic;
signal \N__46425\ : std_logic;
signal \N__46424\ : std_logic;
signal \N__46421\ : std_logic;
signal \N__46418\ : std_logic;
signal \N__46417\ : std_logic;
signal \N__46412\ : std_logic;
signal \N__46409\ : std_logic;
signal \N__46406\ : std_logic;
signal \N__46401\ : std_logic;
signal \N__46400\ : std_logic;
signal \N__46397\ : std_logic;
signal \N__46396\ : std_logic;
signal \N__46395\ : std_logic;
signal \N__46394\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46390\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46377\ : std_logic;
signal \N__46372\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46361\ : std_logic;
signal \N__46356\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46350\ : std_logic;
signal \N__46347\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46340\ : std_logic;
signal \N__46337\ : std_logic;
signal \N__46334\ : std_logic;
signal \N__46333\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46327\ : std_logic;
signal \N__46322\ : std_logic;
signal \N__46319\ : std_logic;
signal \N__46316\ : std_logic;
signal \N__46313\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46307\ : std_logic;
signal \N__46306\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46300\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46291\ : std_logic;
signal \N__46288\ : std_logic;
signal \N__46281\ : std_logic;
signal \N__46278\ : std_logic;
signal \N__46277\ : std_logic;
signal \N__46274\ : std_logic;
signal \N__46271\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46266\ : std_logic;
signal \N__46263\ : std_logic;
signal \N__46260\ : std_logic;
signal \N__46257\ : std_logic;
signal \N__46254\ : std_logic;
signal \N__46251\ : std_logic;
signal \N__46248\ : std_logic;
signal \N__46239\ : std_logic;
signal \N__46236\ : std_logic;
signal \N__46233\ : std_logic;
signal \N__46230\ : std_logic;
signal \N__46227\ : std_logic;
signal \N__46224\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46218\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46212\ : std_logic;
signal \N__46209\ : std_logic;
signal \N__46208\ : std_logic;
signal \N__46205\ : std_logic;
signal \N__46202\ : std_logic;
signal \N__46197\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46188\ : std_logic;
signal \N__46185\ : std_logic;
signal \N__46184\ : std_logic;
signal \N__46179\ : std_logic;
signal \N__46176\ : std_logic;
signal \N__46173\ : std_logic;
signal \N__46170\ : std_logic;
signal \N__46167\ : std_logic;
signal \N__46164\ : std_logic;
signal \N__46161\ : std_logic;
signal \N__46158\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46142\ : std_logic;
signal \N__46139\ : std_logic;
signal \N__46136\ : std_logic;
signal \N__46131\ : std_logic;
signal \N__46128\ : std_logic;
signal \N__46125\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46110\ : std_logic;
signal \N__46107\ : std_logic;
signal \N__46104\ : std_logic;
signal \N__46101\ : std_logic;
signal \N__46100\ : std_logic;
signal \N__46097\ : std_logic;
signal \N__46096\ : std_logic;
signal \N__46093\ : std_logic;
signal \N__46090\ : std_logic;
signal \N__46087\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46068\ : std_logic;
signal \N__46065\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46061\ : std_logic;
signal \N__46058\ : std_logic;
signal \N__46055\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46044\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46033\ : std_logic;
signal \N__46028\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46013\ : std_logic;
signal \N__46012\ : std_logic;
signal \N__46009\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__46003\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45984\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45972\ : std_logic;
signal \N__45969\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45962\ : std_logic;
signal \N__45957\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45951\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45939\ : std_logic;
signal \N__45936\ : std_logic;
signal \N__45933\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45924\ : std_logic;
signal \N__45923\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45917\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45909\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45899\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45893\ : std_logic;
signal \N__45888\ : std_logic;
signal \N__45885\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45879\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45872\ : std_logic;
signal \N__45869\ : std_logic;
signal \N__45864\ : std_logic;
signal \N__45861\ : std_logic;
signal \N__45858\ : std_logic;
signal \N__45855\ : std_logic;
signal \N__45854\ : std_logic;
signal \N__45851\ : std_logic;
signal \N__45850\ : std_logic;
signal \N__45847\ : std_logic;
signal \N__45844\ : std_logic;
signal \N__45841\ : std_logic;
signal \N__45834\ : std_logic;
signal \N__45831\ : std_logic;
signal \N__45828\ : std_logic;
signal \N__45825\ : std_logic;
signal \N__45822\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45816\ : std_logic;
signal \N__45813\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45800\ : std_logic;
signal \N__45799\ : std_logic;
signal \N__45796\ : std_logic;
signal \N__45793\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45784\ : std_logic;
signal \N__45781\ : std_logic;
signal \N__45776\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45758\ : std_logic;
signal \N__45757\ : std_logic;
signal \N__45754\ : std_logic;
signal \N__45751\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45743\ : std_logic;
signal \N__45740\ : std_logic;
signal \N__45737\ : std_logic;
signal \N__45732\ : std_logic;
signal \N__45729\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45723\ : std_logic;
signal \N__45720\ : std_logic;
signal \N__45717\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45702\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45689\ : std_logic;
signal \N__45684\ : std_logic;
signal \N__45681\ : std_logic;
signal \N__45678\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45670\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45664\ : std_logic;
signal \N__45661\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45648\ : std_logic;
signal \N__45645\ : std_logic;
signal \N__45642\ : std_logic;
signal \N__45639\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45633\ : std_logic;
signal \N__45630\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45624\ : std_logic;
signal \N__45621\ : std_logic;
signal \N__45618\ : std_logic;
signal \N__45617\ : std_logic;
signal \N__45616\ : std_logic;
signal \N__45615\ : std_logic;
signal \N__45614\ : std_logic;
signal \N__45613\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45609\ : std_logic;
signal \N__45608\ : std_logic;
signal \N__45605\ : std_logic;
signal \N__45604\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45602\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45598\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45594\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45588\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45586\ : std_logic;
signal \N__45583\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45559\ : std_logic;
signal \N__45550\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45506\ : std_logic;
signal \N__45503\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45500\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45490\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45486\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45484\ : std_logic;
signal \N__45481\ : std_logic;
signal \N__45480\ : std_logic;
signal \N__45477\ : std_logic;
signal \N__45476\ : std_logic;
signal \N__45473\ : std_logic;
signal \N__45468\ : std_logic;
signal \N__45465\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45457\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45417\ : std_logic;
signal \N__45410\ : std_logic;
signal \N__45399\ : std_logic;
signal \N__45396\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45389\ : std_logic;
signal \N__45386\ : std_logic;
signal \N__45383\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45372\ : std_logic;
signal \N__45371\ : std_logic;
signal \N__45368\ : std_logic;
signal \N__45365\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45358\ : std_logic;
signal \N__45355\ : std_logic;
signal \N__45348\ : std_logic;
signal \N__45345\ : std_logic;
signal \N__45342\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45335\ : std_logic;
signal \N__45332\ : std_logic;
signal \N__45329\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45314\ : std_logic;
signal \N__45311\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45307\ : std_logic;
signal \N__45304\ : std_logic;
signal \N__45301\ : std_logic;
signal \N__45294\ : std_logic;
signal \N__45291\ : std_logic;
signal \N__45288\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45282\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45278\ : std_logic;
signal \N__45277\ : std_logic;
signal \N__45274\ : std_logic;
signal \N__45269\ : std_logic;
signal \N__45264\ : std_logic;
signal \N__45261\ : std_logic;
signal \N__45258\ : std_logic;
signal \N__45255\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45249\ : std_logic;
signal \N__45246\ : std_logic;
signal \N__45245\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45239\ : std_logic;
signal \N__45236\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45229\ : std_logic;
signal \N__45226\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45216\ : std_logic;
signal \N__45213\ : std_logic;
signal \N__45210\ : std_logic;
signal \N__45209\ : std_logic;
signal \N__45206\ : std_logic;
signal \N__45203\ : std_logic;
signal \N__45200\ : std_logic;
signal \N__45197\ : std_logic;
signal \N__45196\ : std_logic;
signal \N__45193\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45171\ : std_logic;
signal \N__45168\ : std_logic;
signal \N__45167\ : std_logic;
signal \N__45164\ : std_logic;
signal \N__45161\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45152\ : std_logic;
signal \N__45149\ : std_logic;
signal \N__45146\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45129\ : std_logic;
signal \N__45126\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45111\ : std_logic;
signal \N__45108\ : std_logic;
signal \N__45105\ : std_logic;
signal \N__45102\ : std_logic;
signal \N__45099\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45093\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45084\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45059\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45050\ : std_logic;
signal \N__45049\ : std_logic;
signal \N__45046\ : std_logic;
signal \N__45039\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45030\ : std_logic;
signal \N__45027\ : std_logic;
signal \N__45024\ : std_logic;
signal \N__45021\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45000\ : std_logic;
signal \N__44997\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44988\ : std_logic;
signal \N__44985\ : std_logic;
signal \N__44982\ : std_logic;
signal \N__44979\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44970\ : std_logic;
signal \N__44967\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44958\ : std_logic;
signal \N__44955\ : std_logic;
signal \N__44954\ : std_logic;
signal \N__44951\ : std_logic;
signal \N__44948\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44910\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44904\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44892\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44880\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44875\ : std_logic;
signal \N__44870\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44856\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44850\ : std_logic;
signal \N__44847\ : std_logic;
signal \N__44844\ : std_logic;
signal \N__44841\ : std_logic;
signal \N__44838\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44829\ : std_logic;
signal \N__44826\ : std_logic;
signal \N__44823\ : std_logic;
signal \N__44820\ : std_logic;
signal \N__44819\ : std_logic;
signal \N__44816\ : std_logic;
signal \N__44813\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44807\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44796\ : std_logic;
signal \N__44793\ : std_logic;
signal \N__44790\ : std_logic;
signal \N__44789\ : std_logic;
signal \N__44788\ : std_logic;
signal \N__44785\ : std_logic;
signal \N__44782\ : std_logic;
signal \N__44779\ : std_logic;
signal \N__44774\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44766\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44747\ : std_logic;
signal \N__44744\ : std_logic;
signal \N__44741\ : std_logic;
signal \N__44738\ : std_logic;
signal \N__44733\ : std_logic;
signal \N__44732\ : std_logic;
signal \N__44729\ : std_logic;
signal \N__44726\ : std_logic;
signal \N__44721\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44711\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44700\ : std_logic;
signal \N__44697\ : std_logic;
signal \N__44696\ : std_logic;
signal \N__44691\ : std_logic;
signal \N__44688\ : std_logic;
signal \N__44685\ : std_logic;
signal \N__44682\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44678\ : std_logic;
signal \N__44677\ : std_logic;
signal \N__44674\ : std_logic;
signal \N__44669\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44658\ : std_logic;
signal \N__44655\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44643\ : std_logic;
signal \N__44640\ : std_logic;
signal \N__44639\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44633\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44622\ : std_logic;
signal \N__44619\ : std_logic;
signal \N__44618\ : std_logic;
signal \N__44613\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44604\ : std_logic;
signal \N__44601\ : std_logic;
signal \N__44598\ : std_logic;
signal \N__44595\ : std_logic;
signal \N__44592\ : std_logic;
signal \N__44591\ : std_logic;
signal \N__44588\ : std_logic;
signal \N__44585\ : std_logic;
signal \N__44580\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44574\ : std_logic;
signal \N__44571\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44559\ : std_logic;
signal \N__44556\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44550\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44544\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44537\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44529\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44514\ : std_logic;
signal \N__44511\ : std_logic;
signal \N__44508\ : std_logic;
signal \N__44505\ : std_logic;
signal \N__44502\ : std_logic;
signal \N__44501\ : std_logic;
signal \N__44498\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44490\ : std_logic;
signal \N__44487\ : std_logic;
signal \N__44484\ : std_logic;
signal \N__44483\ : std_logic;
signal \N__44478\ : std_logic;
signal \N__44475\ : std_logic;
signal \N__44472\ : std_logic;
signal \N__44469\ : std_logic;
signal \N__44466\ : std_logic;
signal \N__44463\ : std_logic;
signal \N__44460\ : std_logic;
signal \N__44457\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44451\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44447\ : std_logic;
signal \N__44444\ : std_logic;
signal \N__44439\ : std_logic;
signal \N__44436\ : std_logic;
signal \N__44433\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44424\ : std_logic;
signal \N__44421\ : std_logic;
signal \N__44418\ : std_logic;
signal \N__44415\ : std_logic;
signal \N__44412\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44397\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44391\ : std_logic;
signal \N__44388\ : std_logic;
signal \N__44385\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44370\ : std_logic;
signal \N__44367\ : std_logic;
signal \N__44364\ : std_logic;
signal \N__44361\ : std_logic;
signal \N__44358\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44343\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44337\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44322\ : std_logic;
signal \N__44319\ : std_logic;
signal \N__44316\ : std_logic;
signal \N__44313\ : std_logic;
signal \N__44310\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44306\ : std_logic;
signal \N__44303\ : std_logic;
signal \N__44300\ : std_logic;
signal \N__44297\ : std_logic;
signal \N__44294\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44277\ : std_logic;
signal \N__44274\ : std_logic;
signal \N__44271\ : std_logic;
signal \N__44270\ : std_logic;
signal \N__44267\ : std_logic;
signal \N__44264\ : std_logic;
signal \N__44261\ : std_logic;
signal \N__44258\ : std_logic;
signal \N__44255\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44235\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44231\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44222\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44214\ : std_logic;
signal \N__44211\ : std_logic;
signal \N__44208\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44202\ : std_logic;
signal \N__44201\ : std_logic;
signal \N__44198\ : std_logic;
signal \N__44195\ : std_logic;
signal \N__44192\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44186\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44175\ : std_logic;
signal \N__44172\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44166\ : std_logic;
signal \N__44163\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44154\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44150\ : std_logic;
signal \N__44147\ : std_logic;
signal \N__44144\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44130\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44120\ : std_logic;
signal \N__44117\ : std_logic;
signal \N__44114\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44097\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44093\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44090\ : std_logic;
signal \N__44089\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44076\ : std_logic;
signal \N__44073\ : std_logic;
signal \N__44064\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44057\ : std_logic;
signal \N__44054\ : std_logic;
signal \N__44051\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44043\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44019\ : std_logic;
signal \N__44016\ : std_logic;
signal \N__44013\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43992\ : std_logic;
signal \N__43991\ : std_logic;
signal \N__43988\ : std_logic;
signal \N__43985\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43977\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43971\ : std_logic;
signal \N__43968\ : std_logic;
signal \N__43965\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43958\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43952\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43941\ : std_logic;
signal \N__43938\ : std_logic;
signal \N__43935\ : std_logic;
signal \N__43932\ : std_logic;
signal \N__43929\ : std_logic;
signal \N__43926\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43917\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43913\ : std_logic;
signal \N__43910\ : std_logic;
signal \N__43909\ : std_logic;
signal \N__43906\ : std_logic;
signal \N__43903\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43897\ : std_logic;
signal \N__43894\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43884\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43874\ : std_logic;
signal \N__43871\ : std_logic;
signal \N__43868\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43860\ : std_logic;
signal \N__43857\ : std_logic;
signal \N__43854\ : std_logic;
signal \N__43851\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43839\ : std_logic;
signal \N__43838\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43814\ : std_logic;
signal \N__43809\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43802\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43795\ : std_logic;
signal \N__43792\ : std_logic;
signal \N__43787\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43779\ : std_logic;
signal \N__43776\ : std_logic;
signal \N__43773\ : std_logic;
signal \N__43770\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43764\ : std_logic;
signal \N__43761\ : std_logic;
signal \N__43758\ : std_logic;
signal \N__43755\ : std_logic;
signal \N__43752\ : std_logic;
signal \N__43749\ : std_logic;
signal \N__43748\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43742\ : std_logic;
signal \N__43739\ : std_logic;
signal \N__43736\ : std_logic;
signal \N__43735\ : std_logic;
signal \N__43730\ : std_logic;
signal \N__43727\ : std_logic;
signal \N__43724\ : std_logic;
signal \N__43719\ : std_logic;
signal \N__43716\ : std_logic;
signal \N__43713\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43698\ : std_logic;
signal \N__43695\ : std_logic;
signal \N__43692\ : std_logic;
signal \N__43689\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43684\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43671\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43665\ : std_logic;
signal \N__43662\ : std_logic;
signal \N__43659\ : std_logic;
signal \N__43656\ : std_logic;
signal \N__43655\ : std_logic;
signal \N__43652\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43639\ : std_logic;
signal \N__43634\ : std_logic;
signal \N__43631\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43623\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43610\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43604\ : std_logic;
signal \N__43599\ : std_logic;
signal \N__43596\ : std_logic;
signal \N__43593\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43557\ : std_logic;
signal \N__43554\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43530\ : std_logic;
signal \N__43527\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43512\ : std_logic;
signal \N__43509\ : std_logic;
signal \N__43506\ : std_logic;
signal \N__43503\ : std_logic;
signal \N__43500\ : std_logic;
signal \N__43497\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43487\ : std_logic;
signal \N__43484\ : std_logic;
signal \N__43483\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43477\ : std_logic;
signal \N__43474\ : std_logic;
signal \N__43467\ : std_logic;
signal \N__43464\ : std_logic;
signal \N__43461\ : std_logic;
signal \N__43458\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43437\ : std_logic;
signal \N__43434\ : std_logic;
signal \N__43431\ : std_logic;
signal \N__43428\ : std_logic;
signal \N__43425\ : std_logic;
signal \N__43422\ : std_logic;
signal \N__43419\ : std_logic;
signal \N__43418\ : std_logic;
signal \N__43415\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43407\ : std_logic;
signal \N__43404\ : std_logic;
signal \N__43401\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43391\ : std_logic;
signal \N__43390\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43368\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43356\ : std_logic;
signal \N__43353\ : std_logic;
signal \N__43350\ : std_logic;
signal \N__43347\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43338\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43332\ : std_logic;
signal \N__43329\ : std_logic;
signal \N__43326\ : std_logic;
signal \N__43323\ : std_logic;
signal \N__43320\ : std_logic;
signal \N__43317\ : std_logic;
signal \N__43314\ : std_logic;
signal \N__43311\ : std_logic;
signal \N__43310\ : std_logic;
signal \N__43307\ : std_logic;
signal \N__43304\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43297\ : std_logic;
signal \N__43294\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43278\ : std_logic;
signal \N__43275\ : std_logic;
signal \N__43272\ : std_logic;
signal \N__43271\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43262\ : std_logic;
signal \N__43259\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43251\ : std_logic;
signal \N__43248\ : std_logic;
signal \N__43245\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43224\ : std_logic;
signal \N__43221\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43215\ : std_logic;
signal \N__43212\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43203\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43197\ : std_logic;
signal \N__43194\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43169\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43162\ : std_logic;
signal \N__43159\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43142\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43135\ : std_logic;
signal \N__43132\ : std_logic;
signal \N__43129\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43116\ : std_logic;
signal \N__43113\ : std_logic;
signal \N__43112\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43105\ : std_logic;
signal \N__43102\ : std_logic;
signal \N__43099\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43086\ : std_logic;
signal \N__43083\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43075\ : std_logic;
signal \N__43072\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43058\ : std_logic;
signal \N__43057\ : std_logic;
signal \N__43054\ : std_logic;
signal \N__43051\ : std_logic;
signal \N__43046\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43040\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43032\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43028\ : std_logic;
signal \N__43027\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43015\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43005\ : std_logic;
signal \N__43002\ : std_logic;
signal \N__42999\ : std_logic;
signal \N__42996\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42990\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42980\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42972\ : std_logic;
signal \N__42969\ : std_logic;
signal \N__42966\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42964\ : std_logic;
signal \N__42961\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42955\ : std_logic;
signal \N__42952\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42942\ : std_logic;
signal \N__42939\ : std_logic;
signal \N__42936\ : std_logic;
signal \N__42933\ : std_logic;
signal \N__42930\ : std_logic;
signal \N__42929\ : std_logic;
signal \N__42926\ : std_logic;
signal \N__42923\ : std_logic;
signal \N__42920\ : std_logic;
signal \N__42917\ : std_logic;
signal \N__42914\ : std_logic;
signal \N__42911\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42903\ : std_logic;
signal \N__42900\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42896\ : std_logic;
signal \N__42891\ : std_logic;
signal \N__42888\ : std_logic;
signal \N__42885\ : std_logic;
signal \N__42882\ : std_logic;
signal \N__42879\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42875\ : std_logic;
signal \N__42872\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42861\ : std_logic;
signal \N__42858\ : std_logic;
signal \N__42855\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42845\ : std_logic;
signal \N__42842\ : std_logic;
signal \N__42841\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42825\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42783\ : std_logic;
signal \N__42780\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42774\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42756\ : std_logic;
signal \N__42753\ : std_logic;
signal \N__42750\ : std_logic;
signal \N__42747\ : std_logic;
signal \N__42744\ : std_logic;
signal \N__42741\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42735\ : std_logic;
signal \N__42732\ : std_logic;
signal \N__42729\ : std_logic;
signal \N__42726\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42714\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42704\ : std_logic;
signal \N__42703\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42693\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42678\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42669\ : std_logic;
signal \N__42666\ : std_logic;
signal \N__42663\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42651\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42642\ : std_logic;
signal \N__42639\ : std_logic;
signal \N__42636\ : std_logic;
signal \N__42633\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42609\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42597\ : std_logic;
signal \N__42594\ : std_logic;
signal \N__42591\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42582\ : std_logic;
signal \N__42579\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42573\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42534\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42528\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42501\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42492\ : std_logic;
signal \N__42489\ : std_logic;
signal \N__42486\ : std_logic;
signal \N__42483\ : std_logic;
signal \N__42480\ : std_logic;
signal \N__42477\ : std_logic;
signal \N__42474\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42441\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42427\ : std_logic;
signal \N__42424\ : std_logic;
signal \N__42421\ : std_logic;
signal \N__42418\ : std_logic;
signal \N__42415\ : std_logic;
signal \N__42410\ : std_logic;
signal \N__42407\ : std_logic;
signal \N__42404\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42378\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42371\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42348\ : std_logic;
signal \N__42347\ : std_logic;
signal \N__42344\ : std_logic;
signal \N__42341\ : std_logic;
signal \N__42340\ : std_logic;
signal \N__42337\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42323\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42316\ : std_logic;
signal \N__42313\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42307\ : std_logic;
signal \N__42304\ : std_logic;
signal \N__42301\ : std_logic;
signal \N__42298\ : std_logic;
signal \N__42295\ : std_logic;
signal \N__42292\ : std_logic;
signal \N__42289\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42278\ : std_logic;
signal \N__42275\ : std_logic;
signal \N__42272\ : std_logic;
signal \N__42269\ : std_logic;
signal \N__42264\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42257\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42244\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42238\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42228\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42201\ : std_logic;
signal \N__42198\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42193\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42185\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42175\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42159\ : std_logic;
signal \N__42156\ : std_logic;
signal \N__42155\ : std_logic;
signal \N__42152\ : std_logic;
signal \N__42151\ : std_logic;
signal \N__42148\ : std_logic;
signal \N__42145\ : std_logic;
signal \N__42142\ : std_logic;
signal \N__42135\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42118\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42099\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42074\ : std_logic;
signal \N__42073\ : std_logic;
signal \N__42070\ : std_logic;
signal \N__42067\ : std_logic;
signal \N__42064\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42036\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42030\ : std_logic;
signal \N__42027\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42020\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42016\ : std_logic;
signal \N__42013\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41995\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41970\ : std_logic;
signal \N__41967\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41954\ : std_logic;
signal \N__41951\ : std_logic;
signal \N__41950\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41922\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41918\ : std_logic;
signal \N__41917\ : std_logic;
signal \N__41914\ : std_logic;
signal \N__41909\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41898\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41871\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41865\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41859\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41846\ : std_logic;
signal \N__41843\ : std_logic;
signal \N__41840\ : std_logic;
signal \N__41835\ : std_logic;
signal \N__41832\ : std_logic;
signal \N__41829\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41818\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41814\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41796\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41787\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41784\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41767\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41757\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41748\ : std_logic;
signal \N__41745\ : std_logic;
signal \N__41744\ : std_logic;
signal \N__41741\ : std_logic;
signal \N__41738\ : std_logic;
signal \N__41735\ : std_logic;
signal \N__41732\ : std_logic;
signal \N__41729\ : std_logic;
signal \N__41726\ : std_logic;
signal \N__41725\ : std_logic;
signal \N__41720\ : std_logic;
signal \N__41717\ : std_logic;
signal \N__41712\ : std_logic;
signal \N__41709\ : std_logic;
signal \N__41706\ : std_logic;
signal \N__41703\ : std_logic;
signal \N__41702\ : std_logic;
signal \N__41699\ : std_logic;
signal \N__41696\ : std_logic;
signal \N__41693\ : std_logic;
signal \N__41690\ : std_logic;
signal \N__41687\ : std_logic;
signal \N__41684\ : std_logic;
signal \N__41683\ : std_logic;
signal \N__41680\ : std_logic;
signal \N__41677\ : std_logic;
signal \N__41674\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41666\ : std_logic;
signal \N__41665\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41654\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41637\ : std_logic;
signal \N__41636\ : std_logic;
signal \N__41633\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41627\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41621\ : std_logic;
signal \N__41618\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41610\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41600\ : std_logic;
signal \N__41597\ : std_logic;
signal \N__41596\ : std_logic;
signal \N__41593\ : std_logic;
signal \N__41590\ : std_logic;
signal \N__41587\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41581\ : std_logic;
signal \N__41578\ : std_logic;
signal \N__41571\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41563\ : std_logic;
signal \N__41560\ : std_logic;
signal \N__41557\ : std_logic;
signal \N__41554\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41532\ : std_logic;
signal \N__41529\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41520\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41516\ : std_logic;
signal \N__41515\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41513\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41509\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41505\ : std_logic;
signal \N__41504\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41502\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41491\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41489\ : std_logic;
signal \N__41486\ : std_logic;
signal \N__41483\ : std_logic;
signal \N__41482\ : std_logic;
signal \N__41477\ : std_logic;
signal \N__41472\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41455\ : std_logic;
signal \N__41446\ : std_logic;
signal \N__41439\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41421\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41411\ : std_logic;
signal \N__41408\ : std_logic;
signal \N__41405\ : std_logic;
signal \N__41402\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41394\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41388\ : std_logic;
signal \N__41385\ : std_logic;
signal \N__41382\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41374\ : std_logic;
signal \N__41371\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41369\ : std_logic;
signal \N__41368\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41359\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41344\ : std_logic;
signal \N__41343\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41341\ : std_logic;
signal \N__41340\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41334\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41317\ : std_logic;
signal \N__41314\ : std_logic;
signal \N__41311\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41289\ : std_logic;
signal \N__41274\ : std_logic;
signal \N__41273\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41260\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41254\ : std_logic;
signal \N__41251\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41240\ : std_logic;
signal \N__41237\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41228\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41209\ : std_logic;
signal \N__41206\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41200\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41187\ : std_logic;
signal \N__41184\ : std_logic;
signal \N__41181\ : std_logic;
signal \N__41178\ : std_logic;
signal \N__41175\ : std_logic;
signal \N__41172\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41154\ : std_logic;
signal \N__41151\ : std_logic;
signal \N__41148\ : std_logic;
signal \N__41145\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41126\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41117\ : std_logic;
signal \N__41114\ : std_logic;
signal \N__41111\ : std_logic;
signal \N__41106\ : std_logic;
signal \N__41103\ : std_logic;
signal \N__41100\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41091\ : std_logic;
signal \N__41088\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41075\ : std_logic;
signal \N__41070\ : std_logic;
signal \N__41067\ : std_logic;
signal \N__41064\ : std_logic;
signal \N__41061\ : std_logic;
signal \N__41058\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41043\ : std_logic;
signal \N__41040\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41034\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41016\ : std_logic;
signal \N__41013\ : std_logic;
signal \N__41010\ : std_logic;
signal \N__41007\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40990\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40977\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40967\ : std_logic;
signal \N__40964\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40953\ : std_logic;
signal \N__40950\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40948\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40939\ : std_logic;
signal \N__40934\ : std_logic;
signal \N__40931\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40920\ : std_logic;
signal \N__40917\ : std_logic;
signal \N__40914\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40910\ : std_logic;
signal \N__40907\ : std_logic;
signal \N__40904\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40898\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40890\ : std_logic;
signal \N__40887\ : std_logic;
signal \N__40884\ : std_logic;
signal \N__40883\ : std_logic;
signal \N__40880\ : std_logic;
signal \N__40879\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40873\ : std_logic;
signal \N__40870\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40848\ : std_logic;
signal \N__40847\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40841\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40833\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40818\ : std_logic;
signal \N__40815\ : std_logic;
signal \N__40812\ : std_logic;
signal \N__40809\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40797\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40791\ : std_logic;
signal \N__40788\ : std_logic;
signal \N__40785\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40781\ : std_logic;
signal \N__40780\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40772\ : std_logic;
signal \N__40767\ : std_logic;
signal \N__40764\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40762\ : std_logic;
signal \N__40757\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40749\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40743\ : std_logic;
signal \N__40742\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40736\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40719\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40713\ : std_logic;
signal \N__40710\ : std_logic;
signal \N__40707\ : std_logic;
signal \N__40704\ : std_logic;
signal \N__40701\ : std_logic;
signal \N__40698\ : std_logic;
signal \N__40695\ : std_logic;
signal \N__40692\ : std_logic;
signal \N__40689\ : std_logic;
signal \N__40686\ : std_logic;
signal \N__40683\ : std_logic;
signal \N__40680\ : std_logic;
signal \N__40677\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40668\ : std_logic;
signal \N__40665\ : std_logic;
signal \N__40662\ : std_logic;
signal \N__40659\ : std_logic;
signal \N__40656\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40650\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40635\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40608\ : std_logic;
signal \N__40605\ : std_logic;
signal \N__40602\ : std_logic;
signal \N__40599\ : std_logic;
signal \N__40596\ : std_logic;
signal \N__40593\ : std_logic;
signal \N__40590\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40584\ : std_logic;
signal \N__40581\ : std_logic;
signal \N__40578\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40572\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40566\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40559\ : std_logic;
signal \N__40556\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40548\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40542\ : std_logic;
signal \N__40541\ : std_logic;
signal \N__40538\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40526\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40523\ : std_logic;
signal \N__40522\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40517\ : std_logic;
signal \N__40516\ : std_logic;
signal \N__40515\ : std_logic;
signal \N__40514\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40508\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40504\ : std_logic;
signal \N__40501\ : std_logic;
signal \N__40500\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40496\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40492\ : std_logic;
signal \N__40489\ : std_logic;
signal \N__40488\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40484\ : std_logic;
signal \N__40481\ : std_logic;
signal \N__40480\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40473\ : std_logic;
signal \N__40472\ : std_logic;
signal \N__40469\ : std_logic;
signal \N__40468\ : std_logic;
signal \N__40467\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40460\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40438\ : std_logic;
signal \N__40421\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40389\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40371\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40356\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40350\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40344\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40338\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40311\ : std_logic;
signal \N__40308\ : std_logic;
signal \N__40305\ : std_logic;
signal \N__40304\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40290\ : std_logic;
signal \N__40287\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40272\ : std_logic;
signal \N__40267\ : std_logic;
signal \N__40260\ : std_logic;
signal \N__40257\ : std_logic;
signal \N__40254\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40245\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40236\ : std_logic;
signal \N__40233\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40231\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40228\ : std_logic;
signal \N__40227\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40225\ : std_logic;
signal \N__40224\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40222\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40217\ : std_logic;
signal \N__40214\ : std_logic;
signal \N__40211\ : std_logic;
signal \N__40210\ : std_logic;
signal \N__40207\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40191\ : std_logic;
signal \N__40188\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40174\ : std_logic;
signal \N__40173\ : std_logic;
signal \N__40172\ : std_logic;
signal \N__40171\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40169\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40102\ : std_logic;
signal \N__40095\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40083\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40065\ : std_logic;
signal \N__40062\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40056\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40050\ : std_logic;
signal \N__40047\ : std_logic;
signal \N__40044\ : std_logic;
signal \N__40041\ : std_logic;
signal \N__40038\ : std_logic;
signal \N__40035\ : std_logic;
signal \N__40032\ : std_logic;
signal \N__40029\ : std_logic;
signal \N__40026\ : std_logic;
signal \N__40023\ : std_logic;
signal \N__40020\ : std_logic;
signal \N__40017\ : std_logic;
signal \N__40014\ : std_logic;
signal \N__40011\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39997\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39978\ : std_logic;
signal \N__39975\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39970\ : std_logic;
signal \N__39967\ : std_logic;
signal \N__39964\ : std_logic;
signal \N__39961\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39955\ : std_logic;
signal \N__39952\ : std_logic;
signal \N__39949\ : std_logic;
signal \N__39946\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39936\ : std_logic;
signal \N__39933\ : std_logic;
signal \N__39930\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39928\ : std_logic;
signal \N__39925\ : std_logic;
signal \N__39922\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39916\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39906\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39885\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39858\ : std_logic;
signal \N__39855\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39846\ : std_logic;
signal \N__39843\ : std_logic;
signal \N__39840\ : std_logic;
signal \N__39837\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39831\ : std_logic;
signal \N__39828\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39826\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39810\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39790\ : std_logic;
signal \N__39787\ : std_logic;
signal \N__39780\ : std_logic;
signal \N__39777\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39764\ : std_logic;
signal \N__39761\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39748\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39731\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39718\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39709\ : std_logic;
signal \N__39702\ : std_logic;
signal \N__39699\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39692\ : std_logic;
signal \N__39691\ : std_logic;
signal \N__39688\ : std_logic;
signal \N__39685\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39675\ : std_logic;
signal \N__39672\ : std_logic;
signal \N__39671\ : std_logic;
signal \N__39668\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39664\ : std_logic;
signal \N__39661\ : std_logic;
signal \N__39658\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39639\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39633\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39622\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39609\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39602\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39592\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39575\ : std_logic;
signal \N__39572\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39562\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39506\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39502\ : std_logic;
signal \N__39499\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39490\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39473\ : std_logic;
signal \N__39470\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39460\ : std_logic;
signal \N__39453\ : std_logic;
signal \N__39450\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39439\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39430\ : std_logic;
signal \N__39427\ : std_logic;
signal \N__39424\ : std_logic;
signal \N__39417\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39373\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39367\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39353\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39340\ : std_logic;
signal \N__39337\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39320\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39295\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39281\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39277\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39271\ : std_logic;
signal \N__39268\ : std_logic;
signal \N__39265\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39246\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39242\ : std_logic;
signal \N__39239\ : std_logic;
signal \N__39236\ : std_logic;
signal \N__39233\ : std_logic;
signal \N__39230\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39224\ : std_logic;
signal \N__39221\ : std_logic;
signal \N__39218\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39211\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39187\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39185\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39182\ : std_logic;
signal \N__39181\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39141\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39126\ : std_logic;
signal \N__39123\ : std_logic;
signal \N__39122\ : std_logic;
signal \N__39119\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39106\ : std_logic;
signal \N__39103\ : std_logic;
signal \N__39100\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39054\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39043\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39025\ : std_logic;
signal \N__39022\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39009\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39003\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38974\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38966\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38950\ : std_logic;
signal \N__38947\ : std_logic;
signal \N__38942\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38907\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38898\ : std_logic;
signal \N__38895\ : std_logic;
signal \N__38892\ : std_logic;
signal \N__38889\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38885\ : std_logic;
signal \N__38882\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38864\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38857\ : std_logic;
signal \N__38854\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38841\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38795\ : std_logic;
signal \N__38792\ : std_logic;
signal \N__38791\ : std_logic;
signal \N__38788\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38721\ : std_logic;
signal \N__38718\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38667\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38661\ : std_logic;
signal \N__38658\ : std_logic;
signal \N__38655\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38562\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38544\ : std_logic;
signal \N__38541\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38526\ : std_logic;
signal \N__38523\ : std_logic;
signal \N__38520\ : std_logic;
signal \N__38517\ : std_logic;
signal \N__38514\ : std_logic;
signal \N__38511\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38484\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38478\ : std_logic;
signal \N__38475\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38439\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38424\ : std_logic;
signal \N__38421\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38400\ : std_logic;
signal \N__38397\ : std_logic;
signal \N__38394\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38382\ : std_logic;
signal \N__38379\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38349\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38345\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38330\ : std_logic;
signal \N__38327\ : std_logic;
signal \N__38324\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38307\ : std_logic;
signal \N__38304\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38286\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38244\ : std_logic;
signal \N__38241\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38235\ : std_logic;
signal \N__38232\ : std_logic;
signal \N__38229\ : std_logic;
signal \N__38226\ : std_logic;
signal \N__38223\ : std_logic;
signal \N__38220\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38211\ : std_logic;
signal \N__38210\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38197\ : std_logic;
signal \N__38194\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38159\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38153\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38142\ : std_logic;
signal \N__38139\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38111\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38102\ : std_logic;
signal \N__38099\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38087\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38052\ : std_logic;
signal \N__38049\ : std_logic;
signal \N__38046\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38040\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38027\ : std_logic;
signal \N__38024\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38016\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37971\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37952\ : std_logic;
signal \N__37949\ : std_logic;
signal \N__37946\ : std_logic;
signal \N__37943\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37925\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37914\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37908\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37906\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37897\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37872\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37863\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37857\ : std_logic;
signal \N__37854\ : std_logic;
signal \N__37851\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37806\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37755\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37747\ : std_logic;
signal \N__37744\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37711\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37677\ : std_logic;
signal \N__37674\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37659\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37639\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37621\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37591\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37566\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37546\ : std_logic;
signal \N__37543\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37465\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37429\ : std_logic;
signal \N__37426\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37407\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37399\ : std_logic;
signal \N__37396\ : std_logic;
signal \N__37393\ : std_logic;
signal \N__37390\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37377\ : std_logic;
signal \N__37374\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37333\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37311\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37248\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37201\ : std_logic;
signal \N__37198\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37185\ : std_logic;
signal \N__37182\ : std_logic;
signal \N__37179\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37173\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37123\ : std_logic;
signal \N__37120\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37104\ : std_logic;
signal \N__37101\ : std_logic;
signal \N__37098\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37084\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37074\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37029\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37023\ : std_logic;
signal \N__37020\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37012\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36976\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36923\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36879\ : std_logic;
signal \N__36876\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36793\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36771\ : std_logic;
signal \N__36768\ : std_logic;
signal \N__36765\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36654\ : std_logic;
signal \N__36651\ : std_logic;
signal \N__36648\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36642\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36624\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36614\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36592\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36583\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36528\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36498\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36468\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36457\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36445\ : std_logic;
signal \N__36442\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36427\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36424\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36411\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36408\ : std_logic;
signal \N__36405\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36360\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36354\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36289\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36279\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36240\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36189\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36094\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36048\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35968\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35945\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35918\ : std_logic;
signal \N__35913\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35870\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35727\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35703\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35687\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35670\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35518\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35475\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35373\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35343\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35282\ : std_logic;
signal \N__35281\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35266\ : std_logic;
signal \N__35263\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35244\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35068\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35040\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34912\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34714\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34653\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34510\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34321\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34306\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34272\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34151\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34142\ : std_logic;
signal \N__34139\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33862\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33839\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33256\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33009\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32722\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32012\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31266\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30976\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30903\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30851\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30385\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30252\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29336\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29076\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28922\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28438\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27366\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26747\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26262\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26034\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_1_19_0_\ : std_logic;
signal n12696 : std_logic;
signal n12697 : std_logic;
signal n12698 : std_logic;
signal n12699 : std_logic;
signal n12700 : std_logic;
signal n12701 : std_logic;
signal n12702 : std_logic;
signal n12703 : std_logic;
signal \bfn_1_20_0_\ : std_logic;
signal n12704 : std_logic;
signal n12705 : std_logic;
signal n12706 : std_logic;
signal n12707 : std_logic;
signal n12708 : std_logic;
signal n12709 : std_logic;
signal n12710 : std_logic;
signal n12711 : std_logic;
signal \bfn_1_21_0_\ : std_logic;
signal n12712 : std_logic;
signal n12713 : std_logic;
signal n12714 : std_logic;
signal n12715 : std_logic;
signal n12716 : std_logic;
signal \bfn_1_22_0_\ : std_logic;
signal n12811 : std_logic;
signal n12812 : std_logic;
signal n12813 : std_logic;
signal n12814 : std_logic;
signal n12815 : std_logic;
signal n12816 : std_logic;
signal n12817 : std_logic;
signal n12818 : std_logic;
signal \bfn_1_23_0_\ : std_logic;
signal n12819 : std_logic;
signal n12820 : std_logic;
signal n12821 : std_logic;
signal n12822 : std_logic;
signal n12823 : std_logic;
signal n12824 : std_logic;
signal n12825 : std_logic;
signal n12826 : std_logic;
signal \bfn_1_24_0_\ : std_logic;
signal n12827 : std_logic;
signal n12828 : std_logic;
signal n12829 : std_logic;
signal n12830 : std_logic;
signal n12831 : std_logic;
signal n12832 : std_logic;
signal n12833 : std_logic;
signal n12834 : std_logic;
signal \bfn_1_25_0_\ : std_logic;
signal n12835 : std_logic;
signal n12836 : std_logic;
signal n2882 : std_logic;
signal n2900 : std_logic;
signal n2876 : std_logic;
signal \n2908_cascade_\ : std_logic;
signal n2895 : std_logic;
signal \n2927_cascade_\ : std_logic;
signal \n3024_cascade_\ : std_logic;
signal \n14730_cascade_\ : std_logic;
signal \n3021_cascade_\ : std_logic;
signal n14728 : std_logic;
signal \n14150_cascade_\ : std_logic;
signal \n3128_cascade_\ : std_logic;
signal n14148 : std_logic;
signal \n3120_cascade_\ : std_logic;
signal \n3122_cascade_\ : std_logic;
signal n14146 : std_logic;
signal \debounce.reg_A_2\ : std_logic;
signal \debounce.reg_A_1\ : std_logic;
signal \debounce.reg_A_0\ : std_logic;
signal \reg_B_0\ : std_logic;
signal \debounce.n6_cascade_\ : std_logic;
signal \debounce.n16_cascade_\ : std_logic;
signal \debounce.n17\ : std_logic;
signal \reg_B_2\ : std_logic;
signal \n14129_cascade_\ : std_logic;
signal \debounce.cnt_reg_0\ : std_logic;
signal \bfn_1_31_0_\ : std_logic;
signal \debounce.cnt_reg_1\ : std_logic;
signal \debounce.n13013\ : std_logic;
signal \debounce.cnt_reg_2\ : std_logic;
signal \debounce.n13014\ : std_logic;
signal \debounce.cnt_reg_3\ : std_logic;
signal \debounce.n13015\ : std_logic;
signal \debounce.cnt_reg_4\ : std_logic;
signal \debounce.n13016\ : std_logic;
signal \debounce.cnt_reg_5\ : std_logic;
signal \debounce.n13017\ : std_logic;
signal \debounce.cnt_reg_6\ : std_logic;
signal \debounce.n13018\ : std_logic;
signal \debounce.cnt_reg_7\ : std_logic;
signal \debounce.n13019\ : std_logic;
signal \debounce.n13020\ : std_logic;
signal \debounce.cnt_reg_8\ : std_logic;
signal \bfn_1_32_0_\ : std_logic;
signal \debounce.n13021\ : std_logic;
signal \debounce.cnt_reg_9\ : std_logic;
signal \debounce.cnt_next_9__N_424\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal n12762 : std_logic;
signal n12763 : std_logic;
signal n12764 : std_logic;
signal n12765 : std_logic;
signal n12766 : std_logic;
signal n12767 : std_logic;
signal n12768 : std_logic;
signal n12769 : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal n12770 : std_logic;
signal n12771 : std_logic;
signal n12772 : std_logic;
signal n12773 : std_logic;
signal n12774 : std_logic;
signal n12775 : std_logic;
signal n12776 : std_logic;
signal n12777 : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal n12778 : std_logic;
signal n12779 : std_logic;
signal n2682 : std_logic;
signal n12780 : std_logic;
signal n12781 : std_logic;
signal n12782 : std_logic;
signal n12783 : std_logic;
signal n12784 : std_logic;
signal n12785 : std_logic;
signal \bfn_2_16_0_\ : std_logic;
signal n2801 : std_logic;
signal \bfn_2_17_0_\ : std_logic;
signal n12786 : std_logic;
signal n12787 : std_logic;
signal n12788 : std_logic;
signal n12789 : std_logic;
signal n12790 : std_logic;
signal n12791 : std_logic;
signal n12792 : std_logic;
signal n12793 : std_logic;
signal \bfn_2_18_0_\ : std_logic;
signal n12794 : std_logic;
signal n12795 : std_logic;
signal n12796 : std_logic;
signal n12797 : std_logic;
signal n12798 : std_logic;
signal n12799 : std_logic;
signal n12800 : std_logic;
signal n12801 : std_logic;
signal \bfn_2_19_0_\ : std_logic;
signal n12802 : std_logic;
signal n2783 : std_logic;
signal n12803 : std_logic;
signal n12804 : std_logic;
signal n12805 : std_logic;
signal n12806 : std_logic;
signal n12807 : std_logic;
signal n12808 : std_logic;
signal n12809 : std_logic;
signal \bfn_2_20_0_\ : std_logic;
signal n12810 : std_logic;
signal n2683 : std_logic;
signal n2677 : std_logic;
signal n2678 : std_logic;
signal n2797 : std_logic;
signal n2694 : std_logic;
signal n2793 : std_logic;
signal \n2726_cascade_\ : std_logic;
signal \n2621_cascade_\ : std_logic;
signal n2688 : std_logic;
signal n2696 : std_logic;
signal n2795 : std_logic;
signal \n2728_cascade_\ : std_logic;
signal n2691 : std_logic;
signal n2723 : std_logic;
signal n2790 : std_logic;
signal \n2723_cascade_\ : std_logic;
signal n2693 : std_logic;
signal n2697 : std_logic;
signal n2681 : std_logic;
signal n2794 : std_logic;
signal \n2826_cascade_\ : std_logic;
signal \n14362_cascade_\ : std_logic;
signal n2789 : std_logic;
signal n14346 : std_logic;
signal \n14350_cascade_\ : std_logic;
signal n14356 : std_logic;
signal n2782 : std_logic;
signal n2715 : std_logic;
signal n2785 : std_logic;
signal n2684 : std_logic;
signal n2716 : std_logic;
signal n2679 : std_logic;
signal n2709 : std_logic;
signal \n2711_cascade_\ : std_logic;
signal n14368 : std_logic;
signal n2796 : std_logic;
signal \n2742_cascade_\ : std_logic;
signal n2828 : std_logic;
signal n2788 : std_logic;
signal n2687 : std_logic;
signal n2792 : std_logic;
signal n2725 : std_logic;
signal n2791 : std_logic;
signal \bfn_2_25_0_\ : std_logic;
signal n12837 : std_logic;
signal n12838 : std_logic;
signal n12839 : std_logic;
signal n12840 : std_logic;
signal n12841 : std_logic;
signal n12842 : std_logic;
signal n2994 : std_logic;
signal n12843 : std_logic;
signal n12844 : std_logic;
signal n2993 : std_logic;
signal \bfn_2_26_0_\ : std_logic;
signal n2992 : std_logic;
signal n12845 : std_logic;
signal n12846 : std_logic;
signal n2990 : std_logic;
signal n12847 : std_logic;
signal n2989 : std_logic;
signal n12848 : std_logic;
signal n12849 : std_logic;
signal n12850 : std_logic;
signal n12851 : std_logic;
signal n12852 : std_logic;
signal n2985 : std_logic;
signal \bfn_2_27_0_\ : std_logic;
signal n12853 : std_logic;
signal n12854 : std_logic;
signal n12855 : std_logic;
signal n12856 : std_logic;
signal n12857 : std_logic;
signal n12858 : std_logic;
signal n12859 : std_logic;
signal n12860 : std_logic;
signal n2977 : std_logic;
signal \bfn_2_28_0_\ : std_logic;
signal n12861 : std_logic;
signal n2975 : std_logic;
signal n12862 : std_logic;
signal n12863 : std_logic;
signal \bfn_2_29_0_\ : std_logic;
signal n12892 : std_logic;
signal n12893 : std_logic;
signal n12894 : std_logic;
signal n12895 : std_logic;
signal n12896 : std_logic;
signal n12897 : std_logic;
signal n12898 : std_logic;
signal n12899 : std_logic;
signal \bfn_2_30_0_\ : std_logic;
signal n12900 : std_logic;
signal n12901 : std_logic;
signal n12902 : std_logic;
signal n12903 : std_logic;
signal n12904 : std_logic;
signal n3120 : std_logic;
signal n3187 : std_logic;
signal n12905 : std_logic;
signal n12906 : std_logic;
signal n12907 : std_logic;
signal \bfn_2_31_0_\ : std_logic;
signal n12908 : std_logic;
signal n12909 : std_logic;
signal n12910 : std_logic;
signal n12911 : std_logic;
signal n12912 : std_logic;
signal n12913 : std_logic;
signal n12914 : std_logic;
signal n12915 : std_logic;
signal \bfn_2_32_0_\ : std_logic;
signal n12916 : std_logic;
signal n12917 : std_logic;
signal n12918 : std_logic;
signal n12919 : std_logic;
signal n12920 : std_logic;
signal \bfn_3_14_0_\ : std_logic;
signal n12676 : std_logic;
signal n12677 : std_logic;
signal n12678 : std_logic;
signal n12679 : std_logic;
signal n12680 : std_logic;
signal n12681 : std_logic;
signal n12682 : std_logic;
signal n12683 : std_logic;
signal \bfn_3_15_0_\ : std_logic;
signal n12684 : std_logic;
signal n12685 : std_logic;
signal n12686 : std_logic;
signal n12687 : std_logic;
signal n12688 : std_logic;
signal n12689 : std_logic;
signal n12690 : std_logic;
signal n12691 : std_logic;
signal \bfn_3_16_0_\ : std_logic;
signal n12692 : std_logic;
signal n12693 : std_logic;
signal n12694 : std_logic;
signal n12695 : std_logic;
signal n2233 : std_logic;
signal n2300 : std_logic;
signal \n2233_cascade_\ : std_logic;
signal n2299 : std_logic;
signal \n2331_cascade_\ : std_logic;
signal n2301 : std_logic;
signal n2222 : std_logic;
signal \n2222_cascade_\ : std_logic;
signal n2289 : std_logic;
signal n2291 : std_logic;
signal \n2323_cascade_\ : std_logic;
signal \n2219_cascade_\ : std_logic;
signal n2286 : std_logic;
signal n2290 : std_logic;
signal n2293 : std_logic;
signal n2298 : std_logic;
signal n2295 : std_logic;
signal n2296 : std_logic;
signal n11977 : std_logic;
signal \n14808_cascade_\ : std_logic;
signal n14594 : std_logic;
signal n2219 : std_logic;
signal \n14598_cascade_\ : std_logic;
signal \n14604_cascade_\ : std_logic;
signal \n2247_cascade_\ : std_logic;
signal n2297 : std_logic;
signal n2288 : std_logic;
signal n2391 : std_logic;
signal n2287 : std_logic;
signal n2386 : std_logic;
signal \n2319_cascade_\ : std_logic;
signal n11971 : std_logic;
signal n2292 : std_logic;
signal n2324 : std_logic;
signal \n2324_cascade_\ : std_logic;
signal n2319 : std_logic;
signal \n14384_cascade_\ : std_logic;
signal n14382 : std_logic;
signal n14390 : std_logic;
signal n2689 : std_logic;
signal \n2622_cascade_\ : std_logic;
signal n2721 : std_logic;
signal n2728 : std_logic;
signal n2726 : std_logic;
signal \n2721_cascade_\ : std_logic;
signal n14348 : std_logic;
signal n2383 : std_logic;
signal n2622 : std_logic;
signal \n2628_cascade_\ : std_logic;
signal n2692 : std_logic;
signal n2724 : std_logic;
signal n2695 : std_logic;
signal n2628 : std_logic;
signal n2727 : std_logic;
signal n2700 : std_logic;
signal \n2732_cascade_\ : std_logic;
signal n2729 : std_logic;
signal \n11957_cascade_\ : std_logic;
signal n13808 : std_logic;
signal n2621 : std_logic;
signal n14668 : std_logic;
signal n2698 : std_logic;
signal n2730 : std_logic;
signal n2699 : std_logic;
signal n2701 : std_logic;
signal \n14650_cascade_\ : std_logic;
signal \n14654_cascade_\ : std_logic;
signal \n14660_cascade_\ : std_logic;
signal n14674 : std_logic;
signal \n2643_cascade_\ : std_logic;
signal n2686 : std_logic;
signal n2718 : std_logic;
signal n2690 : std_logic;
signal n2623 : std_logic;
signal n2722 : std_logic;
signal n2732 : std_logic;
signal n2799 : std_logic;
signal n2711 : std_logic;
signal n2778 : std_logic;
signal n2786 : std_logic;
signal n2719 : std_logic;
signal n2685 : std_logic;
signal n2717 : std_logic;
signal n2784 : std_logic;
signal \n2717_cascade_\ : std_logic;
signal n2713 : std_logic;
signal n2780 : std_logic;
signal n2798 : std_logic;
signal n2731 : std_logic;
signal n2680 : std_logic;
signal n2887 : std_logic;
signal n2820 : std_logic;
signal \n14690_cascade_\ : std_logic;
signal n14688 : std_logic;
signal \n14696_cascade_\ : std_logic;
signal n2714 : std_logic;
signal n2781 : std_logic;
signal n2720 : std_logic;
signal n2787 : std_logic;
signal n2823 : std_logic;
signal n2890 : std_logic;
signal n2827 : std_logic;
signal n2894 : std_logic;
signal n2822 : std_logic;
signal n2889 : std_logic;
signal n2982 : std_logic;
signal n2986 : std_logic;
signal n2879 : std_logic;
signal n2710 : std_logic;
signal n2777 : std_logic;
signal n2996 : std_logic;
signal \n3028_cascade_\ : std_logic;
signal n2988 : std_logic;
signal n2880 : std_logic;
signal n2979 : std_logic;
signal \n2912_cascade_\ : std_logic;
signal n2983 : std_logic;
signal \bfn_3_28_0_\ : std_logic;
signal n12864 : std_logic;
signal n12865 : std_logic;
signal n12866 : std_logic;
signal n12867 : std_logic;
signal n3096 : std_logic;
signal n12868 : std_logic;
signal n3028 : std_logic;
signal n3095 : std_logic;
signal n12869 : std_logic;
signal n3094 : std_logic;
signal n12870 : std_logic;
signal n12871 : std_logic;
signal n3026 : std_logic;
signal n3093 : std_logic;
signal \bfn_3_29_0_\ : std_logic;
signal n3025 : std_logic;
signal n3092 : std_logic;
signal n12872 : std_logic;
signal n3024 : std_logic;
signal n3091 : std_logic;
signal n12873 : std_logic;
signal n3090 : std_logic;
signal n12874 : std_logic;
signal n3022 : std_logic;
signal n3089 : std_logic;
signal n12875 : std_logic;
signal n3021 : std_logic;
signal n3088 : std_logic;
signal n12876 : std_logic;
signal n3020 : std_logic;
signal n3087 : std_logic;
signal n12877 : std_logic;
signal n3086 : std_logic;
signal n12878 : std_logic;
signal n12879 : std_logic;
signal \bfn_3_30_0_\ : std_logic;
signal n3017 : std_logic;
signal n3084 : std_logic;
signal n12880 : std_logic;
signal n12881 : std_logic;
signal n12882 : std_logic;
signal n12883 : std_logic;
signal n12884 : std_logic;
signal n12885 : std_logic;
signal n12886 : std_logic;
signal n12887 : std_logic;
signal \bfn_3_31_0_\ : std_logic;
signal n12888 : std_logic;
signal n12889 : std_logic;
signal n12890 : std_logic;
signal n12891 : std_logic;
signal n3075 : std_logic;
signal n3082 : std_logic;
signal n3074 : std_logic;
signal n3173 : std_logic;
signal n3174 : std_logic;
signal n3079 : std_logic;
signal n3078 : std_logic;
signal n3076 : std_logic;
signal n3175 : std_logic;
signal \n3108_cascade_\ : std_logic;
signal n2232 : std_logic;
signal n2231 : std_logic;
signal n2221 : std_logic;
signal n2229 : std_logic;
signal \n2129_cascade_\ : std_logic;
signal n2228 : std_logic;
signal n2226 : std_logic;
signal n2225 : std_logic;
signal \n2228_cascade_\ : std_logic;
signal n14588 : std_logic;
signal n2201 : std_logic;
signal \bfn_4_17_0_\ : std_logic;
signal n2200 : std_logic;
signal n12657 : std_logic;
signal n2199 : std_logic;
signal n12658 : std_logic;
signal n12659 : std_logic;
signal n2197 : std_logic;
signal n12660 : std_logic;
signal n2129 : std_logic;
signal n2196 : std_logic;
signal n12661 : std_logic;
signal n12662 : std_logic;
signal n2194 : std_logic;
signal n12663 : std_logic;
signal n12664 : std_logic;
signal n2193 : std_logic;
signal \bfn_4_18_0_\ : std_logic;
signal n12665 : std_logic;
signal n12666 : std_logic;
signal n2190 : std_logic;
signal n12667 : std_logic;
signal n2189 : std_logic;
signal n12668 : std_logic;
signal n12669 : std_logic;
signal n2187 : std_logic;
signal n12670 : std_logic;
signal n12671 : std_logic;
signal n12672 : std_logic;
signal \bfn_4_19_0_\ : std_logic;
signal n12673 : std_logic;
signal n12674 : std_logic;
signal n12675 : std_logic;
signal n2214 : std_logic;
signal n2294 : std_logic;
signal n2186 : std_logic;
signal n2218 : std_logic;
signal n2285 : std_logic;
signal \n2218_cascade_\ : std_logic;
signal n2188 : std_logic;
signal n2220 : std_logic;
signal n14392 : std_logic;
signal n2313 : std_logic;
signal \n14398_cascade_\ : std_logic;
signal n2327 : std_logic;
signal \n2346_cascade_\ : std_logic;
signal n2394 : std_logic;
signal n2284 : std_logic;
signal n2316 : std_logic;
signal n2282 : std_logic;
signal n2314 : std_logic;
signal \n2314_cascade_\ : std_logic;
signal n2381 : std_logic;
signal n2392 : std_logic;
signal n2325 : std_logic;
signal n2320 : std_logic;
signal n2387 : std_logic;
signal n2382 : std_logic;
signal n2396 : std_logic;
signal n2329 : std_logic;
signal n2328 : std_logic;
signal n2395 : std_logic;
signal \n2427_cascade_\ : std_logic;
signal \n14620_cascade_\ : std_logic;
signal \n2526_cascade_\ : std_logic;
signal n14816 : std_logic;
signal \n2524_cascade_\ : std_logic;
signal \n14574_cascade_\ : std_logic;
signal \n2523_cascade_\ : std_logic;
signal n14576 : std_logic;
signal \n2527_cascade_\ : std_logic;
signal n2626 : std_logic;
signal n2617 : std_logic;
signal n2625 : std_logic;
signal \n2617_cascade_\ : std_logic;
signal n14812 : std_logic;
signal n2633 : std_logic;
signal \n2633_cascade_\ : std_logic;
signal n12059 : std_logic;
signal n2618 : std_logic;
signal n2614 : std_logic;
signal n2613 : std_logic;
signal n2619 : std_logic;
signal n2897 : std_logic;
signal n2712 : std_logic;
signal n2779 : std_logic;
signal n2878 : std_logic;
signal \n2811_cascade_\ : std_logic;
signal n2733 : std_logic;
signal n2800 : std_logic;
signal \n2832_cascade_\ : std_logic;
signal n2833 : std_logic;
signal n2830 : std_logic;
signal \n11953_cascade_\ : std_logic;
signal n13857 : std_logic;
signal n2815 : std_logic;
signal n14702 : std_logic;
signal n2812 : std_logic;
signal n2813 : std_logic;
signal \n14708_cascade_\ : std_logic;
signal n2811 : std_logic;
signal n2809 : std_logic;
signal \n14714_cascade_\ : std_logic;
signal n2808 : std_logic;
signal n2816 : std_logic;
signal \n2841_cascade_\ : std_logic;
signal n2883 : std_logic;
signal n2885 : std_logic;
signal n2818 : std_logic;
signal n3081 : std_logic;
signal n2810 : std_logic;
signal n2877 : std_logic;
signal n2976 : std_logic;
signal n2886 : std_logic;
signal n2819 : std_logic;
signal n2918 : std_logic;
signal n2927 : std_logic;
signal n2926 : std_logic;
signal \n2918_cascade_\ : std_logic;
signal n2825 : std_logic;
signal n2892 : std_logic;
signal n2921 : std_logic;
signal n2922 : std_logic;
signal \n2924_cascade_\ : std_logic;
signal n2919 : std_logic;
signal \n14212_cascade_\ : std_logic;
signal n14216 : std_logic;
signal n2817 : std_logic;
signal n2884 : std_logic;
signal n2916 : std_logic;
signal n2981 : std_logic;
signal n2929 : std_logic;
signal n14222 : std_logic;
signal n2915 : std_logic;
signal \n14224_cascade_\ : std_logic;
signal n2914 : std_logic;
signal n2910 : std_logic;
signal \n14230_cascade_\ : std_logic;
signal n2912 : std_logic;
signal n2908 : std_logic;
signal n2907 : std_logic;
signal \n14236_cascade_\ : std_logic;
signal n2909 : std_logic;
signal \n2940_cascade_\ : std_logic;
signal n2997 : std_logic;
signal n2911 : std_logic;
signal n2978 : std_logic;
signal n2995 : std_logic;
signal n3000 : std_logic;
signal n3015 : std_logic;
signal n14736 : std_logic;
signal n3014 : std_logic;
signal \n14742_cascade_\ : std_logic;
signal n3011 : std_logic;
signal n3009 : std_logic;
signal \n14748_cascade_\ : std_logic;
signal n3006 : std_logic;
signal n3008 : std_logic;
signal \n14754_cascade_\ : std_logic;
signal n3007 : std_logic;
signal n3099 : std_logic;
signal \n3039_cascade_\ : std_logic;
signal n3018 : std_logic;
signal n3085 : std_logic;
signal n3098 : std_logic;
signal \n3130_cascade_\ : std_logic;
signal n3101 : std_logic;
signal n3097 : std_logic;
signal n3100 : std_logic;
signal \n3132_cascade_\ : std_logic;
signal n11945 : std_logic;
signal n3080 : std_logic;
signal n3013 : std_logic;
signal \n23_adj_715_cascade_\ : std_logic;
signal n3123 : std_logic;
signal n3190 : std_logic;
signal n3121 : std_logic;
signal n3188 : std_logic;
signal n3192 : std_logic;
signal n3125 : std_logic;
signal n3127 : std_logic;
signal n3194 : std_logic;
signal \n3226_cascade_\ : std_logic;
signal n3119 : std_logic;
signal n3186 : std_logic;
signal \n3218_cascade_\ : std_logic;
signal n3180 : std_logic;
signal \n3212_cascade_\ : std_logic;
signal n14798 : std_logic;
signal n3107 : std_logic;
signal n3106 : std_logic;
signal n3105 : std_logic;
signal n3195 : std_logic;
signal \n3138_cascade_\ : std_logic;
signal n3128 : std_logic;
signal n3181 : std_logic;
signal n3184 : std_logic;
signal n3117 : std_logic;
signal n3083 : std_logic;
signal n13831 : std_logic;
signal n3114 : std_logic;
signal \n3115_cascade_\ : std_logic;
signal n14156 : std_logic;
signal n3113 : std_logic;
signal \n14162_cascade_\ : std_logic;
signal \n14168_cascade_\ : std_logic;
signal n3108 : std_logic;
signal n14174 : std_logic;
signal n3010 : std_logic;
signal n3077 : std_logic;
signal n14264 : std_logic;
signal n14260 : std_logic;
signal n2130 : std_logic;
signal \n14324_cascade_\ : std_logic;
signal n13787 : std_logic;
signal n2127 : std_logic;
signal \n2127_cascade_\ : std_logic;
signal n14318 : std_logic;
signal n2131 : std_logic;
signal n2198 : std_logic;
signal \n2131_cascade_\ : std_logic;
signal n2230 : std_logic;
signal n14584 : std_logic;
signal n2191 : std_logic;
signal n2223 : std_logic;
signal n2192 : std_logic;
signal n2224 : std_logic;
signal n14330 : std_logic;
signal \n2116_cascade_\ : std_logic;
signal \n2148_cascade_\ : std_logic;
signal n2195 : std_logic;
signal n2227 : std_logic;
signal n2128 : std_logic;
signal n2126 : std_logic;
signal \n2128_cascade_\ : std_logic;
signal n14316 : std_logic;
signal n2125 : std_logic;
signal n2185 : std_logic;
signal n2217 : std_logic;
signal n2183 : std_logic;
signal n2116 : std_logic;
signal n2215 : std_logic;
signal n2184 : std_logic;
signal n2122 : std_logic;
signal n2124 : std_logic;
signal n2401 : std_logic;
signal n2390 : std_logic;
signal n2323 : std_logic;
signal n2118 : std_logic;
signal n2393 : std_logic;
signal n2326 : std_logic;
signal n2330 : std_logic;
signal n2397 : std_logic;
signal n2322 : std_logic;
signal n2389 : std_logic;
signal n2399 : std_logic;
signal n2332 : std_logic;
signal n2388 : std_logic;
signal n2321 : std_logic;
signal \n2420_cascade_\ : std_logic;
signal n14622 : std_logic;
signal n2398 : std_logic;
signal n2331 : std_logic;
signal \n2430_cascade_\ : std_logic;
signal n2400 : std_logic;
signal n2333 : std_logic;
signal \n2432_cascade_\ : std_logic;
signal n11967 : std_logic;
signal \n2528_cascade_\ : std_logic;
signal n2627 : std_logic;
signal n2384 : std_logic;
signal n2317 : std_logic;
signal n13828 : std_logic;
signal n14628 : std_logic;
signal n2318 : std_logic;
signal n2385 : std_logic;
signal \n2417_cascade_\ : std_logic;
signal n14634 : std_logic;
signal \n14640_cascade_\ : std_logic;
signal \n2445_cascade_\ : std_logic;
signal \n2530_cascade_\ : std_logic;
signal n14646 : std_logic;
signal \n2533_cascade_\ : std_logic;
signal n12063 : std_logic;
signal n2632 : std_logic;
signal n14188 : std_logic;
signal \n2515_cascade_\ : std_logic;
signal n14117 : std_logic;
signal \n14194_cascade_\ : std_logic;
signal \n2544_cascade_\ : std_logic;
signal n2631 : std_logic;
signal \n2513_cascade_\ : std_logic;
signal n2612 : std_logic;
signal n2629 : std_logic;
signal n2899 : std_logic;
signal n2832 : std_logic;
signal n2630 : std_logic;
signal n2620 : std_logic;
signal n2901 : std_logic;
signal n2824 : std_logic;
signal n2891 : std_logic;
signal n2923 : std_logic;
signal \n2923_cascade_\ : std_logic;
signal n14214 : std_logic;
signal n2896 : std_logic;
signal n2829 : std_logic;
signal n2928 : std_logic;
signal n2821 : std_logic;
signal n2888 : std_logic;
signal n2881 : std_logic;
signal n2814 : std_logic;
signal n2893 : std_logic;
signal n2826 : std_logic;
signal n2925 : std_logic;
signal n2615 : std_logic;
signal n2831 : std_logic;
signal n2898 : std_logic;
signal n2930 : std_logic;
signal n2991 : std_logic;
signal n2924 : std_logic;
signal n2913 : std_logic;
signal n2980 : std_logic;
signal n3012 : std_logic;
signal n2933 : std_logic;
signal n12053 : std_logic;
signal n2987 : std_logic;
signal n2920 : std_logic;
signal n2999 : std_logic;
signal n2932 : std_logic;
signal n3001 : std_logic;
signal n3033 : std_logic;
signal \n3033_cascade_\ : std_logic;
signal n3032 : std_logic;
signal n3182 : std_logic;
signal n3115 : std_logic;
signal n2998 : std_logic;
signal n2931 : std_logic;
signal n3030 : std_logic;
signal n3029 : std_logic;
signal n3031 : std_logic;
signal \n3030_cascade_\ : std_logic;
signal n11947 : std_logic;
signal n3019 : std_logic;
signal n3027 : std_logic;
signal \n13871_cascade_\ : std_logic;
signal n3023 : std_logic;
signal n14078 : std_logic;
signal n3199 : std_logic;
signal n3132 : std_logic;
signal n3129 : std_logic;
signal n3196 : std_logic;
signal \n3228_cascade_\ : std_logic;
signal n14768 : std_logic;
signal n3200 : std_logic;
signal n3133 : std_logic;
signal n3198 : std_logic;
signal n3131 : std_logic;
signal n2917 : std_logic;
signal n2984 : std_logic;
signal n3016 : std_logic;
signal n3124 : std_logic;
signal n3191 : std_logic;
signal n14804 : std_logic;
signal n14025 : std_logic;
signal \n3237_cascade_\ : std_logic;
signal n13_adj_713 : std_logic;
signal n3179 : std_logic;
signal n3112 : std_logic;
signal n14770 : std_logic;
signal \n14776_cascade_\ : std_logic;
signal n3122 : std_logic;
signal n3189 : std_logic;
signal n3116 : std_logic;
signal n3183 : std_logic;
signal n3185 : std_logic;
signal n3118 : std_logic;
signal \n27_adj_716_cascade_\ : std_logic;
signal n14266 : std_logic;
signal n35_adj_719 : std_logic;
signal \n17_adj_714_cascade_\ : std_logic;
signal n3109 : std_logic;
signal n3176 : std_logic;
signal \n33_adj_718_cascade_\ : std_logic;
signal n14272 : std_logic;
signal n14268 : std_logic;
signal \n14262_cascade_\ : std_logic;
signal n14282 : std_logic;
signal n3111 : std_logic;
signal n3178 : std_logic;
signal n3110 : std_logic;
signal n3177 : std_logic;
signal n2283 : std_logic;
signal n2216 : std_logic;
signal n2315 : std_logic;
signal \bfn_6_17_0_\ : std_logic;
signal n12639 : std_logic;
signal n2099 : std_logic;
signal n12640 : std_logic;
signal n2098 : std_logic;
signal n12641 : std_logic;
signal n2097 : std_logic;
signal n12642 : std_logic;
signal n2096 : std_logic;
signal n12643 : std_logic;
signal n2095 : std_logic;
signal n12644 : std_logic;
signal n2094 : std_logic;
signal n12645 : std_logic;
signal n12646 : std_logic;
signal n2093 : std_logic;
signal \bfn_6_18_0_\ : std_logic;
signal n2092 : std_logic;
signal n12647 : std_logic;
signal n12648 : std_logic;
signal n2090 : std_logic;
signal n12649 : std_logic;
signal n12650 : std_logic;
signal n12651 : std_logic;
signal n12652 : std_logic;
signal n2086 : std_logic;
signal n12653 : std_logic;
signal n12654 : std_logic;
signal \bfn_6_19_0_\ : std_logic;
signal n2084 : std_logic;
signal n12655 : std_logic;
signal n12656 : std_logic;
signal n2115 : std_logic;
signal n2091 : std_logic;
signal n2123 : std_logic;
signal \n14558_cascade_\ : std_logic;
signal n2101 : std_logic;
signal \n2049_cascade_\ : std_logic;
signal n2018 : std_logic;
signal n2085 : std_logic;
signal \n2018_cascade_\ : std_logic;
signal n2117 : std_logic;
signal n2089 : std_logic;
signal n2121 : std_logic;
signal n2501 : std_logic;
signal \bfn_6_21_0_\ : std_logic;
signal n12717 : std_logic;
signal n2432 : std_logic;
signal n2499 : std_logic;
signal n12718 : std_logic;
signal n2431 : std_logic;
signal n2498 : std_logic;
signal n12719 : std_logic;
signal n2430 : std_logic;
signal n2497 : std_logic;
signal n12720 : std_logic;
signal n2429 : std_logic;
signal n2496 : std_logic;
signal n12721 : std_logic;
signal n2428 : std_logic;
signal n2495 : std_logic;
signal n12722 : std_logic;
signal n2427 : std_logic;
signal n2494 : std_logic;
signal n12723 : std_logic;
signal n12724 : std_logic;
signal \bfn_6_22_0_\ : std_logic;
signal n2425 : std_logic;
signal n2492 : std_logic;
signal n12725 : std_logic;
signal n2424 : std_logic;
signal n2491 : std_logic;
signal n12726 : std_logic;
signal n12727 : std_logic;
signal n12728 : std_logic;
signal n2421 : std_logic;
signal n2488 : std_logic;
signal n12729 : std_logic;
signal n2420 : std_logic;
signal n2487 : std_logic;
signal n12730 : std_logic;
signal n12731 : std_logic;
signal n12732 : std_logic;
signal \bfn_6_23_0_\ : std_logic;
signal n2417 : std_logic;
signal n2484 : std_logic;
signal n12733 : std_logic;
signal n2416 : std_logic;
signal n2483 : std_logic;
signal n12734 : std_logic;
signal n2415 : std_logic;
signal n2482 : std_logic;
signal n12735 : std_logic;
signal n2414 : std_logic;
signal n2481 : std_logic;
signal n12736 : std_logic;
signal n2413 : std_logic;
signal n2480 : std_logic;
signal n12737 : std_logic;
signal n2412 : std_logic;
signal n12738 : std_logic;
signal n2433 : std_logic;
signal n2500 : std_logic;
signal n2601 : std_logic;
signal \bfn_6_24_0_\ : std_logic;
signal n2533 : std_logic;
signal n2600 : std_logic;
signal n12739 : std_logic;
signal n2532 : std_logic;
signal n2599 : std_logic;
signal n12740 : std_logic;
signal n2531 : std_logic;
signal n2598 : std_logic;
signal n12741 : std_logic;
signal n2530 : std_logic;
signal n2597 : std_logic;
signal n12742 : std_logic;
signal n2529 : std_logic;
signal n2596 : std_logic;
signal n12743 : std_logic;
signal n2528 : std_logic;
signal n2595 : std_logic;
signal n12744 : std_logic;
signal n2527 : std_logic;
signal n2594 : std_logic;
signal n12745 : std_logic;
signal n12746 : std_logic;
signal n2526 : std_logic;
signal n2593 : std_logic;
signal \bfn_6_25_0_\ : std_logic;
signal n12747 : std_logic;
signal n2524 : std_logic;
signal n2591 : std_logic;
signal n12748 : std_logic;
signal n2523 : std_logic;
signal n2590 : std_logic;
signal n12749 : std_logic;
signal n2589 : std_logic;
signal n12750 : std_logic;
signal n2588 : std_logic;
signal n12751 : std_logic;
signal n2520 : std_logic;
signal n2587 : std_logic;
signal n12752 : std_logic;
signal n2519 : std_logic;
signal n2586 : std_logic;
signal n12753 : std_logic;
signal n12754 : std_logic;
signal n2585 : std_logic;
signal \bfn_6_26_0_\ : std_logic;
signal n12755 : std_logic;
signal n2516 : std_logic;
signal n2583 : std_logic;
signal n12756 : std_logic;
signal n2515 : std_logic;
signal n2582 : std_logic;
signal n12757 : std_logic;
signal n2514 : std_logic;
signal n2581 : std_logic;
signal n12758 : std_logic;
signal n2513 : std_logic;
signal n2580 : std_logic;
signal n12759 : std_logic;
signal n12760 : std_logic;
signal n2511 : std_logic;
signal n12761 : std_logic;
signal n2610 : std_logic;
signal n2418 : std_logic;
signal n2485 : std_logic;
signal n2517 : std_logic;
signal n2584 : std_logic;
signal \n2517_cascade_\ : std_logic;
signal n2616 : std_logic;
signal n2512 : std_logic;
signal n2579 : std_logic;
signal n2611 : std_logic;
signal n3130 : std_logic;
signal n3197 : std_logic;
signal n3193 : std_logic;
signal n3126 : std_logic;
signal n3201 : std_logic;
signal \n3233_cascade_\ : std_logic;
signal \n11943_cascade_\ : std_logic;
signal n13875 : std_logic;
signal \n29_adj_717_cascade_\ : std_logic;
signal n14270 : std_logic;
signal \n11941_cascade_\ : std_logic;
signal n11878 : std_logic;
signal n14782 : std_logic;
signal n14788 : std_logic;
signal \n14300_cascade_\ : std_logic;
signal \n14302_cascade_\ : std_logic;
signal \n14304_cascade_\ : std_logic;
signal \n14306_cascade_\ : std_logic;
signal n14308 : std_logic;
signal n5_adj_704 : std_logic;
signal n12039 : std_logic;
signal \n14292_cascade_\ : std_logic;
signal n14284 : std_logic;
signal \n14286_cascade_\ : std_logic;
signal n14288 : std_logic;
signal n14294 : std_logic;
signal \n14296_cascade_\ : std_logic;
signal n14298 : std_logic;
signal n45_adj_720 : std_logic;
signal \ENCODER0_A_N\ : std_logic;
signal \n1922_cascade_\ : std_logic;
signal n2021 : std_logic;
signal n2088 : std_logic;
signal \n2021_cascade_\ : std_logic;
signal n2120 : std_logic;
signal n2020 : std_logic;
signal n2087 : std_logic;
signal \n2020_cascade_\ : std_logic;
signal n2119 : std_logic;
signal \n14446_cascade_\ : std_logic;
signal n11985 : std_logic;
signal \n14450_cascade_\ : std_logic;
signal \n1950_cascade_\ : std_logic;
signal n2017 : std_logic;
signal n2025 : std_logic;
signal n2028 : std_logic;
signal n2026 : std_logic;
signal \n2025_cascade_\ : std_logic;
signal n2027 : std_logic;
signal n2032 : std_logic;
signal n2031 : std_logic;
signal \n2032_cascade_\ : std_logic;
signal n2022 : std_logic;
signal n2024 : std_logic;
signal n2023 : std_logic;
signal n14544 : std_logic;
signal n11981 : std_logic;
signal n2029 : std_logic;
signal \n14550_cascade_\ : std_logic;
signal n2030 : std_logic;
signal n14552 : std_logic;
signal n2100 : std_logic;
signal n2033 : std_logic;
signal n2132 : std_logic;
signal \n2132_cascade_\ : std_logic;
signal n2133 : std_logic;
signal n11909 : std_logic;
signal n307 : std_logic;
signal n310 : std_logic;
signal n312 : std_logic;
signal n313 : std_logic;
signal n314 : std_logic;
signal n317 : std_logic;
signal n14184 : std_logic;
signal n2490 : std_logic;
signal n2423 : std_logic;
signal n2522 : std_logic;
signal n2489 : std_logic;
signal n2422 : std_logic;
signal n2521 : std_logic;
signal n2426 : std_logic;
signal n2493 : std_logic;
signal n2525 : std_logic;
signal n2592 : std_logic;
signal \n2525_cascade_\ : std_logic;
signal n2624 : std_logic;
signal n2486 : std_logic;
signal n2419 : std_logic;
signal n2518 : std_logic;
signal n315 : std_logic;
signal n311 : std_logic;
signal \bfn_7_25_0_\ : std_logic;
signal n15485 : std_logic;
signal n3237 : std_logic;
signal n12952 : std_logic;
signal n15451 : std_logic;
signal n3138 : std_logic;
signal n12953 : std_logic;
signal n15418 : std_logic;
signal n3039 : std_logic;
signal n12954 : std_logic;
signal n15384 : std_logic;
signal n2940 : std_logic;
signal n12955 : std_logic;
signal n15352 : std_logic;
signal n2841 : std_logic;
signal n12956 : std_logic;
signal n15322 : std_logic;
signal n2742 : std_logic;
signal n12957 : std_logic;
signal n15292 : std_logic;
signal n2643 : std_logic;
signal encoder0_position_scaled_7 : std_logic;
signal n12958 : std_logic;
signal n12959 : std_logic;
signal n15830 : std_logic;
signal n2544 : std_logic;
signal \bfn_7_26_0_\ : std_logic;
signal n15802 : std_logic;
signal n2445 : std_logic;
signal n12960 : std_logic;
signal n15775 : std_logic;
signal n2346 : std_logic;
signal n12961 : std_logic;
signal n15748 : std_logic;
signal n2247 : std_logic;
signal n12962 : std_logic;
signal n15722 : std_logic;
signal n2148 : std_logic;
signal n12963 : std_logic;
signal n15697 : std_logic;
signal n2049 : std_logic;
signal n12964 : std_logic;
signal n12965 : std_logic;
signal n15652 : std_logic;
signal n12966 : std_logic;
signal n12967 : std_logic;
signal \bfn_7_27_0_\ : std_logic;
signal n12968 : std_logic;
signal n12969 : std_logic;
signal n12970 : std_logic;
signal n12971 : std_logic;
signal n12972 : std_logic;
signal n12973 : std_logic;
signal n12974 : std_logic;
signal n12051 : std_logic;
signal n15490 : std_logic;
signal n319 : std_logic;
signal \bfn_7_29_0_\ : std_logic;
signal n318 : std_logic;
signal n3301 : std_logic;
signal n12921 : std_logic;
signal n3233 : std_logic;
signal n3300 : std_logic;
signal n12922 : std_logic;
signal n3232 : std_logic;
signal n3299 : std_logic;
signal n12923 : std_logic;
signal n3231 : std_logic;
signal n12924 : std_logic;
signal n3298 : std_logic;
signal n3230 : std_logic;
signal n15079 : std_logic;
signal n12925 : std_logic;
signal n3229 : std_logic;
signal n3296 : std_logic;
signal n12926 : std_logic;
signal n3228 : std_logic;
signal n3295 : std_logic;
signal n12927 : std_logic;
signal n12928 : std_logic;
signal n3227 : std_logic;
signal n3294 : std_logic;
signal \bfn_7_30_0_\ : std_logic;
signal n3226 : std_logic;
signal n3293 : std_logic;
signal n12929 : std_logic;
signal n3225 : std_logic;
signal n3292 : std_logic;
signal n12930 : std_logic;
signal n3224 : std_logic;
signal n3291 : std_logic;
signal n12931 : std_logic;
signal n3223 : std_logic;
signal n3290 : std_logic;
signal n12932 : std_logic;
signal n3222 : std_logic;
signal n3289 : std_logic;
signal n12933 : std_logic;
signal n3221 : std_logic;
signal n3288 : std_logic;
signal n12934 : std_logic;
signal n3220 : std_logic;
signal n3287 : std_logic;
signal n12935 : std_logic;
signal n12936 : std_logic;
signal n3219 : std_logic;
signal n3286 : std_logic;
signal \bfn_7_31_0_\ : std_logic;
signal n3218 : std_logic;
signal n3285 : std_logic;
signal n12937 : std_logic;
signal n3217 : std_logic;
signal n3284 : std_logic;
signal n12938 : std_logic;
signal n3216 : std_logic;
signal n3283 : std_logic;
signal n12939 : std_logic;
signal n3215 : std_logic;
signal n3282 : std_logic;
signal n12940 : std_logic;
signal n3214 : std_logic;
signal n3281 : std_logic;
signal n12941 : std_logic;
signal n3213 : std_logic;
signal n3280 : std_logic;
signal n12942 : std_logic;
signal n3212 : std_logic;
signal n3279 : std_logic;
signal n12943 : std_logic;
signal n12944 : std_logic;
signal n3211 : std_logic;
signal n3278 : std_logic;
signal \bfn_7_32_0_\ : std_logic;
signal n3210 : std_logic;
signal n3277 : std_logic;
signal n12945 : std_logic;
signal n3209 : std_logic;
signal n3276 : std_logic;
signal n12946 : std_logic;
signal n3208 : std_logic;
signal n3275 : std_logic;
signal n12947 : std_logic;
signal n3207 : std_logic;
signal n3274 : std_logic;
signal n12948 : std_logic;
signal n3206 : std_logic;
signal n3273 : std_logic;
signal n12949 : std_logic;
signal n3205 : std_logic;
signal n3272 : std_logic;
signal n12950 : std_logic;
signal n3204 : std_logic;
signal n12951 : std_logic;
signal n3271 : std_logic;
signal n2001 : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal n2000 : std_logic;
signal n12622 : std_logic;
signal n1999 : std_logic;
signal n12623 : std_logic;
signal n1998 : std_logic;
signal n12624 : std_logic;
signal n1997 : std_logic;
signal n12625 : std_logic;
signal n1996 : std_logic;
signal n12626 : std_logic;
signal n1995 : std_logic;
signal n12627 : std_logic;
signal n1994 : std_logic;
signal n12628 : std_logic;
signal n12629 : std_logic;
signal n1993 : std_logic;
signal \bfn_9_17_0_\ : std_logic;
signal n1992 : std_logic;
signal n12630 : std_logic;
signal n1991 : std_logic;
signal n12631 : std_logic;
signal n1990 : std_logic;
signal n12632 : std_logic;
signal n1922 : std_logic;
signal n1989 : std_logic;
signal n12633 : std_logic;
signal n1988 : std_logic;
signal n12634 : std_logic;
signal n12635 : std_logic;
signal n1986 : std_logic;
signal n12636 : std_logic;
signal n12637 : std_logic;
signal n1985 : std_logic;
signal \bfn_9_18_0_\ : std_logic;
signal n15674 : std_logic;
signal n12638 : std_logic;
signal n2016 : std_logic;
signal n1921 : std_logic;
signal n14530 : std_logic;
signal n1918 : std_logic;
signal n1919 : std_logic;
signal n305 : std_logic;
signal n306 : std_logic;
signal n308 : std_logic;
signal n309 : std_logic;
signal n33_adj_651 : std_logic;
signal n33 : std_logic;
signal \bfn_9_22_0_\ : std_logic;
signal n32 : std_logic;
signal n12975 : std_logic;
signal n31_adj_649 : std_logic;
signal n31 : std_logic;
signal n12976 : std_logic;
signal n30_adj_648 : std_logic;
signal n12977 : std_logic;
signal n29_adj_647 : std_logic;
signal n29 : std_logic;
signal n12978 : std_logic;
signal n28_adj_646 : std_logic;
signal n28 : std_logic;
signal n12979 : std_logic;
signal n27_adj_645 : std_logic;
signal n27 : std_logic;
signal n12980 : std_logic;
signal n26_adj_644 : std_logic;
signal n26 : std_logic;
signal n12981 : std_logic;
signal n12982 : std_logic;
signal n25_adj_643 : std_logic;
signal n25 : std_logic;
signal \bfn_9_23_0_\ : std_logic;
signal n24_adj_642 : std_logic;
signal n24 : std_logic;
signal n12983 : std_logic;
signal n23_adj_641 : std_logic;
signal n23 : std_logic;
signal n12984 : std_logic;
signal n22 : std_logic;
signal n12985 : std_logic;
signal n21 : std_logic;
signal n12986 : std_logic;
signal n20 : std_logic;
signal n12987 : std_logic;
signal n19_adj_637 : std_logic;
signal n19 : std_logic;
signal n12988 : std_logic;
signal n18_adj_636 : std_logic;
signal n18 : std_logic;
signal n12989 : std_logic;
signal n12990 : std_logic;
signal \bfn_9_24_0_\ : std_logic;
signal n12991 : std_logic;
signal n12992 : std_logic;
signal n14_adj_632 : std_logic;
signal n14 : std_logic;
signal n12993 : std_logic;
signal n12994 : std_logic;
signal n12995 : std_logic;
signal n12996 : std_logic;
signal n12997 : std_logic;
signal n12998 : std_logic;
signal \bfn_9_25_0_\ : std_logic;
signal n12999 : std_logic;
signal n13000 : std_logic;
signal n13001 : std_logic;
signal n13002 : std_logic;
signal n4_adj_622 : std_logic;
signal n13003 : std_logic;
signal n13004 : std_logic;
signal n13005 : std_logic;
signal encoder0_position_scaled_8 : std_logic;
signal encoder0_position_scaled_14 : std_logic;
signal encoder0_position_scaled_10 : std_logic;
signal encoder0_position_scaled_12 : std_logic;
signal encoder0_position_scaled_13 : std_logic;
signal encoder0_position_scaled_15 : std_logic;
signal n15508 : std_logic;
signal encoder0_position_scaled_18 : std_logic;
signal encoder0_position_scaled_23 : std_logic;
signal encoder0_position_scaled_17 : std_logic;
signal \dti_N_333_cascade_\ : std_logic;
signal \reg_B_1\ : std_logic;
signal n14129 : std_logic;
signal n1377 : std_logic;
signal \bfn_9_29_0_\ : std_logic;
signal n13006 : std_logic;
signal n13007 : std_logic;
signal n13008 : std_logic;
signal n13009 : std_logic;
signal n15072 : std_logic;
signal n13010 : std_logic;
signal n13011 : std_logic;
signal n11526 : std_logic;
signal n13012 : std_logic;
signal n15075 : std_logic;
signal n15071 : std_logic;
signal dti_counter_5 : std_logic;
signal dti_counter_6 : std_logic;
signal \n14_adj_705_cascade_\ : std_logic;
signal dti_counter_2 : std_logic;
signal n10_adj_706 : std_logic;
signal dti_counter_0 : std_logic;
signal n15081 : std_logic;
signal dti_counter_3 : std_logic;
signal n15074 : std_logic;
signal dti_counter_4 : std_logic;
signal n15073 : std_logic;
signal dti_counter_7 : std_logic;
signal n15070 : std_logic;
signal dti_counter_1 : std_logic;
signal n15076 : std_logic;
signal commutation_state_prev_0 : std_logic;
signal n14929 : std_logic;
signal n14928 : std_logic;
signal \LED_c\ : std_logic;
signal \n1831_cascade_\ : std_logic;
signal n1930 : std_logic;
signal n1931 : std_logic;
signal n1933 : std_logic;
signal n1929 : std_logic;
signal \n14524_cascade_\ : std_logic;
signal \n14526_cascade_\ : std_logic;
signal \n1851_cascade_\ : std_logic;
signal n1928 : std_logic;
signal n1925 : std_logic;
signal \n1928_cascade_\ : std_logic;
signal n1923 : std_logic;
signal n14440 : std_logic;
signal n1932 : std_logic;
signal encoder0_position_0 : std_logic;
signal \bfn_10_18_0_\ : std_logic;
signal \quad_counter0.n13095\ : std_logic;
signal encoder0_position_2 : std_logic;
signal \quad_counter0.n13096\ : std_logic;
signal \quad_counter0.n13097\ : std_logic;
signal encoder0_position_4 : std_logic;
signal \quad_counter0.n13098\ : std_logic;
signal encoder0_position_5 : std_logic;
signal \quad_counter0.n13099\ : std_logic;
signal encoder0_position_6 : std_logic;
signal \quad_counter0.n13100\ : std_logic;
signal encoder0_position_7 : std_logic;
signal \quad_counter0.n13101\ : std_logic;
signal \quad_counter0.n13102\ : std_logic;
signal encoder0_position_8 : std_logic;
signal \bfn_10_19_0_\ : std_logic;
signal encoder0_position_9 : std_logic;
signal \quad_counter0.n13103\ : std_logic;
signal encoder0_position_10 : std_logic;
signal \quad_counter0.n13104\ : std_logic;
signal \quad_counter0.n13105\ : std_logic;
signal \quad_counter0.n13106\ : std_logic;
signal \quad_counter0.n13107\ : std_logic;
signal encoder0_position_14 : std_logic;
signal \quad_counter0.n13108\ : std_logic;
signal encoder0_position_15 : std_logic;
signal \quad_counter0.n13109\ : std_logic;
signal \quad_counter0.n13110\ : std_logic;
signal \bfn_10_20_0_\ : std_logic;
signal \quad_counter0.n13111\ : std_logic;
signal \quad_counter0.n13112\ : std_logic;
signal encoder0_position_19 : std_logic;
signal \quad_counter0.n13113\ : std_logic;
signal \quad_counter0.n13114\ : std_logic;
signal \quad_counter0.n13115\ : std_logic;
signal \quad_counter0.n13116\ : std_logic;
signal \quad_counter0.n13117\ : std_logic;
signal \quad_counter0.n13118\ : std_logic;
signal \bfn_10_21_0_\ : std_logic;
signal \quad_counter0.n13119\ : std_logic;
signal \quad_counter0.n13120\ : std_logic;
signal \quad_counter0.n13121\ : std_logic;
signal \quad_counter0.n13122\ : std_logic;
signal \quad_counter0.n13123\ : std_logic;
signal \quad_counter0.n13124\ : std_logic;
signal \quad_counter0.n13125\ : std_logic;
signal \bfn_10_22_0_\ : std_logic;
signal n12496 : std_logic;
signal n12497 : std_logic;
signal n12498 : std_logic;
signal n12499 : std_logic;
signal n12500 : std_logic;
signal n2563 : std_logic;
signal n13656 : std_logic;
signal n403 : std_logic;
signal n13_adj_631 : std_logic;
signal n38 : std_logic;
signal n402 : std_logic;
signal n39 : std_logic;
signal n2562 : std_logic;
signal n5187 : std_logic;
signal encoder0_position_11 : std_logic;
signal n22_adj_640 : std_logic;
signal encoder0_position_12 : std_logic;
signal n21_adj_639 : std_logic;
signal encoder0_position_13 : std_logic;
signal n20_adj_638 : std_logic;
signal n15_adj_633 : std_logic;
signal n6_adj_624 : std_logic;
signal \direction_N_537\ : std_logic;
signal \direction_N_537_cascade_\ : std_logic;
signal n1302 : std_logic;
signal n8_adj_626 : std_logic;
signal n5_adj_623 : std_logic;
signal n2_adj_620 : std_logic;
signal n9_adj_627 : std_logic;
signal encoder0_position_scaled_5 : std_logic;
signal encoder0_position_scaled_1 : std_logic;
signal \quad_counter0.direction_N_540\ : std_logic;
signal encoder0_position_scaled_9 : std_logic;
signal encoder0_position_scaled_20 : std_logic;
signal encoder0_position_scaled_11 : std_logic;
signal encoder0_position_scaled_21 : std_logic;
signal encoder0_position_scaled_19 : std_logic;
signal pwm_setpoint_4 : std_logic;
signal encoder0_position_scaled_22 : std_logic;
signal \quad_counter0.a_prev\ : std_logic;
signal \quad_counter0.direction_N_536\ : std_logic;
signal n26_adj_703 : std_logic;
signal \bfn_10_29_0_\ : std_logic;
signal n25_adj_702 : std_logic;
signal n13070 : std_logic;
signal n24_adj_701 : std_logic;
signal n13071 : std_logic;
signal n23_adj_700 : std_logic;
signal n13072 : std_logic;
signal n22_adj_699 : std_logic;
signal n13073 : std_logic;
signal n21_adj_698 : std_logic;
signal n13074 : std_logic;
signal n20_adj_697 : std_logic;
signal n13075 : std_logic;
signal n19_adj_696 : std_logic;
signal n13076 : std_logic;
signal n13077 : std_logic;
signal n18_adj_695 : std_logic;
signal \bfn_10_30_0_\ : std_logic;
signal n17_adj_694 : std_logic;
signal n13078 : std_logic;
signal n16_adj_693 : std_logic;
signal n13079 : std_logic;
signal n15_adj_692 : std_logic;
signal n13080 : std_logic;
signal n14_adj_691 : std_logic;
signal n13081 : std_logic;
signal n13_adj_690 : std_logic;
signal n13082 : std_logic;
signal n12_adj_689 : std_logic;
signal n13083 : std_logic;
signal n11_adj_688 : std_logic;
signal n13084 : std_logic;
signal n13085 : std_logic;
signal n10_adj_687 : std_logic;
signal \bfn_10_31_0_\ : std_logic;
signal n9_adj_686 : std_logic;
signal n13086 : std_logic;
signal n8_adj_685 : std_logic;
signal n13087 : std_logic;
signal n7_adj_684 : std_logic;
signal n13088 : std_logic;
signal n6_adj_683 : std_logic;
signal n13089 : std_logic;
signal blink_counter_21 : std_logic;
signal n13090 : std_logic;
signal blink_counter_22 : std_logic;
signal n13091 : std_logic;
signal blink_counter_23 : std_logic;
signal n13092 : std_logic;
signal n13093 : std_logic;
signal blink_counter_24 : std_logic;
signal \bfn_10_32_0_\ : std_logic;
signal n13094 : std_logic;
signal blink_counter_25 : std_logic;
signal \n1833_cascade_\ : std_logic;
signal n11989 : std_logic;
signal n304 : std_logic;
signal n1901 : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal n1833 : std_logic;
signal n1900 : std_logic;
signal n12606 : std_logic;
signal n1832 : std_logic;
signal n1899 : std_logic;
signal n12607 : std_logic;
signal n1831 : std_logic;
signal n1898 : std_logic;
signal n12608 : std_logic;
signal n1897 : std_logic;
signal n12609 : std_logic;
signal n1896 : std_logic;
signal n12610 : std_logic;
signal n12611 : std_logic;
signal n12612 : std_logic;
signal n12613 : std_logic;
signal n1893 : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal n12614 : std_logic;
signal n1891 : std_logic;
signal n12615 : std_logic;
signal n1890 : std_logic;
signal n12616 : std_logic;
signal n1889 : std_logic;
signal n12617 : std_logic;
signal n12618 : std_logic;
signal n1887 : std_logic;
signal n12619 : std_logic;
signal n1886 : std_logic;
signal n12620 : std_logic;
signal n12621 : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal n1892 : std_logic;
signal n1924 : std_logic;
signal \n1924_cascade_\ : std_logic;
signal n14438 : std_logic;
signal n1822 : std_logic;
signal \n1822_cascade_\ : std_logic;
signal n14534 : std_logic;
signal n1895 : std_logic;
signal n1927 : std_logic;
signal n1894 : std_logic;
signal n1926 : std_logic;
signal n1829 : std_logic;
signal n1885 : std_logic;
signal n1917 : std_logic;
signal n30 : std_logic;
signal encoder0_position_3 : std_logic;
signal n316 : std_logic;
signal n1888 : std_logic;
signal n1851 : std_logic;
signal n1920 : std_logic;
signal n1987 : std_logic;
signal \n1920_cascade_\ : std_logic;
signal n1950 : std_logic;
signal n2019 : std_logic;
signal n1819 : std_logic;
signal n16 : std_logic;
signal encoder0_position_29 : std_logic;
signal n404 : std_logic;
signal encoder0_position_17 : std_logic;
signal n16_adj_634 : std_logic;
signal n7_adj_625 : std_logic;
signal n3_adj_621 : std_logic;
signal n2566 : std_logic;
signal n7 : std_logic;
signal \n13662_cascade_\ : std_logic;
signal encoder0_position_26 : std_logic;
signal n2565 : std_logic;
signal encoder0_position_27 : std_logic;
signal \n13660_cascade_\ : std_logic;
signal \n832_cascade_\ : std_logic;
signal n2564 : std_logic;
signal \n13658_cascade_\ : std_logic;
signal encoder0_position_28 : std_logic;
signal encoder0_position_scaled_4 : std_logic;
signal \n929_cascade_\ : std_logic;
signal encoder0_position_30 : std_logic;
signal n13654 : std_logic;
signal \n829_cascade_\ : std_logic;
signal n12027 : std_logic;
signal \n861_cascade_\ : std_logic;
signal n6 : std_logic;
signal n4 : std_logic;
signal n40 : std_logic;
signal n5 : std_logic;
signal n5_adj_682 : std_logic;
signal n3 : std_logic;
signal \n5_adj_682_cascade_\ : std_logic;
signal n13653 : std_logic;
signal \bfn_11_24_0_\ : std_logic;
signal n12501 : std_logic;
signal n12502 : std_logic;
signal n831 : std_logic;
signal n898 : std_logic;
signal n12503 : std_logic;
signal n830 : std_logic;
signal n897 : std_logic;
signal n12504 : std_logic;
signal n12505 : std_logic;
signal n12506 : std_logic;
signal n2 : std_logic;
signal n14568 : std_logic;
signal n2561 : std_logic;
signal n828 : std_logic;
signal encoder0_position_scaled_3 : std_logic;
signal encoder0_position_scaled_6 : std_logic;
signal encoder0_position_scaled_2 : std_logic;
signal n25_adj_597 : std_logic;
signal \bfn_11_26_0_\ : std_logic;
signal n12426 : std_logic;
signal n12427 : std_logic;
signal n22_adj_594 : std_logic;
signal n12428 : std_logic;
signal n21_adj_593 : std_logic;
signal \pwm_setpoint_23_N_171_4\ : std_logic;
signal n12429 : std_logic;
signal n20_adj_592 : std_logic;
signal \pwm_setpoint_23_N_171_5\ : std_logic;
signal n12430 : std_logic;
signal n12431 : std_logic;
signal n18_adj_590 : std_logic;
signal \pwm_setpoint_23_N_171_7\ : std_logic;
signal n12432 : std_logic;
signal n12433 : std_logic;
signal n17_adj_589 : std_logic;
signal \pwm_setpoint_23_N_171_8\ : std_logic;
signal \bfn_11_27_0_\ : std_logic;
signal n16_adj_588 : std_logic;
signal n12434 : std_logic;
signal n15_adj_587 : std_logic;
signal n12435 : std_logic;
signal n14_adj_586 : std_logic;
signal \pwm_setpoint_23_N_171_11\ : std_logic;
signal n12436 : std_logic;
signal n12437 : std_logic;
signal n12_adj_584 : std_logic;
signal \pwm_setpoint_23_N_171_13\ : std_logic;
signal n12438 : std_logic;
signal n11_adj_583 : std_logic;
signal n12439 : std_logic;
signal n10_adj_582 : std_logic;
signal n12440 : std_logic;
signal n12441 : std_logic;
signal n9_adj_581 : std_logic;
signal \bfn_11_28_0_\ : std_logic;
signal n12442 : std_logic;
signal \pwm_setpoint_23_N_171_18\ : std_logic;
signal n12443 : std_logic;
signal n12444 : std_logic;
signal n12445 : std_logic;
signal n12446 : std_logic;
signal n12447 : std_logic;
signal n12448 : std_logic;
signal \n16_adj_664_cascade_\ : std_logic;
signal \n24_adj_669_cascade_\ : std_logic;
signal n8_adj_657 : std_logic;
signal n15144 : std_logic;
signal \pwm_setpoint_23_N_171_21\ : std_logic;
signal \pwm_setpoint_23_N_171_9\ : std_logic;
signal pwm_setpoint_9 : std_logic;
signal \pwm_setpoint_23_N_171_14\ : std_logic;
signal \pwm_setpoint_23_N_171_22\ : std_logic;
signal n9_adj_658 : std_logic;
signal pwm_setpoint_8 : std_logic;
signal n17_adj_665 : std_logic;
signal n19_adj_666 : std_logic;
signal n15178 : std_logic;
signal \n17_adj_665_cascade_\ : std_logic;
signal \pwm_setpoint_23_N_171_16\ : std_logic;
signal n15174 : std_logic;
signal \pwm_setpoint_23_N_171_17\ : std_logic;
signal pwm_setpoint_16 : std_logic;
signal pwm_setpoint_7 : std_logic;
signal \pwm_setpoint_23_N_171_10\ : std_logic;
signal pwm_setpoint_11 : std_logic;
signal n15204 : std_logic;
signal pwm_setpoint_17 : std_logic;
signal \n35_cascade_\ : std_logic;
signal n12_adj_661 : std_logic;
signal n1825 : std_logic;
signal \n1825_cascade_\ : std_logic;
signal n14520 : std_logic;
signal n1828 : std_logic;
signal n1830 : std_logic;
signal \n1752_cascade_\ : std_logic;
signal n1826 : std_logic;
signal n1824 : std_logic;
signal n1823 : std_logic;
signal \n1726_cascade_\ : std_logic;
signal \n14244_cascade_\ : std_logic;
signal \n14250_cascade_\ : std_logic;
signal n14254 : std_logic;
signal \n1721_cascade_\ : std_logic;
signal n1820 : std_logic;
signal n1827 : std_logic;
signal \n1722_cascade_\ : std_logic;
signal n1821 : std_logic;
signal \n1731_cascade_\ : std_logic;
signal n11991 : std_logic;
signal n1801 : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal n1800 : std_logic;
signal n12591 : std_logic;
signal n1732 : std_logic;
signal n1799 : std_logic;
signal n12592 : std_logic;
signal n1731 : std_logic;
signal n1798 : std_logic;
signal n12593 : std_logic;
signal n1797 : std_logic;
signal n12594 : std_logic;
signal n1796 : std_logic;
signal n12595 : std_logic;
signal n1795 : std_logic;
signal n12596 : std_logic;
signal n1794 : std_logic;
signal n12597 : std_logic;
signal n12598 : std_logic;
signal n1726 : std_logic;
signal n1793 : std_logic;
signal \bfn_12_21_0_\ : std_logic;
signal n1792 : std_logic;
signal n12599 : std_logic;
signal n1791 : std_logic;
signal n12600 : std_logic;
signal n1723 : std_logic;
signal n1790 : std_logic;
signal n12601 : std_logic;
signal n1722 : std_logic;
signal n1789 : std_logic;
signal n12602 : std_logic;
signal n1721 : std_logic;
signal n1788 : std_logic;
signal n12603 : std_logic;
signal n1720 : std_logic;
signal n1787 : std_logic;
signal n12604 : std_logic;
signal n12605 : std_logic;
signal n1818 : std_logic;
signal n10_adj_628 : std_logic;
signal n17 : std_logic;
signal n303 : std_logic;
signal n15 : std_logic;
signal encoder0_position_18 : std_logic;
signal n899 : std_logic;
signal n832 : std_logic;
signal n900 : std_logic;
signal n833 : std_logic;
signal \n932_cascade_\ : std_logic;
signal encoder0_position_25 : std_logic;
signal n8 : std_logic;
signal n41 : std_logic;
signal n901 : std_logic;
signal \n41_cascade_\ : std_logic;
signal \n933_cascade_\ : std_logic;
signal n10 : std_logic;
signal encoder0_position_23 : std_logic;
signal encoder0_position_24 : std_logic;
signal n9 : std_logic;
signal \n295_cascade_\ : std_logic;
signal \n11955_cascade_\ : std_logic;
signal n14460 : std_logic;
signal \n960_cascade_\ : std_logic;
signal n861 : std_logic;
signal n829 : std_logic;
signal n896 : std_logic;
signal \bfn_12_25_0_\ : std_logic;
signal n24_adj_552 : std_logic;
signal n12473 : std_logic;
signal n23_adj_553 : std_logic;
signal n12474 : std_logic;
signal n22_adj_554 : std_logic;
signal n12475 : std_logic;
signal n21_adj_555 : std_logic;
signal duty_4 : std_logic;
signal n12476 : std_logic;
signal n20_adj_556 : std_logic;
signal duty_5 : std_logic;
signal n12477 : std_logic;
signal n19_adj_557 : std_logic;
signal n12478 : std_logic;
signal n18_adj_558 : std_logic;
signal duty_7 : std_logic;
signal n12479 : std_logic;
signal n12480 : std_logic;
signal n17_adj_559 : std_logic;
signal duty_8 : std_logic;
signal \bfn_12_26_0_\ : std_logic;
signal n16_adj_560 : std_logic;
signal duty_9 : std_logic;
signal n12481 : std_logic;
signal n15_adj_561 : std_logic;
signal duty_10 : std_logic;
signal n12482 : std_logic;
signal n14_adj_562 : std_logic;
signal duty_11 : std_logic;
signal n12483 : std_logic;
signal n13_adj_563 : std_logic;
signal n12484 : std_logic;
signal n12_adj_564 : std_logic;
signal duty_13 : std_logic;
signal n12485 : std_logic;
signal n11_adj_565 : std_logic;
signal duty_14 : std_logic;
signal n12486 : std_logic;
signal n10_adj_566 : std_logic;
signal n12487 : std_logic;
signal n12488 : std_logic;
signal duty_16 : std_logic;
signal \bfn_12_27_0_\ : std_logic;
signal n8_adj_568 : std_logic;
signal n12489 : std_logic;
signal n7_adj_569 : std_logic;
signal n12490 : std_logic;
signal n6_adj_570 : std_logic;
signal n12491 : std_logic;
signal n5_adj_571 : std_logic;
signal n12492 : std_logic;
signal n4_adj_572 : std_logic;
signal n12493 : std_logic;
signal n3_adj_573 : std_logic;
signal n12494 : std_logic;
signal n2_adj_574 : std_logic;
signal n12495 : std_logic;
signal duty_17 : std_logic;
signal n8_adj_580 : std_logic;
signal duty_21 : std_logic;
signal n4_adj_576 : std_logic;
signal duty_18 : std_logic;
signal n7_adj_579 : std_logic;
signal \pwm_setpoint_23_N_171_19\ : std_logic;
signal \pwm_setpoint_23_N_171_20\ : std_logic;
signal \pwm_setpoint_23_N_171_0\ : std_logic;
signal duty_0 : std_logic;
signal pwm_setpoint_0 : std_logic;
signal duty_20 : std_logic;
signal n5_adj_577 : std_logic;
signal pwm_setpoint_22 : std_logic;
signal \n45_cascade_\ : std_logic;
signal pwm_setpoint_20 : std_logic;
signal \n41_adj_678_cascade_\ : std_logic;
signal n40_adj_677 : std_logic;
signal n45 : std_logic;
signal n15223 : std_logic;
signal n15165 : std_logic;
signal n15243 : std_logic;
signal duty_22 : std_logic;
signal n3_adj_575 : std_logic;
signal pwm_setpoint_19 : std_logic;
signal \n39_adj_676_cascade_\ : std_logic;
signal n15254 : std_logic;
signal pwm_setpoint_21 : std_logic;
signal \pwm_setpoint_23_N_171_12\ : std_logic;
signal n39_adj_676 : std_logic;
signal n41_adj_678 : std_logic;
signal n15091 : std_logic;
signal n4_adj_655 : std_logic;
signal pwm_setpoint_12 : std_logic;
signal n25_adj_670 : std_logic;
signal n15110 : std_logic;
signal n23_adj_668 : std_logic;
signal \n25_adj_670_cascade_\ : std_logic;
signal n43 : std_logic;
signal n15146 : std_logic;
signal n13_adj_662 : std_logic;
signal n15_adj_663 : std_logic;
signal n15229 : std_logic;
signal duty_12 : std_logic;
signal n13_adj_585 : std_logic;
signal \n31_adj_674_cascade_\ : std_logic;
signal n15230 : std_logic;
signal n15237 : std_logic;
signal \n15195_cascade_\ : std_logic;
signal n15241 : std_logic;
signal n15097 : std_logic;
signal n10_adj_659 : std_logic;
signal n30_adj_673 : std_logic;
signal n33_adj_675 : std_logic;
signal n15104 : std_logic;
signal n31_adj_674 : std_logic;
signal n35 : std_logic;
signal n15247 : std_logic;
signal \n15099_cascade_\ : std_logic;
signal n15220 : std_logic;
signal pwm_setpoint_18 : std_logic;
signal \n15257_cascade_\ : std_logic;
signal n37 : std_logic;
signal n15258 : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal n1700 : std_logic;
signal n12577 : std_logic;
signal n1699 : std_logic;
signal n12578 : std_logic;
signal n12579 : std_logic;
signal n12580 : std_logic;
signal n12581 : std_logic;
signal n12582 : std_logic;
signal n1694 : std_logic;
signal n12583 : std_logic;
signal n12584 : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal n12585 : std_logic;
signal n1691 : std_logic;
signal n12586 : std_logic;
signal n1690 : std_logic;
signal n12587 : std_logic;
signal n1689 : std_logic;
signal n12588 : std_logic;
signal n1688 : std_logic;
signal n12589 : std_logic;
signal n12590 : std_logic;
signal n1719 : std_logic;
signal n1695 : std_logic;
signal n1727 : std_logic;
signal n1696 : std_logic;
signal \n1653_cascade_\ : std_logic;
signal n1728 : std_logic;
signal n1697 : std_logic;
signal n1692 : std_logic;
signal n1724 : std_logic;
signal n1693_adj_614 : std_logic;
signal n1725 : std_logic;
signal n15611 : std_logic;
signal n1625_adj_605 : std_logic;
signal \n1625_adj_605_cascade_\ : std_logic;
signal n1698 : std_logic;
signal n1730 : std_logic;
signal \n1730_cascade_\ : std_logic;
signal n1729 : std_logic;
signal n14514 : std_logic;
signal n11_adj_629 : std_logic;
signal n1701 : std_logic;
signal n1653 : std_logic;
signal n1733 : std_logic;
signal n1752 : std_logic;
signal n15630 : std_logic;
signal n1621_adj_601 : std_logic;
signal \ENCODER0_B_N\ : std_logic;
signal encoder0_position_1 : std_logic;
signal n32_adj_650 : std_logic;
signal encoder0_position_16 : std_logic;
signal n17_adj_635 : std_logic;
signal \n1129_cascade_\ : std_logic;
signal \n11933_cascade_\ : std_logic;
signal \n13728_cascade_\ : std_logic;
signal \n1059_cascade_\ : std_logic;
signal \n1132_cascade_\ : std_logic;
signal n295 : std_logic;
signal n1001 : std_logic;
signal \bfn_13_24_0_\ : std_logic;
signal n933 : std_logic;
signal n1000 : std_logic;
signal n12507 : std_logic;
signal n932 : std_logic;
signal n999 : std_logic;
signal n12508 : std_logic;
signal n931 : std_logic;
signal n998 : std_logic;
signal n12509 : std_logic;
signal n930 : std_logic;
signal n997 : std_logic;
signal n12510 : std_logic;
signal n929 : std_logic;
signal n996 : std_logic;
signal n12511 : std_logic;
signal n928 : std_logic;
signal n995 : std_logic;
signal n12512 : std_logic;
signal n960 : std_logic;
signal n927 : std_logic;
signal n12513 : std_logic;
signal encoder0_position_scaled_0 : std_logic;
signal n25_adj_551 : std_logic;
signal \n11872_cascade_\ : std_logic;
signal \n14034_cascade_\ : std_logic;
signal \n14116_cascade_\ : std_logic;
signal n10_adj_598 : std_logic;
signal \pwm_setpoint_23_N_171_2\ : std_logic;
signal \pwm_setpoint_23_N_171_3\ : std_logic;
signal duty_3 : std_logic;
signal n10_adj_681 : std_logic;
signal \n16_adj_710_cascade_\ : std_logic;
signal n15_adj_711 : std_logic;
signal duty_2 : std_logic;
signal n23_adj_595 : std_logic;
signal duty_15 : std_logic;
signal \pwm_setpoint_23_N_171_15\ : std_logic;
signal pwm_setpoint_15 : std_logic;
signal \quad_counter0.a_new_0\ : std_logic;
signal \quad_counter0.b_new_0\ : std_logic;
signal a_new_1 : std_logic;
signal \quad_counter0.a_prev_N_543\ : std_logic;
signal \quad_counter0.b_new_1\ : std_logic;
signal \quad_counter0.debounce_cnt\ : std_logic;
signal \quad_counter0.a_prev_N_543_cascade_\ : std_logic;
signal b_prev : std_logic;
signal n15121 : std_logic;
signal \pwm_setpoint_23_N_171_6\ : std_logic;
signal pwm_setpoint_6 : std_logic;
signal pwm_setpoint_2 : std_logic;
signal pwm_setpoint_3 : std_logic;
signal duty_19 : std_logic;
signal n6_adj_578 : std_logic;
signal \PWM.n13991\ : std_logic;
signal n4_adj_599 : std_logic;
signal commutation_state_prev_1 : std_logic;
signal n5137 : std_logic;
signal dti : std_logic;
signal \n5201_cascade_\ : std_logic;
signal pwm_setpoint_13 : std_logic;
signal n27_adj_671 : std_logic;
signal \PWM.n17\ : std_logic;
signal \PWM.n26_cascade_\ : std_logic;
signal \PWM.n27\ : std_logic;
signal \PWM.n29_cascade_\ : std_logic;
signal \PWM.n28\ : std_logic;
signal commutation_state_prev_2 : std_logic;
signal h2 : std_logic;
signal h3 : std_logic;
signal h1 : std_logic;
signal n6_adj_721 : std_logic;
signal \commutation_state_7__N_261\ : std_logic;
signal pwm_setpoint_5 : std_logic;
signal n11_adj_660 : std_logic;
signal pwm_setpoint_14 : std_logic;
signal n29_adj_672 : std_logic;
signal n21_adj_667 : std_logic;
signal pwm_setpoint_10 : std_logic;
signal \n21_adj_667_cascade_\ : std_logic;
signal n6_adj_656 : std_logic;
signal n15203 : std_logic;
signal \n14420_cascade_\ : std_logic;
signal n1630_adj_610 : std_logic;
signal n1629_adj_609 : std_logic;
signal \n1630_adj_610_cascade_\ : std_logic;
signal n1624_adj_604 : std_logic;
signal n14502 : std_logic;
signal n1623_adj_603 : std_logic;
signal \n1624_adj_604_cascade_\ : std_logic;
signal n13748 : std_logic;
signal n14508 : std_logic;
signal n1627_adj_607 : std_logic;
signal \n1523_cascade_\ : std_logic;
signal n1622_adj_602 : std_logic;
signal n14426 : std_logic;
signal \n14428_cascade_\ : std_logic;
signal \n1554_cascade_\ : std_logic;
signal \n1427_cascade_\ : std_logic;
signal n1628_adj_608 : std_logic;
signal n11 : std_logic;
signal encoder0_position_22 : std_logic;
signal n1626_adj_606 : std_logic;
signal duty_6 : std_logic;
signal n19_adj_591 : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal n12541 : std_logic;
signal n12542 : std_logic;
signal n12543 : std_logic;
signal n12544 : std_logic;
signal n1396 : std_logic;
signal n12545 : std_logic;
signal n1395 : std_logic;
signal n12546 : std_logic;
signal n12547 : std_logic;
signal n12548 : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal n1392 : std_logic;
signal n12549 : std_logic;
signal n12550 : std_logic;
signal n12551 : std_logic;
signal n15553 : std_logic;
signal n1401 : std_logic;
signal n12019 : std_logic;
signal \n14406_cascade_\ : std_logic;
signal n14464 : std_logic;
signal \n1233_cascade_\ : std_logic;
signal n297 : std_logic;
signal n1201 : std_logic;
signal \bfn_14_23_0_\ : std_logic;
signal n1133 : std_logic;
signal n1200 : std_logic;
signal n12522 : std_logic;
signal n12523 : std_logic;
signal n1131 : std_logic;
signal n1198 : std_logic;
signal n12524 : std_logic;
signal n1130 : std_logic;
signal n1197 : std_logic;
signal n12525 : std_logic;
signal n12526 : std_logic;
signal n12527 : std_logic;
signal n12528 : std_logic;
signal n12529 : std_logic;
signal \bfn_14_24_0_\ : std_logic;
signal n12530 : std_logic;
signal n15522 : std_logic;
signal n13 : std_logic;
signal encoder0_position_20 : std_logic;
signal n1125 : std_logic;
signal \n20_adj_618_cascade_\ : std_logic;
signal n13197 : std_logic;
signal \n13197_cascade_\ : std_logic;
signal n24_adj_653 : std_logic;
signal \direction_N_342_cascade_\ : std_logic;
signal \direction_N_342\ : std_logic;
signal n13675 : std_logic;
signal \n23_adj_709_cascade_\ : std_logic;
signal n25_adj_707 : std_logic;
signal \direction_N_340\ : std_logic;
signal n24_adj_708 : std_logic;
signal n23_adj_654 : std_logic;
signal \pwm_setpoint_23_N_171_1\ : std_logic;
signal pwm_setpoint_1 : std_logic;
signal \n16_adj_679_cascade_\ : std_logic;
signal n15_adj_680 : std_logic;
signal n25_adj_652 : std_logic;
signal \n16_adj_619_cascade_\ : std_logic;
signal n22_adj_617 : std_logic;
signal n24_adj_616 : std_logic;
signal encoder0_position_scaled_16 : std_logic;
signal n9_adj_567 : std_logic;
signal duty_1 : std_logic;
signal n24_adj_596 : std_logic;
signal \pwm_setpoint_23__N_195\ : std_logic;
signal pwm_counter_0 : std_logic;
signal \bfn_14_28_0_\ : std_logic;
signal pwm_counter_1 : std_logic;
signal \PWM.n13022\ : std_logic;
signal pwm_counter_2 : std_logic;
signal \PWM.n13023\ : std_logic;
signal pwm_counter_3 : std_logic;
signal \PWM.n13024\ : std_logic;
signal pwm_counter_4 : std_logic;
signal \PWM.n13025\ : std_logic;
signal pwm_counter_5 : std_logic;
signal \PWM.n13026\ : std_logic;
signal pwm_counter_6 : std_logic;
signal \PWM.n13027\ : std_logic;
signal pwm_counter_7 : std_logic;
signal \PWM.n13028\ : std_logic;
signal \PWM.n13029\ : std_logic;
signal pwm_counter_8 : std_logic;
signal \bfn_14_29_0_\ : std_logic;
signal pwm_counter_9 : std_logic;
signal \PWM.n13030\ : std_logic;
signal pwm_counter_10 : std_logic;
signal \PWM.n13031\ : std_logic;
signal pwm_counter_11 : std_logic;
signal \PWM.n13032\ : std_logic;
signal pwm_counter_12 : std_logic;
signal \PWM.n13033\ : std_logic;
signal pwm_counter_13 : std_logic;
signal \PWM.n13034\ : std_logic;
signal pwm_counter_14 : std_logic;
signal \PWM.n13035\ : std_logic;
signal pwm_counter_15 : std_logic;
signal \PWM.n13036\ : std_logic;
signal \PWM.n13037\ : std_logic;
signal pwm_counter_16 : std_logic;
signal \bfn_14_30_0_\ : std_logic;
signal pwm_counter_17 : std_logic;
signal \PWM.n13038\ : std_logic;
signal pwm_counter_18 : std_logic;
signal \PWM.n13039\ : std_logic;
signal pwm_counter_19 : std_logic;
signal \PWM.n13040\ : std_logic;
signal pwm_counter_20 : std_logic;
signal \PWM.n13041\ : std_logic;
signal pwm_counter_21 : std_logic;
signal \PWM.n13042\ : std_logic;
signal pwm_counter_22 : std_logic;
signal \PWM.n13043\ : std_logic;
signal \PWM.n13044\ : std_logic;
signal \PWM.n13045\ : std_logic;
signal \bfn_14_31_0_\ : std_logic;
signal \PWM.n13046\ : std_logic;
signal \PWM.n13047\ : std_logic;
signal \PWM.n13048\ : std_logic;
signal \PWM.n13049\ : std_logic;
signal \PWM.n13050\ : std_logic;
signal \PWM.n13051\ : std_logic;
signal \PWM.n13052\ : std_logic;
signal \PWM.pwm_counter_31__N_407\ : std_logic;
signal pwm_counter_24 : std_logic;
signal pwm_counter_29 : std_logic;
signal pwm_counter_27 : std_logic;
signal pwm_counter_26 : std_logic;
signal pwm_counter_30 : std_logic;
signal pwm_counter_25 : std_logic;
signal \n12_adj_615_cascade_\ : std_logic;
signal pwm_counter_28 : std_logic;
signal n1631_adj_611 : std_logic;
signal n1554 : std_logic;
signal n1632_adj_612 : std_logic;
signal n302 : std_logic;
signal \n1632_adj_612_cascade_\ : std_logic;
signal n1633_adj_613 : std_logic;
signal n11919 : std_logic;
signal n1393 : std_logic;
signal \n1425_cascade_\ : std_logic;
signal n14484 : std_logic;
signal \n14490_cascade_\ : std_logic;
signal \n1455_cascade_\ : std_logic;
signal \n1531_cascade_\ : std_logic;
signal n11997 : std_logic;
signal n1455 : std_logic;
signal n1394 : std_logic;
signal n1391 : std_logic;
signal n299 : std_logic;
signal \n11925_cascade_\ : std_logic;
signal n1398 : std_logic;
signal \n1430_cascade_\ : std_logic;
signal n13739 : std_logic;
signal n13720 : std_logic;
signal n1400 : std_logic;
signal \n1356_cascade_\ : std_logic;
signal n1333 : std_logic;
signal \n1432_cascade_\ : std_logic;
signal n11923 : std_logic;
signal n1328 : std_logic;
signal \n1328_cascade_\ : std_logic;
signal n14414 : std_logic;
signal n1327 : std_logic;
signal n1331 : std_logic;
signal n1332 : std_logic;
signal n1399 : std_logic;
signal \n1332_cascade_\ : std_logic;
signal n1329 : std_logic;
signal n11927 : std_logic;
signal \n13723_cascade_\ : std_logic;
signal \n1257_cascade_\ : std_logic;
signal n1325 : std_logic;
signal n12 : std_logic;
signal encoder0_position_31 : std_logic;
signal n1326 : std_logic;
signal n1195 : std_logic;
signal \n1227_cascade_\ : std_logic;
signal n14476 : std_logic;
signal n1199 : std_logic;
signal n1132 : std_logic;
signal n1127 : std_logic;
signal n1194 : std_logic;
signal \n1127_cascade_\ : std_logic;
signal n1126 : std_logic;
signal n1193 : std_logic;
signal \n1225_cascade_\ : std_logic;
signal n1324 : std_logic;
signal n1129 : std_logic;
signal n1196 : std_logic;
signal n1158 : std_logic;
signal n1059 : std_logic;
signal n1128 : std_logic;
signal \bfn_15_25_0_\ : std_logic;
signal n1693 : std_logic;
signal encoder0_position_target_0 : std_logic;
signal n12449 : std_logic;
signal encoder0_position_target_1 : std_logic;
signal n12450 : std_logic;
signal encoder0_position_target_2 : std_logic;
signal n12451 : std_logic;
signal encoder0_position_target_3 : std_logic;
signal n12452 : std_logic;
signal encoder0_position_target_4 : std_logic;
signal n12453 : std_logic;
signal encoder0_position_target_5 : std_logic;
signal n12454 : std_logic;
signal encoder0_position_target_6 : std_logic;
signal n12455 : std_logic;
signal n12456 : std_logic;
signal encoder0_position_target_7 : std_logic;
signal \bfn_15_26_0_\ : std_logic;
signal encoder0_position_target_8 : std_logic;
signal n12457 : std_logic;
signal encoder0_position_target_9 : std_logic;
signal n12458 : std_logic;
signal encoder0_position_target_10 : std_logic;
signal n12459 : std_logic;
signal encoder0_position_target_11 : std_logic;
signal n12460 : std_logic;
signal encoder0_position_target_12 : std_logic;
signal n12461 : std_logic;
signal encoder0_position_target_13 : std_logic;
signal n12462 : std_logic;
signal encoder0_position_target_14 : std_logic;
signal n12463 : std_logic;
signal n12464 : std_logic;
signal encoder0_position_target_15 : std_logic;
signal \bfn_15_27_0_\ : std_logic;
signal encoder0_position_target_16 : std_logic;
signal n12465 : std_logic;
signal encoder0_position_target_17 : std_logic;
signal n12466 : std_logic;
signal encoder0_position_target_18 : std_logic;
signal n12467 : std_logic;
signal encoder0_position_target_19 : std_logic;
signal n12468 : std_logic;
signal encoder0_position_target_20 : std_logic;
signal n12469 : std_logic;
signal encoder0_position_target_21 : std_logic;
signal n12470 : std_logic;
signal encoder0_position_target_22 : std_logic;
signal n12471 : std_logic;
signal n12472 : std_logic;
signal direction_c : std_logic;
signal \bfn_15_28_0_\ : std_logic;
signal encoder0_position_target_23 : std_logic;
signal pwm_setpoint_23 : std_logic;
signal pwm_counter_23 : std_logic;
signal n15245 : std_logic;
signal pwm_counter_31 : std_logic;
signal n5180 : std_logic;
signal n5182 : std_logic;
signal duty_23 : std_logic;
signal n300 : std_logic;
signal n1501 : std_logic;
signal \bfn_16_17_0_\ : std_logic;
signal n1433 : std_logic;
signal n1500 : std_logic;
signal n12552 : std_logic;
signal n1432 : std_logic;
signal n1499 : std_logic;
signal n12553 : std_logic;
signal n1431 : std_logic;
signal n1498 : std_logic;
signal n12554 : std_logic;
signal n1430 : std_logic;
signal n1497 : std_logic;
signal n12555 : std_logic;
signal n1496 : std_logic;
signal n12556 : std_logic;
signal n1428 : std_logic;
signal n1495 : std_logic;
signal n12557 : std_logic;
signal n1427 : std_logic;
signal n1494 : std_logic;
signal n12558 : std_logic;
signal n12559 : std_logic;
signal n1426 : std_logic;
signal n1493 : std_logic;
signal \bfn_16_18_0_\ : std_logic;
signal n1425 : std_logic;
signal n1492 : std_logic;
signal n12560 : std_logic;
signal n1424 : std_logic;
signal n1491 : std_logic;
signal n12561 : std_logic;
signal n1423 : std_logic;
signal n1490 : std_logic;
signal n12562 : std_logic;
signal n15572 : std_logic;
signal n1422 : std_logic;
signal n12563 : std_logic;
signal n301 : std_logic;
signal n1601 : std_logic;
signal \bfn_16_19_0_\ : std_logic;
signal n1533 : std_logic;
signal n1600 : std_logic;
signal n12564 : std_logic;
signal n1532 : std_logic;
signal n1599 : std_logic;
signal n12565 : std_logic;
signal n1531 : std_logic;
signal n1598 : std_logic;
signal n12566 : std_logic;
signal n1530 : std_logic;
signal n1597 : std_logic;
signal n12567 : std_logic;
signal n1529 : std_logic;
signal n1596 : std_logic;
signal n12568 : std_logic;
signal n1528 : std_logic;
signal n1595 : std_logic;
signal n12569 : std_logic;
signal n1527 : std_logic;
signal n1594 : std_logic;
signal n12570 : std_logic;
signal n12571 : std_logic;
signal n1526 : std_logic;
signal n1593 : std_logic;
signal \bfn_16_20_0_\ : std_logic;
signal n1525 : std_logic;
signal n1592 : std_logic;
signal n12572 : std_logic;
signal n1524 : std_logic;
signal n1591 : std_logic;
signal n12573 : std_logic;
signal n1523 : std_logic;
signal n1590 : std_logic;
signal n12574 : std_logic;
signal n1522 : std_logic;
signal n1589 : std_logic;
signal n12575 : std_logic;
signal n1521 : std_logic;
signal n15591 : std_logic;
signal n12576 : std_logic;
signal n1620_adj_600 : std_logic;
signal encoder0_position_21 : std_logic;
signal n12_adj_630 : std_logic;
signal n1397 : std_logic;
signal n1356 : std_logic;
signal n1429 : std_logic;
signal n298 : std_logic;
signal n1301 : std_logic;
signal \bfn_16_21_0_\ : std_logic;
signal n1233 : std_logic;
signal n1300 : std_logic;
signal n12531 : std_logic;
signal n1232 : std_logic;
signal n1299 : std_logic;
signal n12532 : std_logic;
signal n12533 : std_logic;
signal n1230 : std_logic;
signal n1297 : std_logic;
signal n12534 : std_logic;
signal n1229 : std_logic;
signal n1296 : std_logic;
signal n12535 : std_logic;
signal n1228 : std_logic;
signal n1295 : std_logic;
signal n12536 : std_logic;
signal n1227 : std_logic;
signal n1294 : std_logic;
signal n12537 : std_logic;
signal n12538 : std_logic;
signal n1226 : std_logic;
signal n1293 : std_logic;
signal \bfn_16_22_0_\ : std_logic;
signal n1225 : std_logic;
signal n1292 : std_logic;
signal n12539 : std_logic;
signal n15537 : std_logic;
signal n1224 : std_logic;
signal n12540 : std_logic;
signal n1323 : std_logic;
signal n1298 : std_logic;
signal n1231 : std_logic;
signal n1257 : std_logic;
signal n1330 : std_logic;
signal n296 : std_logic;
signal n1101 : std_logic;
signal \bfn_16_23_0_\ : std_logic;
signal n1033 : std_logic;
signal n1100 : std_logic;
signal n12514 : std_logic;
signal n1032 : std_logic;
signal n1099 : std_logic;
signal n12515 : std_logic;
signal n1031 : std_logic;
signal n1098 : std_logic;
signal n12516 : std_logic;
signal n1030 : std_logic;
signal n1097 : std_logic;
signal n12517 : std_logic;
signal n1029 : std_logic;
signal n1096 : std_logic;
signal n12518 : std_logic;
signal n1028 : std_logic;
signal n1095 : std_logic;
signal n12519 : std_logic;
signal n1027 : std_logic;
signal n1094 : std_logic;
signal n12520 : std_logic;
signal n12521 : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal n1026 : std_logic;
signal \bfn_16_24_0_\ : std_logic;
signal n1093 : std_logic;
signal sweep_counter_0 : std_logic;
signal \bfn_16_25_0_\ : std_logic;
signal sweep_counter_1 : std_logic;
signal n13053 : std_logic;
signal sweep_counter_2 : std_logic;
signal n13054 : std_logic;
signal sweep_counter_3 : std_logic;
signal n13055 : std_logic;
signal sweep_counter_4 : std_logic;
signal n13056 : std_logic;
signal sweep_counter_5 : std_logic;
signal n13057 : std_logic;
signal sweep_counter_6 : std_logic;
signal n13058 : std_logic;
signal sweep_counter_7 : std_logic;
signal n13059 : std_logic;
signal n13060 : std_logic;
signal \bfn_16_26_0_\ : std_logic;
signal sweep_counter_9 : std_logic;
signal n13061 : std_logic;
signal sweep_counter_10 : std_logic;
signal n13062 : std_logic;
signal sweep_counter_11 : std_logic;
signal n13063 : std_logic;
signal n13064 : std_logic;
signal n13065 : std_logic;
signal n13066 : std_logic;
signal sweep_counter_15 : std_logic;
signal n13067 : std_logic;
signal n13068 : std_logic;
signal sweep_counter_16 : std_logic;
signal \bfn_16_27_0_\ : std_logic;
signal n13069 : std_logic;
signal n5215 : std_logic;
signal sweep_counter_8 : std_logic;
signal sweep_counter_14 : std_logic;
signal sweep_counter_13 : std_logic;
signal sweep_counter_17 : std_logic;
signal \n6_adj_712_cascade_\ : std_logic;
signal sweep_counter_12 : std_logic;
signal n13968 : std_logic;
signal \GHC\ : std_logic;
signal \INHC_c_0\ : std_logic;
signal \GHB\ : std_logic;
signal \INHB_c_0\ : std_logic;
signal \INLA_c_0\ : std_logic;
signal \INLB_c_0\ : std_logic;
signal commutation_state_0 : std_logic;
signal commutation_state_2 : std_logic;
signal dir : std_logic;
signal commutation_state_1 : std_logic;
signal \INLC_c_0\ : std_logic;
signal \CLK_N\ : std_logic;
signal n5201 : std_logic;
signal n5253 : std_logic;
signal \GHA\ : std_logic;
signal pwm_out : std_logic;
signal \INHA_c_0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CS_CLK_wire\ : std_logic;
signal \CS_wire\ : std_logic;
signal \DE_wire\ : std_logic;
signal \ENCODER0_A_wire\ : std_logic;
signal \ENCODER0_B_wire\ : std_logic;
signal \INHA_wire\ : std_logic;
signal \INHB_wire\ : std_logic;
signal \INHC_wire\ : std_logic;
signal \INLA_wire\ : std_logic;
signal \INLB_wire\ : std_logic;
signal \INLC_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \NEOPXL_wire\ : std_logic;
signal \TX_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \HALL1_wire\ : std_logic;
signal \HALL2_wire\ : std_logic;
signal \HALL3_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    CS_CLK <= \CS_CLK_wire\;
    CS <= \CS_wire\;
    DE <= \DE_wire\;
    \ENCODER0_A_wire\ <= ENCODER0_A;
    \ENCODER0_B_wire\ <= ENCODER0_B;
    INHA <= \INHA_wire\;
    INHB <= \INHB_wire\;
    INHC <= \INHC_wire\;
    INLA <= \INLA_wire\;
    INLB <= \INLB_wire\;
    INLC <= \INLC_wire\;
    LED <= \LED_wire\;
    NEOPXL <= \NEOPXL_wire\;
    TX <= \TX_wire\;
    USBPU <= \USBPU_wire\;
    \HALL1_wire\ <= HALL1;
    \HALL2_wire\ <= HALL2;
    \HALL3_wire\ <= HALL3;
    \CLK_wire\ <= CLK;

    \CS_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56752\,
            DIN => \N__56751\,
            DOUT => \N__56750\,
            PACKAGEPIN => \CS_CLK_wire\
        );

    \CS_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56752\,
            PADOUT => \N__56751\,
            PADIN => \N__56750\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \CS_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56743\,
            DIN => \N__56742\,
            DOUT => \N__56741\,
            PACKAGEPIN => \CS_wire\
        );

    \CS_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56743\,
            PADOUT => \N__56742\,
            PADIN => \N__56741\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \DE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56734\,
            DIN => \N__56733\,
            DOUT => \N__56732\,
            PACKAGEPIN => \DE_wire\
        );

    \DE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56734\,
            PADOUT => \N__56733\,
            PADIN => \N__56732\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \ENCODER0_A_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56725\,
            DIN => \N__56724\,
            DOUT => \N__56723\,
            PACKAGEPIN => \ENCODER0_A_wire\
        );

    \ENCODER0_A_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56725\,
            PADOUT => \N__56724\,
            PADIN => \N__56723\,
            CLOCKENABLE => 'H',
            DIN0 => \ENCODER0_A_N\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \ENCODER0_B_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56716\,
            DIN => \N__56715\,
            DOUT => \N__56714\,
            PACKAGEPIN => \ENCODER0_B_wire\
        );

    \ENCODER0_B_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56716\,
            PADOUT => \N__56715\,
            PADIN => \N__56714\,
            CLOCKENABLE => 'H',
            DIN0 => \ENCODER0_B_N\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHA_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56707\,
            DIN => \N__56706\,
            DOUT => \N__56705\,
            PACKAGEPIN => \INHA_wire\
        );

    \INHA_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56707\,
            PADOUT => \N__56706\,
            PADIN => \N__56705\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__55974\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHB_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56698\,
            DIN => \N__56697\,
            DOUT => \N__56696\,
            PACKAGEPIN => \INHB_wire\
        );

    \INHB_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56698\,
            PADOUT => \N__56697\,
            PADIN => \N__56696\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__56565\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56689\,
            DIN => \N__56688\,
            DOUT => \N__56687\,
            PACKAGEPIN => \INHC_wire\
        );

    \INHC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56689\,
            PADOUT => \N__56688\,
            PADIN => \N__56687\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__55728\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLA_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56680\,
            DIN => \N__56679\,
            DOUT => \N__56678\,
            PACKAGEPIN => \INLA_wire\
        );

    \INLA_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56680\,
            PADOUT => \N__56679\,
            PADIN => \N__56678\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__56553\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLB_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56671\,
            DIN => \N__56670\,
            DOUT => \N__56669\,
            PACKAGEPIN => \INLB_wire\
        );

    \INLB_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56671\,
            PADOUT => \N__56670\,
            PADIN => \N__56669\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__56538\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56662\,
            DIN => \N__56661\,
            DOUT => \N__56660\,
            PACKAGEPIN => \INLC_wire\
        );

    \INLC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56662\,
            PADOUT => \N__56661\,
            PADIN => \N__56660\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__56277\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56653\,
            DIN => \N__56652\,
            DOUT => \N__56651\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56653\,
            PADOUT => \N__56652\,
            PADIN => \N__56651\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__39138\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \NEOPXL_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56644\,
            DIN => \N__56643\,
            DOUT => \N__56642\,
            PACKAGEPIN => \NEOPXL_wire\
        );

    \NEOPXL_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56644\,
            PADOUT => \N__56643\,
            PADIN => \N__56642\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \TX_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56635\,
            DIN => \N__56634\,
            DOUT => \N__56633\,
            PACKAGEPIN => \TX_wire\
        );

    \TX_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56635\,
            PADOUT => \N__56634\,
            PADIN => \N__56633\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56626\,
            DIN => \N__56625\,
            DOUT => \N__56624\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56626\,
            PADOUT => \N__56625\,
            PADIN => \N__56624\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall1_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__56617\,
            DIN => \N__56616\,
            DOUT => \N__56615\,
            PACKAGEPIN => \HALL1_wire\
        );

    \hall1_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56617\,
            PADOUT => \N__56616\,
            PADIN => \N__56615\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => \debounce.reg_A_2\,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => \N__56204\,
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall2_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__56608\,
            DIN => \N__56607\,
            DOUT => \N__56606\,
            PACKAGEPIN => \HALL2_wire\
        );

    \hall2_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56608\,
            PADOUT => \N__56607\,
            PADIN => \N__56606\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => \debounce.reg_A_1\,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => \N__56200\,
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hall3_input_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__56599\,
            DIN => \N__56598\,
            DOUT => \N__56597\,
            PACKAGEPIN => \HALL3_wire\
        );

    \hall3_input_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56599\,
            PADOUT => \N__56598\,
            PADIN => \N__56597\,
            CLOCKENABLE => \VCCG0\,
            DIN0 => \debounce.reg_A_0\,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => \GNDG0\,
            INPUTCLK => \N__56200\,
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__56590\,
            DIN => \N__56589\,
            DOUT => \N__56588\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__56590\,
            PADOUT => \N__56589\,
            PADIN => \N__56588\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__13452\ : InMux
    port map (
            O => \N__56571\,
            I => \N__56568\
        );

    \I__13451\ : LocalMux
    port map (
            O => \N__56568\,
            I => \GHB\
        );

    \I__13450\ : IoInMux
    port map (
            O => \N__56565\,
            I => \N__56562\
        );

    \I__13449\ : LocalMux
    port map (
            O => \N__56562\,
            I => \N__56559\
        );

    \I__13448\ : Span12Mux_s0_v
    port map (
            O => \N__56559\,
            I => \N__56556\
        );

    \I__13447\ : Odrv12
    port map (
            O => \N__56556\,
            I => \INHB_c_0\
        );

    \I__13446\ : IoInMux
    port map (
            O => \N__56553\,
            I => \N__56550\
        );

    \I__13445\ : LocalMux
    port map (
            O => \N__56550\,
            I => \N__56547\
        );

    \I__13444\ : Span4Mux_s1_v
    port map (
            O => \N__56547\,
            I => \N__56544\
        );

    \I__13443\ : Span4Mux_h
    port map (
            O => \N__56544\,
            I => \N__56541\
        );

    \I__13442\ : Odrv4
    port map (
            O => \N__56541\,
            I => \INLA_c_0\
        );

    \I__13441\ : IoInMux
    port map (
            O => \N__56538\,
            I => \N__56535\
        );

    \I__13440\ : LocalMux
    port map (
            O => \N__56535\,
            I => \N__56532\
        );

    \I__13439\ : Span4Mux_s1_v
    port map (
            O => \N__56532\,
            I => \N__56529\
        );

    \I__13438\ : Span4Mux_h
    port map (
            O => \N__56529\,
            I => \N__56526\
        );

    \I__13437\ : Odrv4
    port map (
            O => \N__56526\,
            I => \INLB_c_0\
        );

    \I__13436\ : InMux
    port map (
            O => \N__56523\,
            I => \N__56497\
        );

    \I__13435\ : InMux
    port map (
            O => \N__56522\,
            I => \N__56497\
        );

    \I__13434\ : InMux
    port map (
            O => \N__56521\,
            I => \N__56497\
        );

    \I__13433\ : InMux
    port map (
            O => \N__56520\,
            I => \N__56497\
        );

    \I__13432\ : InMux
    port map (
            O => \N__56519\,
            I => \N__56497\
        );

    \I__13431\ : InMux
    port map (
            O => \N__56518\,
            I => \N__56494\
        );

    \I__13430\ : InMux
    port map (
            O => \N__56517\,
            I => \N__56491\
        );

    \I__13429\ : InMux
    port map (
            O => \N__56516\,
            I => \N__56488\
        );

    \I__13428\ : InMux
    port map (
            O => \N__56515\,
            I => \N__56485\
        );

    \I__13427\ : InMux
    port map (
            O => \N__56514\,
            I => \N__56476\
        );

    \I__13426\ : InMux
    port map (
            O => \N__56513\,
            I => \N__56476\
        );

    \I__13425\ : InMux
    port map (
            O => \N__56512\,
            I => \N__56476\
        );

    \I__13424\ : InMux
    port map (
            O => \N__56511\,
            I => \N__56476\
        );

    \I__13423\ : InMux
    port map (
            O => \N__56510\,
            I => \N__56469\
        );

    \I__13422\ : InMux
    port map (
            O => \N__56509\,
            I => \N__56469\
        );

    \I__13421\ : InMux
    port map (
            O => \N__56508\,
            I => \N__56469\
        );

    \I__13420\ : LocalMux
    port map (
            O => \N__56497\,
            I => \N__56466\
        );

    \I__13419\ : LocalMux
    port map (
            O => \N__56494\,
            I => \N__56461\
        );

    \I__13418\ : LocalMux
    port map (
            O => \N__56491\,
            I => \N__56461\
        );

    \I__13417\ : LocalMux
    port map (
            O => \N__56488\,
            I => \N__56450\
        );

    \I__13416\ : LocalMux
    port map (
            O => \N__56485\,
            I => \N__56450\
        );

    \I__13415\ : LocalMux
    port map (
            O => \N__56476\,
            I => \N__56450\
        );

    \I__13414\ : LocalMux
    port map (
            O => \N__56469\,
            I => \N__56450\
        );

    \I__13413\ : Span12Mux_v
    port map (
            O => \N__56466\,
            I => \N__56450\
        );

    \I__13412\ : Span4Mux_h
    port map (
            O => \N__56461\,
            I => \N__56447\
        );

    \I__13411\ : Odrv12
    port map (
            O => \N__56450\,
            I => commutation_state_0
        );

    \I__13410\ : Odrv4
    port map (
            O => \N__56447\,
            I => commutation_state_0
        );

    \I__13409\ : CascadeMux
    port map (
            O => \N__56442\,
            I => \N__56436\
        );

    \I__13408\ : CascadeMux
    port map (
            O => \N__56441\,
            I => \N__56433\
        );

    \I__13407\ : CascadeMux
    port map (
            O => \N__56440\,
            I => \N__56428\
        );

    \I__13406\ : CascadeMux
    port map (
            O => \N__56439\,
            I => \N__56425\
        );

    \I__13405\ : InMux
    port map (
            O => \N__56436\,
            I => \N__56416\
        );

    \I__13404\ : InMux
    port map (
            O => \N__56433\,
            I => \N__56416\
        );

    \I__13403\ : InMux
    port map (
            O => \N__56432\,
            I => \N__56416\
        );

    \I__13402\ : InMux
    port map (
            O => \N__56431\,
            I => \N__56416\
        );

    \I__13401\ : InMux
    port map (
            O => \N__56428\,
            I => \N__56413\
        );

    \I__13400\ : InMux
    port map (
            O => \N__56425\,
            I => \N__56410\
        );

    \I__13399\ : LocalMux
    port map (
            O => \N__56416\,
            I => \N__56407\
        );

    \I__13398\ : LocalMux
    port map (
            O => \N__56413\,
            I => \N__56398\
        );

    \I__13397\ : LocalMux
    port map (
            O => \N__56410\,
            I => \N__56398\
        );

    \I__13396\ : Span4Mux_s2_v
    port map (
            O => \N__56407\,
            I => \N__56395\
        );

    \I__13395\ : CascadeMux
    port map (
            O => \N__56406\,
            I => \N__56392\
        );

    \I__13394\ : CascadeMux
    port map (
            O => \N__56405\,
            I => \N__56389\
        );

    \I__13393\ : InMux
    port map (
            O => \N__56404\,
            I => \N__56384\
        );

    \I__13392\ : InMux
    port map (
            O => \N__56403\,
            I => \N__56384\
        );

    \I__13391\ : Span4Mux_s2_v
    port map (
            O => \N__56398\,
            I => \N__56381\
        );

    \I__13390\ : Span4Mux_h
    port map (
            O => \N__56395\,
            I => \N__56378\
        );

    \I__13389\ : InMux
    port map (
            O => \N__56392\,
            I => \N__56373\
        );

    \I__13388\ : InMux
    port map (
            O => \N__56389\,
            I => \N__56373\
        );

    \I__13387\ : LocalMux
    port map (
            O => \N__56384\,
            I => commutation_state_2
        );

    \I__13386\ : Odrv4
    port map (
            O => \N__56381\,
            I => commutation_state_2
        );

    \I__13385\ : Odrv4
    port map (
            O => \N__56378\,
            I => commutation_state_2
        );

    \I__13384\ : LocalMux
    port map (
            O => \N__56373\,
            I => commutation_state_2
        );

    \I__13383\ : CascadeMux
    port map (
            O => \N__56364\,
            I => \N__56360\
        );

    \I__13382\ : CascadeMux
    port map (
            O => \N__56363\,
            I => \N__56356\
        );

    \I__13381\ : InMux
    port map (
            O => \N__56360\,
            I => \N__56344\
        );

    \I__13380\ : InMux
    port map (
            O => \N__56359\,
            I => \N__56344\
        );

    \I__13379\ : InMux
    port map (
            O => \N__56356\,
            I => \N__56344\
        );

    \I__13378\ : InMux
    port map (
            O => \N__56355\,
            I => \N__56344\
        );

    \I__13377\ : InMux
    port map (
            O => \N__56354\,
            I => \N__56341\
        );

    \I__13376\ : InMux
    port map (
            O => \N__56353\,
            I => \N__56338\
        );

    \I__13375\ : LocalMux
    port map (
            O => \N__56344\,
            I => \N__56333\
        );

    \I__13374\ : LocalMux
    port map (
            O => \N__56341\,
            I => \N__56333\
        );

    \I__13373\ : LocalMux
    port map (
            O => \N__56338\,
            I => dir
        );

    \I__13372\ : Odrv12
    port map (
            O => \N__56333\,
            I => dir
        );

    \I__13371\ : InMux
    port map (
            O => \N__56328\,
            I => \N__56316\
        );

    \I__13370\ : InMux
    port map (
            O => \N__56327\,
            I => \N__56307\
        );

    \I__13369\ : InMux
    port map (
            O => \N__56326\,
            I => \N__56307\
        );

    \I__13368\ : InMux
    port map (
            O => \N__56325\,
            I => \N__56307\
        );

    \I__13367\ : InMux
    port map (
            O => \N__56324\,
            I => \N__56307\
        );

    \I__13366\ : InMux
    port map (
            O => \N__56323\,
            I => \N__56304\
        );

    \I__13365\ : InMux
    port map (
            O => \N__56322\,
            I => \N__56297\
        );

    \I__13364\ : InMux
    port map (
            O => \N__56321\,
            I => \N__56297\
        );

    \I__13363\ : InMux
    port map (
            O => \N__56320\,
            I => \N__56297\
        );

    \I__13362\ : InMux
    port map (
            O => \N__56319\,
            I => \N__56294\
        );

    \I__13361\ : LocalMux
    port map (
            O => \N__56316\,
            I => \N__56287\
        );

    \I__13360\ : LocalMux
    port map (
            O => \N__56307\,
            I => \N__56287\
        );

    \I__13359\ : LocalMux
    port map (
            O => \N__56304\,
            I => \N__56287\
        );

    \I__13358\ : LocalMux
    port map (
            O => \N__56297\,
            I => \N__56284\
        );

    \I__13357\ : LocalMux
    port map (
            O => \N__56294\,
            I => commutation_state_1
        );

    \I__13356\ : Odrv12
    port map (
            O => \N__56287\,
            I => commutation_state_1
        );

    \I__13355\ : Odrv4
    port map (
            O => \N__56284\,
            I => commutation_state_1
        );

    \I__13354\ : IoInMux
    port map (
            O => \N__56277\,
            I => \N__56274\
        );

    \I__13353\ : LocalMux
    port map (
            O => \N__56274\,
            I => \N__56271\
        );

    \I__13352\ : Span12Mux_s6_v
    port map (
            O => \N__56271\,
            I => \N__56268\
        );

    \I__13351\ : Span12Mux_h
    port map (
            O => \N__56268\,
            I => \N__56265\
        );

    \I__13350\ : Odrv12
    port map (
            O => \N__56265\,
            I => \INLC_c_0\
        );

    \I__13349\ : ClkMux
    port map (
            O => \N__56262\,
            I => \N__56070\
        );

    \I__13348\ : ClkMux
    port map (
            O => \N__56261\,
            I => \N__56070\
        );

    \I__13347\ : ClkMux
    port map (
            O => \N__56260\,
            I => \N__56070\
        );

    \I__13346\ : ClkMux
    port map (
            O => \N__56259\,
            I => \N__56070\
        );

    \I__13345\ : ClkMux
    port map (
            O => \N__56258\,
            I => \N__56070\
        );

    \I__13344\ : ClkMux
    port map (
            O => \N__56257\,
            I => \N__56070\
        );

    \I__13343\ : ClkMux
    port map (
            O => \N__56256\,
            I => \N__56070\
        );

    \I__13342\ : ClkMux
    port map (
            O => \N__56255\,
            I => \N__56070\
        );

    \I__13341\ : ClkMux
    port map (
            O => \N__56254\,
            I => \N__56070\
        );

    \I__13340\ : ClkMux
    port map (
            O => \N__56253\,
            I => \N__56070\
        );

    \I__13339\ : ClkMux
    port map (
            O => \N__56252\,
            I => \N__56070\
        );

    \I__13338\ : ClkMux
    port map (
            O => \N__56251\,
            I => \N__56070\
        );

    \I__13337\ : ClkMux
    port map (
            O => \N__56250\,
            I => \N__56070\
        );

    \I__13336\ : ClkMux
    port map (
            O => \N__56249\,
            I => \N__56070\
        );

    \I__13335\ : ClkMux
    port map (
            O => \N__56248\,
            I => \N__56070\
        );

    \I__13334\ : ClkMux
    port map (
            O => \N__56247\,
            I => \N__56070\
        );

    \I__13333\ : ClkMux
    port map (
            O => \N__56246\,
            I => \N__56070\
        );

    \I__13332\ : ClkMux
    port map (
            O => \N__56245\,
            I => \N__56070\
        );

    \I__13331\ : ClkMux
    port map (
            O => \N__56244\,
            I => \N__56070\
        );

    \I__13330\ : ClkMux
    port map (
            O => \N__56243\,
            I => \N__56070\
        );

    \I__13329\ : ClkMux
    port map (
            O => \N__56242\,
            I => \N__56070\
        );

    \I__13328\ : ClkMux
    port map (
            O => \N__56241\,
            I => \N__56070\
        );

    \I__13327\ : ClkMux
    port map (
            O => \N__56240\,
            I => \N__56070\
        );

    \I__13326\ : ClkMux
    port map (
            O => \N__56239\,
            I => \N__56070\
        );

    \I__13325\ : ClkMux
    port map (
            O => \N__56238\,
            I => \N__56070\
        );

    \I__13324\ : ClkMux
    port map (
            O => \N__56237\,
            I => \N__56070\
        );

    \I__13323\ : ClkMux
    port map (
            O => \N__56236\,
            I => \N__56070\
        );

    \I__13322\ : ClkMux
    port map (
            O => \N__56235\,
            I => \N__56070\
        );

    \I__13321\ : ClkMux
    port map (
            O => \N__56234\,
            I => \N__56070\
        );

    \I__13320\ : ClkMux
    port map (
            O => \N__56233\,
            I => \N__56070\
        );

    \I__13319\ : ClkMux
    port map (
            O => \N__56232\,
            I => \N__56070\
        );

    \I__13318\ : ClkMux
    port map (
            O => \N__56231\,
            I => \N__56070\
        );

    \I__13317\ : ClkMux
    port map (
            O => \N__56230\,
            I => \N__56070\
        );

    \I__13316\ : ClkMux
    port map (
            O => \N__56229\,
            I => \N__56070\
        );

    \I__13315\ : ClkMux
    port map (
            O => \N__56228\,
            I => \N__56070\
        );

    \I__13314\ : ClkMux
    port map (
            O => \N__56227\,
            I => \N__56070\
        );

    \I__13313\ : ClkMux
    port map (
            O => \N__56226\,
            I => \N__56070\
        );

    \I__13312\ : ClkMux
    port map (
            O => \N__56225\,
            I => \N__56070\
        );

    \I__13311\ : ClkMux
    port map (
            O => \N__56224\,
            I => \N__56070\
        );

    \I__13310\ : ClkMux
    port map (
            O => \N__56223\,
            I => \N__56070\
        );

    \I__13309\ : ClkMux
    port map (
            O => \N__56222\,
            I => \N__56070\
        );

    \I__13308\ : ClkMux
    port map (
            O => \N__56221\,
            I => \N__56070\
        );

    \I__13307\ : ClkMux
    port map (
            O => \N__56220\,
            I => \N__56070\
        );

    \I__13306\ : ClkMux
    port map (
            O => \N__56219\,
            I => \N__56070\
        );

    \I__13305\ : ClkMux
    port map (
            O => \N__56218\,
            I => \N__56070\
        );

    \I__13304\ : ClkMux
    port map (
            O => \N__56217\,
            I => \N__56070\
        );

    \I__13303\ : ClkMux
    port map (
            O => \N__56216\,
            I => \N__56070\
        );

    \I__13302\ : ClkMux
    port map (
            O => \N__56215\,
            I => \N__56070\
        );

    \I__13301\ : ClkMux
    port map (
            O => \N__56214\,
            I => \N__56070\
        );

    \I__13300\ : ClkMux
    port map (
            O => \N__56213\,
            I => \N__56070\
        );

    \I__13299\ : ClkMux
    port map (
            O => \N__56212\,
            I => \N__56070\
        );

    \I__13298\ : ClkMux
    port map (
            O => \N__56211\,
            I => \N__56070\
        );

    \I__13297\ : ClkMux
    port map (
            O => \N__56210\,
            I => \N__56070\
        );

    \I__13296\ : ClkMux
    port map (
            O => \N__56209\,
            I => \N__56070\
        );

    \I__13295\ : ClkMux
    port map (
            O => \N__56208\,
            I => \N__56070\
        );

    \I__13294\ : ClkMux
    port map (
            O => \N__56207\,
            I => \N__56070\
        );

    \I__13293\ : ClkMux
    port map (
            O => \N__56206\,
            I => \N__56070\
        );

    \I__13292\ : ClkMux
    port map (
            O => \N__56205\,
            I => \N__56070\
        );

    \I__13291\ : ClkMux
    port map (
            O => \N__56204\,
            I => \N__56070\
        );

    \I__13290\ : ClkMux
    port map (
            O => \N__56203\,
            I => \N__56070\
        );

    \I__13289\ : ClkMux
    port map (
            O => \N__56202\,
            I => \N__56070\
        );

    \I__13288\ : ClkMux
    port map (
            O => \N__56201\,
            I => \N__56070\
        );

    \I__13287\ : ClkMux
    port map (
            O => \N__56200\,
            I => \N__56070\
        );

    \I__13286\ : ClkMux
    port map (
            O => \N__56199\,
            I => \N__56070\
        );

    \I__13285\ : GlobalMux
    port map (
            O => \N__56070\,
            I => \N__56067\
        );

    \I__13284\ : gio2CtrlBuf
    port map (
            O => \N__56067\,
            I => \CLK_N\
        );

    \I__13283\ : CEMux
    port map (
            O => \N__56064\,
            I => \N__56060\
        );

    \I__13282\ : CEMux
    port map (
            O => \N__56063\,
            I => \N__56057\
        );

    \I__13281\ : LocalMux
    port map (
            O => \N__56060\,
            I => \N__56053\
        );

    \I__13280\ : LocalMux
    port map (
            O => \N__56057\,
            I => \N__56050\
        );

    \I__13279\ : CEMux
    port map (
            O => \N__56056\,
            I => \N__56047\
        );

    \I__13278\ : Span4Mux_h
    port map (
            O => \N__56053\,
            I => \N__56040\
        );

    \I__13277\ : Span4Mux_h
    port map (
            O => \N__56050\,
            I => \N__56040\
        );

    \I__13276\ : LocalMux
    port map (
            O => \N__56047\,
            I => \N__56040\
        );

    \I__13275\ : Span4Mux_h
    port map (
            O => \N__56040\,
            I => \N__56037\
        );

    \I__13274\ : Odrv4
    port map (
            O => \N__56037\,
            I => n5201
        );

    \I__13273\ : SRMux
    port map (
            O => \N__56034\,
            I => \N__56031\
        );

    \I__13272\ : LocalMux
    port map (
            O => \N__56031\,
            I => \N__56026\
        );

    \I__13271\ : SRMux
    port map (
            O => \N__56030\,
            I => \N__56023\
        );

    \I__13270\ : SRMux
    port map (
            O => \N__56029\,
            I => \N__56020\
        );

    \I__13269\ : Span4Mux_h
    port map (
            O => \N__56026\,
            I => \N__56015\
        );

    \I__13268\ : LocalMux
    port map (
            O => \N__56023\,
            I => \N__56015\
        );

    \I__13267\ : LocalMux
    port map (
            O => \N__56020\,
            I => \N__56012\
        );

    \I__13266\ : Span4Mux_h
    port map (
            O => \N__56015\,
            I => \N__56009\
        );

    \I__13265\ : Span12Mux_s3_v
    port map (
            O => \N__56012\,
            I => \N__56006\
        );

    \I__13264\ : Odrv4
    port map (
            O => \N__56009\,
            I => n5253
        );

    \I__13263\ : Odrv12
    port map (
            O => \N__56006\,
            I => n5253
        );

    \I__13262\ : InMux
    port map (
            O => \N__56001\,
            I => \N__55998\
        );

    \I__13261\ : LocalMux
    port map (
            O => \N__55998\,
            I => \GHA\
        );

    \I__13260\ : InMux
    port map (
            O => \N__55995\,
            I => \N__55990\
        );

    \I__13259\ : InMux
    port map (
            O => \N__55994\,
            I => \N__55985\
        );

    \I__13258\ : InMux
    port map (
            O => \N__55993\,
            I => \N__55985\
        );

    \I__13257\ : LocalMux
    port map (
            O => \N__55990\,
            I => \N__55980\
        );

    \I__13256\ : LocalMux
    port map (
            O => \N__55985\,
            I => \N__55980\
        );

    \I__13255\ : Span4Mux_s2_v
    port map (
            O => \N__55980\,
            I => \N__55977\
        );

    \I__13254\ : Odrv4
    port map (
            O => \N__55977\,
            I => pwm_out
        );

    \I__13253\ : IoInMux
    port map (
            O => \N__55974\,
            I => \N__55971\
        );

    \I__13252\ : LocalMux
    port map (
            O => \N__55971\,
            I => \N__55968\
        );

    \I__13251\ : IoSpan4Mux
    port map (
            O => \N__55968\,
            I => \N__55965\
        );

    \I__13250\ : Span4Mux_s0_v
    port map (
            O => \N__55965\,
            I => \N__55962\
        );

    \I__13249\ : Odrv4
    port map (
            O => \N__55962\,
            I => \INHA_c_0\
        );

    \I__13248\ : InMux
    port map (
            O => \N__55959\,
            I => \N__55956\
        );

    \I__13247\ : LocalMux
    port map (
            O => \N__55956\,
            I => \N__55952\
        );

    \I__13246\ : InMux
    port map (
            O => \N__55955\,
            I => \N__55949\
        );

    \I__13245\ : Span4Mux_h
    port map (
            O => \N__55952\,
            I => \N__55946\
        );

    \I__13244\ : LocalMux
    port map (
            O => \N__55949\,
            I => sweep_counter_15
        );

    \I__13243\ : Odrv4
    port map (
            O => \N__55946\,
            I => sweep_counter_15
        );

    \I__13242\ : InMux
    port map (
            O => \N__55941\,
            I => n13067
        );

    \I__13241\ : InMux
    port map (
            O => \N__55938\,
            I => \N__55934\
        );

    \I__13240\ : InMux
    port map (
            O => \N__55937\,
            I => \N__55931\
        );

    \I__13239\ : LocalMux
    port map (
            O => \N__55934\,
            I => \N__55928\
        );

    \I__13238\ : LocalMux
    port map (
            O => \N__55931\,
            I => sweep_counter_16
        );

    \I__13237\ : Odrv4
    port map (
            O => \N__55928\,
            I => sweep_counter_16
        );

    \I__13236\ : InMux
    port map (
            O => \N__55923\,
            I => \bfn_16_27_0_\
        );

    \I__13235\ : InMux
    port map (
            O => \N__55920\,
            I => n13069
        );

    \I__13234\ : SRMux
    port map (
            O => \N__55917\,
            I => \N__55913\
        );

    \I__13233\ : CEMux
    port map (
            O => \N__55916\,
            I => \N__55908\
        );

    \I__13232\ : LocalMux
    port map (
            O => \N__55913\,
            I => \N__55905\
        );

    \I__13231\ : SRMux
    port map (
            O => \N__55912\,
            I => \N__55902\
        );

    \I__13230\ : CEMux
    port map (
            O => \N__55911\,
            I => \N__55899\
        );

    \I__13229\ : LocalMux
    port map (
            O => \N__55908\,
            I => \N__55894\
        );

    \I__13228\ : Span4Mux_v
    port map (
            O => \N__55905\,
            I => \N__55891\
        );

    \I__13227\ : LocalMux
    port map (
            O => \N__55902\,
            I => \N__55888\
        );

    \I__13226\ : LocalMux
    port map (
            O => \N__55899\,
            I => \N__55885\
        );

    \I__13225\ : CEMux
    port map (
            O => \N__55898\,
            I => \N__55882\
        );

    \I__13224\ : SRMux
    port map (
            O => \N__55897\,
            I => \N__55878\
        );

    \I__13223\ : Span4Mux_h
    port map (
            O => \N__55894\,
            I => \N__55875\
        );

    \I__13222\ : Span4Mux_v
    port map (
            O => \N__55891\,
            I => \N__55872\
        );

    \I__13221\ : Span4Mux_h
    port map (
            O => \N__55888\,
            I => \N__55869\
        );

    \I__13220\ : Span4Mux_v
    port map (
            O => \N__55885\,
            I => \N__55866\
        );

    \I__13219\ : LocalMux
    port map (
            O => \N__55882\,
            I => \N__55863\
        );

    \I__13218\ : CEMux
    port map (
            O => \N__55881\,
            I => \N__55860\
        );

    \I__13217\ : LocalMux
    port map (
            O => \N__55878\,
            I => \N__55857\
        );

    \I__13216\ : Span4Mux_v
    port map (
            O => \N__55875\,
            I => \N__55850\
        );

    \I__13215\ : Span4Mux_h
    port map (
            O => \N__55872\,
            I => \N__55850\
        );

    \I__13214\ : Span4Mux_v
    port map (
            O => \N__55869\,
            I => \N__55850\
        );

    \I__13213\ : Span4Mux_h
    port map (
            O => \N__55866\,
            I => \N__55841\
        );

    \I__13212\ : Span4Mux_v
    port map (
            O => \N__55863\,
            I => \N__55841\
        );

    \I__13211\ : LocalMux
    port map (
            O => \N__55860\,
            I => \N__55841\
        );

    \I__13210\ : Span4Mux_h
    port map (
            O => \N__55857\,
            I => \N__55841\
        );

    \I__13209\ : Odrv4
    port map (
            O => \N__55850\,
            I => n5215
        );

    \I__13208\ : Odrv4
    port map (
            O => \N__55841\,
            I => n5215
        );

    \I__13207\ : InMux
    port map (
            O => \N__55836\,
            I => \N__55832\
        );

    \I__13206\ : InMux
    port map (
            O => \N__55835\,
            I => \N__55829\
        );

    \I__13205\ : LocalMux
    port map (
            O => \N__55832\,
            I => \N__55826\
        );

    \I__13204\ : LocalMux
    port map (
            O => \N__55829\,
            I => sweep_counter_8
        );

    \I__13203\ : Odrv4
    port map (
            O => \N__55826\,
            I => sweep_counter_8
        );

    \I__13202\ : InMux
    port map (
            O => \N__55821\,
            I => \N__55817\
        );

    \I__13201\ : InMux
    port map (
            O => \N__55820\,
            I => \N__55814\
        );

    \I__13200\ : LocalMux
    port map (
            O => \N__55817\,
            I => \N__55811\
        );

    \I__13199\ : LocalMux
    port map (
            O => \N__55814\,
            I => sweep_counter_14
        );

    \I__13198\ : Odrv4
    port map (
            O => \N__55811\,
            I => sweep_counter_14
        );

    \I__13197\ : InMux
    port map (
            O => \N__55806\,
            I => \N__55802\
        );

    \I__13196\ : InMux
    port map (
            O => \N__55805\,
            I => \N__55799\
        );

    \I__13195\ : LocalMux
    port map (
            O => \N__55802\,
            I => \N__55796\
        );

    \I__13194\ : LocalMux
    port map (
            O => \N__55799\,
            I => sweep_counter_13
        );

    \I__13193\ : Odrv4
    port map (
            O => \N__55796\,
            I => sweep_counter_13
        );

    \I__13192\ : InMux
    port map (
            O => \N__55791\,
            I => \N__55787\
        );

    \I__13191\ : InMux
    port map (
            O => \N__55790\,
            I => \N__55784\
        );

    \I__13190\ : LocalMux
    port map (
            O => \N__55787\,
            I => sweep_counter_17
        );

    \I__13189\ : LocalMux
    port map (
            O => \N__55784\,
            I => sweep_counter_17
        );

    \I__13188\ : CascadeMux
    port map (
            O => \N__55779\,
            I => \n6_adj_712_cascade_\
        );

    \I__13187\ : InMux
    port map (
            O => \N__55776\,
            I => \N__55772\
        );

    \I__13186\ : InMux
    port map (
            O => \N__55775\,
            I => \N__55769\
        );

    \I__13185\ : LocalMux
    port map (
            O => \N__55772\,
            I => \N__55766\
        );

    \I__13184\ : LocalMux
    port map (
            O => \N__55769\,
            I => sweep_counter_12
        );

    \I__13183\ : Odrv4
    port map (
            O => \N__55766\,
            I => sweep_counter_12
        );

    \I__13182\ : InMux
    port map (
            O => \N__55761\,
            I => \N__55757\
        );

    \I__13181\ : InMux
    port map (
            O => \N__55760\,
            I => \N__55754\
        );

    \I__13180\ : LocalMux
    port map (
            O => \N__55757\,
            I => \N__55751\
        );

    \I__13179\ : LocalMux
    port map (
            O => \N__55754\,
            I => \N__55748\
        );

    \I__13178\ : Span4Mux_h
    port map (
            O => \N__55751\,
            I => \N__55745\
        );

    \I__13177\ : Span4Mux_h
    port map (
            O => \N__55748\,
            I => \N__55742\
        );

    \I__13176\ : Span4Mux_v
    port map (
            O => \N__55745\,
            I => \N__55739\
        );

    \I__13175\ : Odrv4
    port map (
            O => \N__55742\,
            I => n13968
        );

    \I__13174\ : Odrv4
    port map (
            O => \N__55739\,
            I => n13968
        );

    \I__13173\ : InMux
    port map (
            O => \N__55734\,
            I => \N__55731\
        );

    \I__13172\ : LocalMux
    port map (
            O => \N__55731\,
            I => \GHC\
        );

    \I__13171\ : IoInMux
    port map (
            O => \N__55728\,
            I => \N__55725\
        );

    \I__13170\ : LocalMux
    port map (
            O => \N__55725\,
            I => \N__55722\
        );

    \I__13169\ : Span12Mux_s0_v
    port map (
            O => \N__55722\,
            I => \N__55719\
        );

    \I__13168\ : Odrv12
    port map (
            O => \N__55719\,
            I => \INHC_c_0\
        );

    \I__13167\ : InMux
    port map (
            O => \N__55716\,
            I => \N__55712\
        );

    \I__13166\ : InMux
    port map (
            O => \N__55715\,
            I => \N__55709\
        );

    \I__13165\ : LocalMux
    port map (
            O => \N__55712\,
            I => \N__55706\
        );

    \I__13164\ : LocalMux
    port map (
            O => \N__55709\,
            I => sweep_counter_6
        );

    \I__13163\ : Odrv4
    port map (
            O => \N__55706\,
            I => sweep_counter_6
        );

    \I__13162\ : InMux
    port map (
            O => \N__55701\,
            I => n13058
        );

    \I__13161\ : InMux
    port map (
            O => \N__55698\,
            I => \N__55695\
        );

    \I__13160\ : LocalMux
    port map (
            O => \N__55695\,
            I => \N__55691\
        );

    \I__13159\ : InMux
    port map (
            O => \N__55694\,
            I => \N__55688\
        );

    \I__13158\ : Span4Mux_h
    port map (
            O => \N__55691\,
            I => \N__55685\
        );

    \I__13157\ : LocalMux
    port map (
            O => \N__55688\,
            I => sweep_counter_7
        );

    \I__13156\ : Odrv4
    port map (
            O => \N__55685\,
            I => sweep_counter_7
        );

    \I__13155\ : InMux
    port map (
            O => \N__55680\,
            I => n13059
        );

    \I__13154\ : InMux
    port map (
            O => \N__55677\,
            I => \bfn_16_26_0_\
        );

    \I__13153\ : CascadeMux
    port map (
            O => \N__55674\,
            I => \N__55671\
        );

    \I__13152\ : InMux
    port map (
            O => \N__55671\,
            I => \N__55668\
        );

    \I__13151\ : LocalMux
    port map (
            O => \N__55668\,
            I => \N__55664\
        );

    \I__13150\ : InMux
    port map (
            O => \N__55667\,
            I => \N__55661\
        );

    \I__13149\ : Span4Mux_h
    port map (
            O => \N__55664\,
            I => \N__55658\
        );

    \I__13148\ : LocalMux
    port map (
            O => \N__55661\,
            I => sweep_counter_9
        );

    \I__13147\ : Odrv4
    port map (
            O => \N__55658\,
            I => sweep_counter_9
        );

    \I__13146\ : InMux
    port map (
            O => \N__55653\,
            I => n13061
        );

    \I__13145\ : InMux
    port map (
            O => \N__55650\,
            I => \N__55647\
        );

    \I__13144\ : LocalMux
    port map (
            O => \N__55647\,
            I => \N__55643\
        );

    \I__13143\ : InMux
    port map (
            O => \N__55646\,
            I => \N__55640\
        );

    \I__13142\ : Span4Mux_h
    port map (
            O => \N__55643\,
            I => \N__55637\
        );

    \I__13141\ : LocalMux
    port map (
            O => \N__55640\,
            I => sweep_counter_10
        );

    \I__13140\ : Odrv4
    port map (
            O => \N__55637\,
            I => sweep_counter_10
        );

    \I__13139\ : InMux
    port map (
            O => \N__55632\,
            I => n13062
        );

    \I__13138\ : InMux
    port map (
            O => \N__55629\,
            I => \N__55626\
        );

    \I__13137\ : LocalMux
    port map (
            O => \N__55626\,
            I => \N__55622\
        );

    \I__13136\ : InMux
    port map (
            O => \N__55625\,
            I => \N__55619\
        );

    \I__13135\ : Span4Mux_h
    port map (
            O => \N__55622\,
            I => \N__55616\
        );

    \I__13134\ : LocalMux
    port map (
            O => \N__55619\,
            I => sweep_counter_11
        );

    \I__13133\ : Odrv4
    port map (
            O => \N__55616\,
            I => sweep_counter_11
        );

    \I__13132\ : InMux
    port map (
            O => \N__55611\,
            I => n13063
        );

    \I__13131\ : InMux
    port map (
            O => \N__55608\,
            I => n13064
        );

    \I__13130\ : InMux
    port map (
            O => \N__55605\,
            I => n13065
        );

    \I__13129\ : InMux
    port map (
            O => \N__55602\,
            I => n13066
        );

    \I__13128\ : CascadeMux
    port map (
            O => \N__55599\,
            I => \N__55596\
        );

    \I__13127\ : InMux
    port map (
            O => \N__55596\,
            I => \N__55593\
        );

    \I__13126\ : LocalMux
    port map (
            O => \N__55593\,
            I => \N__55588\
        );

    \I__13125\ : InMux
    port map (
            O => \N__55592\,
            I => \N__55583\
        );

    \I__13124\ : InMux
    port map (
            O => \N__55591\,
            I => \N__55583\
        );

    \I__13123\ : Span4Mux_v
    port map (
            O => \N__55588\,
            I => \N__55580\
        );

    \I__13122\ : LocalMux
    port map (
            O => \N__55583\,
            I => n1027
        );

    \I__13121\ : Odrv4
    port map (
            O => \N__55580\,
            I => n1027
        );

    \I__13120\ : InMux
    port map (
            O => \N__55575\,
            I => \N__55572\
        );

    \I__13119\ : LocalMux
    port map (
            O => \N__55572\,
            I => \N__55569\
        );

    \I__13118\ : Odrv4
    port map (
            O => \N__55569\,
            I => n1094
        );

    \I__13117\ : InMux
    port map (
            O => \N__55566\,
            I => n12520
        );

    \I__13116\ : CascadeMux
    port map (
            O => \N__55563\,
            I => \N__55559\
        );

    \I__13115\ : InMux
    port map (
            O => \N__55562\,
            I => \N__55521\
        );

    \I__13114\ : InMux
    port map (
            O => \N__55559\,
            I => \N__55521\
        );

    \I__13113\ : CascadeMux
    port map (
            O => \N__55558\,
            I => \N__55518\
        );

    \I__13112\ : CascadeMux
    port map (
            O => \N__55557\,
            I => \N__55515\
        );

    \I__13111\ : CascadeMux
    port map (
            O => \N__55556\,
            I => \N__55512\
        );

    \I__13110\ : CascadeMux
    port map (
            O => \N__55555\,
            I => \N__55509\
        );

    \I__13109\ : CascadeMux
    port map (
            O => \N__55554\,
            I => \N__55506\
        );

    \I__13108\ : CascadeMux
    port map (
            O => \N__55553\,
            I => \N__55503\
        );

    \I__13107\ : CascadeMux
    port map (
            O => \N__55552\,
            I => \N__55500\
        );

    \I__13106\ : CascadeMux
    port map (
            O => \N__55551\,
            I => \N__55497\
        );

    \I__13105\ : CascadeMux
    port map (
            O => \N__55550\,
            I => \N__55487\
        );

    \I__13104\ : CascadeMux
    port map (
            O => \N__55549\,
            I => \N__55482\
        );

    \I__13103\ : CascadeMux
    port map (
            O => \N__55548\,
            I => \N__55479\
        );

    \I__13102\ : CascadeMux
    port map (
            O => \N__55547\,
            I => \N__55473\
        );

    \I__13101\ : InMux
    port map (
            O => \N__55546\,
            I => \N__55470\
        );

    \I__13100\ : InMux
    port map (
            O => \N__55545\,
            I => \N__55463\
        );

    \I__13099\ : InMux
    port map (
            O => \N__55544\,
            I => \N__55463\
        );

    \I__13098\ : InMux
    port map (
            O => \N__55543\,
            I => \N__55463\
        );

    \I__13097\ : InMux
    port map (
            O => \N__55542\,
            I => \N__55456\
        );

    \I__13096\ : InMux
    port map (
            O => \N__55541\,
            I => \N__55456\
        );

    \I__13095\ : InMux
    port map (
            O => \N__55540\,
            I => \N__55456\
        );

    \I__13094\ : CascadeMux
    port map (
            O => \N__55539\,
            I => \N__55450\
        );

    \I__13093\ : CascadeMux
    port map (
            O => \N__55538\,
            I => \N__55447\
        );

    \I__13092\ : CascadeMux
    port map (
            O => \N__55537\,
            I => \N__55441\
        );

    \I__13091\ : CascadeMux
    port map (
            O => \N__55536\,
            I => \N__55438\
        );

    \I__13090\ : CascadeMux
    port map (
            O => \N__55535\,
            I => \N__55428\
        );

    \I__13089\ : CascadeMux
    port map (
            O => \N__55534\,
            I => \N__55422\
        );

    \I__13088\ : CascadeMux
    port map (
            O => \N__55533\,
            I => \N__55415\
        );

    \I__13087\ : CascadeMux
    port map (
            O => \N__55532\,
            I => \N__55412\
        );

    \I__13086\ : CascadeMux
    port map (
            O => \N__55531\,
            I => \N__55409\
        );

    \I__13085\ : CascadeMux
    port map (
            O => \N__55530\,
            I => \N__55406\
        );

    \I__13084\ : CascadeMux
    port map (
            O => \N__55529\,
            I => \N__55403\
        );

    \I__13083\ : CascadeMux
    port map (
            O => \N__55528\,
            I => \N__55400\
        );

    \I__13082\ : CascadeMux
    port map (
            O => \N__55527\,
            I => \N__55397\
        );

    \I__13081\ : CascadeMux
    port map (
            O => \N__55526\,
            I => \N__55394\
        );

    \I__13080\ : LocalMux
    port map (
            O => \N__55521\,
            I => \N__55389\
        );

    \I__13079\ : InMux
    port map (
            O => \N__55518\,
            I => \N__55380\
        );

    \I__13078\ : InMux
    port map (
            O => \N__55515\,
            I => \N__55380\
        );

    \I__13077\ : InMux
    port map (
            O => \N__55512\,
            I => \N__55380\
        );

    \I__13076\ : InMux
    port map (
            O => \N__55509\,
            I => \N__55380\
        );

    \I__13075\ : InMux
    port map (
            O => \N__55506\,
            I => \N__55371\
        );

    \I__13074\ : InMux
    port map (
            O => \N__55503\,
            I => \N__55371\
        );

    \I__13073\ : InMux
    port map (
            O => \N__55500\,
            I => \N__55371\
        );

    \I__13072\ : InMux
    port map (
            O => \N__55497\,
            I => \N__55371\
        );

    \I__13071\ : InMux
    port map (
            O => \N__55496\,
            I => \N__55368\
        );

    \I__13070\ : InMux
    port map (
            O => \N__55495\,
            I => \N__55361\
        );

    \I__13069\ : InMux
    port map (
            O => \N__55494\,
            I => \N__55361\
        );

    \I__13068\ : InMux
    port map (
            O => \N__55493\,
            I => \N__55361\
        );

    \I__13067\ : CascadeMux
    port map (
            O => \N__55492\,
            I => \N__55358\
        );

    \I__13066\ : CascadeMux
    port map (
            O => \N__55491\,
            I => \N__55352\
        );

    \I__13065\ : CascadeMux
    port map (
            O => \N__55490\,
            I => \N__55341\
        );

    \I__13064\ : InMux
    port map (
            O => \N__55487\,
            I => \N__55333\
        );

    \I__13063\ : InMux
    port map (
            O => \N__55486\,
            I => \N__55333\
        );

    \I__13062\ : InMux
    port map (
            O => \N__55485\,
            I => \N__55333\
        );

    \I__13061\ : InMux
    port map (
            O => \N__55482\,
            I => \N__55322\
        );

    \I__13060\ : InMux
    port map (
            O => \N__55479\,
            I => \N__55322\
        );

    \I__13059\ : InMux
    port map (
            O => \N__55478\,
            I => \N__55322\
        );

    \I__13058\ : InMux
    port map (
            O => \N__55477\,
            I => \N__55322\
        );

    \I__13057\ : InMux
    port map (
            O => \N__55476\,
            I => \N__55322\
        );

    \I__13056\ : InMux
    port map (
            O => \N__55473\,
            I => \N__55319\
        );

    \I__13055\ : LocalMux
    port map (
            O => \N__55470\,
            I => \N__55312\
        );

    \I__13054\ : LocalMux
    port map (
            O => \N__55463\,
            I => \N__55312\
        );

    \I__13053\ : LocalMux
    port map (
            O => \N__55456\,
            I => \N__55312\
        );

    \I__13052\ : InMux
    port map (
            O => \N__55455\,
            I => \N__55305\
        );

    \I__13051\ : InMux
    port map (
            O => \N__55454\,
            I => \N__55305\
        );

    \I__13050\ : InMux
    port map (
            O => \N__55453\,
            I => \N__55305\
        );

    \I__13049\ : InMux
    port map (
            O => \N__55450\,
            I => \N__55294\
        );

    \I__13048\ : InMux
    port map (
            O => \N__55447\,
            I => \N__55294\
        );

    \I__13047\ : InMux
    port map (
            O => \N__55446\,
            I => \N__55294\
        );

    \I__13046\ : InMux
    port map (
            O => \N__55445\,
            I => \N__55294\
        );

    \I__13045\ : InMux
    port map (
            O => \N__55444\,
            I => \N__55294\
        );

    \I__13044\ : InMux
    port map (
            O => \N__55441\,
            I => \N__55289\
        );

    \I__13043\ : InMux
    port map (
            O => \N__55438\,
            I => \N__55289\
        );

    \I__13042\ : InMux
    port map (
            O => \N__55437\,
            I => \N__55270\
        );

    \I__13041\ : InMux
    port map (
            O => \N__55436\,
            I => \N__55270\
        );

    \I__13040\ : InMux
    port map (
            O => \N__55435\,
            I => \N__55263\
        );

    \I__13039\ : InMux
    port map (
            O => \N__55434\,
            I => \N__55263\
        );

    \I__13038\ : InMux
    port map (
            O => \N__55433\,
            I => \N__55263\
        );

    \I__13037\ : InMux
    port map (
            O => \N__55432\,
            I => \N__55252\
        );

    \I__13036\ : InMux
    port map (
            O => \N__55431\,
            I => \N__55252\
        );

    \I__13035\ : InMux
    port map (
            O => \N__55428\,
            I => \N__55252\
        );

    \I__13034\ : InMux
    port map (
            O => \N__55427\,
            I => \N__55252\
        );

    \I__13033\ : InMux
    port map (
            O => \N__55426\,
            I => \N__55252\
        );

    \I__13032\ : InMux
    port map (
            O => \N__55425\,
            I => \N__55241\
        );

    \I__13031\ : InMux
    port map (
            O => \N__55422\,
            I => \N__55241\
        );

    \I__13030\ : InMux
    port map (
            O => \N__55421\,
            I => \N__55241\
        );

    \I__13029\ : InMux
    port map (
            O => \N__55420\,
            I => \N__55241\
        );

    \I__13028\ : InMux
    port map (
            O => \N__55419\,
            I => \N__55241\
        );

    \I__13027\ : InMux
    port map (
            O => \N__55418\,
            I => \N__55237\
        );

    \I__13026\ : InMux
    port map (
            O => \N__55415\,
            I => \N__55228\
        );

    \I__13025\ : InMux
    port map (
            O => \N__55412\,
            I => \N__55228\
        );

    \I__13024\ : InMux
    port map (
            O => \N__55409\,
            I => \N__55228\
        );

    \I__13023\ : InMux
    port map (
            O => \N__55406\,
            I => \N__55228\
        );

    \I__13022\ : InMux
    port map (
            O => \N__55403\,
            I => \N__55219\
        );

    \I__13021\ : InMux
    port map (
            O => \N__55400\,
            I => \N__55219\
        );

    \I__13020\ : InMux
    port map (
            O => \N__55397\,
            I => \N__55219\
        );

    \I__13019\ : InMux
    port map (
            O => \N__55394\,
            I => \N__55219\
        );

    \I__13018\ : CascadeMux
    port map (
            O => \N__55393\,
            I => \N__55215\
        );

    \I__13017\ : CascadeMux
    port map (
            O => \N__55392\,
            I => \N__55206\
        );

    \I__13016\ : Span4Mux_v
    port map (
            O => \N__55389\,
            I => \N__55192\
        );

    \I__13015\ : LocalMux
    port map (
            O => \N__55380\,
            I => \N__55192\
        );

    \I__13014\ : LocalMux
    port map (
            O => \N__55371\,
            I => \N__55192\
        );

    \I__13013\ : LocalMux
    port map (
            O => \N__55368\,
            I => \N__55192\
        );

    \I__13012\ : LocalMux
    port map (
            O => \N__55361\,
            I => \N__55192\
        );

    \I__13011\ : InMux
    port map (
            O => \N__55358\,
            I => \N__55183\
        );

    \I__13010\ : InMux
    port map (
            O => \N__55357\,
            I => \N__55183\
        );

    \I__13009\ : InMux
    port map (
            O => \N__55356\,
            I => \N__55183\
        );

    \I__13008\ : InMux
    port map (
            O => \N__55355\,
            I => \N__55183\
        );

    \I__13007\ : InMux
    port map (
            O => \N__55352\,
            I => \N__55174\
        );

    \I__13006\ : InMux
    port map (
            O => \N__55351\,
            I => \N__55174\
        );

    \I__13005\ : InMux
    port map (
            O => \N__55350\,
            I => \N__55174\
        );

    \I__13004\ : InMux
    port map (
            O => \N__55349\,
            I => \N__55174\
        );

    \I__13003\ : InMux
    port map (
            O => \N__55348\,
            I => \N__55167\
        );

    \I__13002\ : InMux
    port map (
            O => \N__55347\,
            I => \N__55167\
        );

    \I__13001\ : InMux
    port map (
            O => \N__55346\,
            I => \N__55167\
        );

    \I__13000\ : CascadeMux
    port map (
            O => \N__55345\,
            I => \N__55161\
        );

    \I__12999\ : InMux
    port map (
            O => \N__55344\,
            I => \N__55152\
        );

    \I__12998\ : InMux
    port map (
            O => \N__55341\,
            I => \N__55152\
        );

    \I__12997\ : CascadeMux
    port map (
            O => \N__55340\,
            I => \N__55148\
        );

    \I__12996\ : LocalMux
    port map (
            O => \N__55333\,
            I => \N__55141\
        );

    \I__12995\ : LocalMux
    port map (
            O => \N__55322\,
            I => \N__55141\
        );

    \I__12994\ : LocalMux
    port map (
            O => \N__55319\,
            I => \N__55141\
        );

    \I__12993\ : Span4Mux_v
    port map (
            O => \N__55312\,
            I => \N__55132\
        );

    \I__12992\ : LocalMux
    port map (
            O => \N__55305\,
            I => \N__55132\
        );

    \I__12991\ : LocalMux
    port map (
            O => \N__55294\,
            I => \N__55132\
        );

    \I__12990\ : LocalMux
    port map (
            O => \N__55289\,
            I => \N__55132\
        );

    \I__12989\ : CascadeMux
    port map (
            O => \N__55288\,
            I => \N__55122\
        );

    \I__12988\ : InMux
    port map (
            O => \N__55287\,
            I => \N__55110\
        );

    \I__12987\ : InMux
    port map (
            O => \N__55286\,
            I => \N__55110\
        );

    \I__12986\ : InMux
    port map (
            O => \N__55285\,
            I => \N__55110\
        );

    \I__12985\ : InMux
    port map (
            O => \N__55284\,
            I => \N__55101\
        );

    \I__12984\ : InMux
    port map (
            O => \N__55283\,
            I => \N__55101\
        );

    \I__12983\ : InMux
    port map (
            O => \N__55282\,
            I => \N__55101\
        );

    \I__12982\ : InMux
    port map (
            O => \N__55281\,
            I => \N__55101\
        );

    \I__12981\ : InMux
    port map (
            O => \N__55280\,
            I => \N__55098\
        );

    \I__12980\ : CascadeMux
    port map (
            O => \N__55279\,
            I => \N__55093\
        );

    \I__12979\ : CascadeMux
    port map (
            O => \N__55278\,
            I => \N__55088\
        );

    \I__12978\ : CascadeMux
    port map (
            O => \N__55277\,
            I => \N__55073\
        );

    \I__12977\ : CascadeMux
    port map (
            O => \N__55276\,
            I => \N__55070\
        );

    \I__12976\ : CascadeMux
    port map (
            O => \N__55275\,
            I => \N__55067\
        );

    \I__12975\ : LocalMux
    port map (
            O => \N__55270\,
            I => \N__55046\
        );

    \I__12974\ : LocalMux
    port map (
            O => \N__55263\,
            I => \N__55046\
        );

    \I__12973\ : LocalMux
    port map (
            O => \N__55252\,
            I => \N__55046\
        );

    \I__12972\ : LocalMux
    port map (
            O => \N__55241\,
            I => \N__55046\
        );

    \I__12971\ : CascadeMux
    port map (
            O => \N__55240\,
            I => \N__55042\
        );

    \I__12970\ : LocalMux
    port map (
            O => \N__55237\,
            I => \N__55023\
        );

    \I__12969\ : LocalMux
    port map (
            O => \N__55228\,
            I => \N__55023\
        );

    \I__12968\ : LocalMux
    port map (
            O => \N__55219\,
            I => \N__55023\
        );

    \I__12967\ : InMux
    port map (
            O => \N__55218\,
            I => \N__55020\
        );

    \I__12966\ : InMux
    port map (
            O => \N__55215\,
            I => \N__55011\
        );

    \I__12965\ : InMux
    port map (
            O => \N__55214\,
            I => \N__55011\
        );

    \I__12964\ : InMux
    port map (
            O => \N__55213\,
            I => \N__55011\
        );

    \I__12963\ : InMux
    port map (
            O => \N__55212\,
            I => \N__55011\
        );

    \I__12962\ : InMux
    port map (
            O => \N__55211\,
            I => \N__55004\
        );

    \I__12961\ : InMux
    port map (
            O => \N__55210\,
            I => \N__55004\
        );

    \I__12960\ : InMux
    port map (
            O => \N__55209\,
            I => \N__55004\
        );

    \I__12959\ : InMux
    port map (
            O => \N__55206\,
            I => \N__54995\
        );

    \I__12958\ : InMux
    port map (
            O => \N__55205\,
            I => \N__54995\
        );

    \I__12957\ : InMux
    port map (
            O => \N__55204\,
            I => \N__54995\
        );

    \I__12956\ : InMux
    port map (
            O => \N__55203\,
            I => \N__54995\
        );

    \I__12955\ : Span4Mux_v
    port map (
            O => \N__55192\,
            I => \N__54988\
        );

    \I__12954\ : LocalMux
    port map (
            O => \N__55183\,
            I => \N__54988\
        );

    \I__12953\ : LocalMux
    port map (
            O => \N__55174\,
            I => \N__54988\
        );

    \I__12952\ : LocalMux
    port map (
            O => \N__55167\,
            I => \N__54985\
        );

    \I__12951\ : InMux
    port map (
            O => \N__55166\,
            I => \N__54974\
        );

    \I__12950\ : InMux
    port map (
            O => \N__55165\,
            I => \N__54974\
        );

    \I__12949\ : InMux
    port map (
            O => \N__55164\,
            I => \N__54974\
        );

    \I__12948\ : InMux
    port map (
            O => \N__55161\,
            I => \N__54974\
        );

    \I__12947\ : InMux
    port map (
            O => \N__55160\,
            I => \N__54974\
        );

    \I__12946\ : InMux
    port map (
            O => \N__55159\,
            I => \N__54967\
        );

    \I__12945\ : InMux
    port map (
            O => \N__55158\,
            I => \N__54967\
        );

    \I__12944\ : InMux
    port map (
            O => \N__55157\,
            I => \N__54967\
        );

    \I__12943\ : LocalMux
    port map (
            O => \N__55152\,
            I => \N__54964\
        );

    \I__12942\ : InMux
    port map (
            O => \N__55151\,
            I => \N__54959\
        );

    \I__12941\ : InMux
    port map (
            O => \N__55148\,
            I => \N__54959\
        );

    \I__12940\ : Span4Mux_s3_h
    port map (
            O => \N__55141\,
            I => \N__54947\
        );

    \I__12939\ : Span4Mux_v
    port map (
            O => \N__55132\,
            I => \N__54947\
        );

    \I__12938\ : InMux
    port map (
            O => \N__55131\,
            I => \N__54944\
        );

    \I__12937\ : InMux
    port map (
            O => \N__55130\,
            I => \N__54937\
        );

    \I__12936\ : InMux
    port map (
            O => \N__55129\,
            I => \N__54937\
        );

    \I__12935\ : InMux
    port map (
            O => \N__55128\,
            I => \N__54937\
        );

    \I__12934\ : InMux
    port map (
            O => \N__55127\,
            I => \N__54932\
        );

    \I__12933\ : InMux
    port map (
            O => \N__55126\,
            I => \N__54932\
        );

    \I__12932\ : InMux
    port map (
            O => \N__55125\,
            I => \N__54925\
        );

    \I__12931\ : InMux
    port map (
            O => \N__55122\,
            I => \N__54925\
        );

    \I__12930\ : InMux
    port map (
            O => \N__55121\,
            I => \N__54925\
        );

    \I__12929\ : InMux
    port map (
            O => \N__55120\,
            I => \N__54922\
        );

    \I__12928\ : InMux
    port map (
            O => \N__55119\,
            I => \N__54915\
        );

    \I__12927\ : InMux
    port map (
            O => \N__55118\,
            I => \N__54915\
        );

    \I__12926\ : InMux
    port map (
            O => \N__55117\,
            I => \N__54915\
        );

    \I__12925\ : LocalMux
    port map (
            O => \N__55110\,
            I => \N__54908\
        );

    \I__12924\ : LocalMux
    port map (
            O => \N__55101\,
            I => \N__54908\
        );

    \I__12923\ : LocalMux
    port map (
            O => \N__55098\,
            I => \N__54908\
        );

    \I__12922\ : InMux
    port map (
            O => \N__55097\,
            I => \N__54903\
        );

    \I__12921\ : InMux
    port map (
            O => \N__55096\,
            I => \N__54903\
        );

    \I__12920\ : InMux
    port map (
            O => \N__55093\,
            I => \N__54894\
        );

    \I__12919\ : InMux
    port map (
            O => \N__55092\,
            I => \N__54894\
        );

    \I__12918\ : InMux
    port map (
            O => \N__55091\,
            I => \N__54894\
        );

    \I__12917\ : InMux
    port map (
            O => \N__55088\,
            I => \N__54894\
        );

    \I__12916\ : InMux
    port map (
            O => \N__55087\,
            I => \N__54887\
        );

    \I__12915\ : InMux
    port map (
            O => \N__55086\,
            I => \N__54884\
        );

    \I__12914\ : CascadeMux
    port map (
            O => \N__55085\,
            I => \N__54857\
        );

    \I__12913\ : CascadeMux
    port map (
            O => \N__55084\,
            I => \N__54854\
        );

    \I__12912\ : CascadeMux
    port map (
            O => \N__55083\,
            I => \N__54851\
        );

    \I__12911\ : CascadeMux
    port map (
            O => \N__55082\,
            I => \N__54848\
        );

    \I__12910\ : CascadeMux
    port map (
            O => \N__55081\,
            I => \N__54845\
        );

    \I__12909\ : CascadeMux
    port map (
            O => \N__55080\,
            I => \N__54842\
        );

    \I__12908\ : CascadeMux
    port map (
            O => \N__55079\,
            I => \N__54839\
        );

    \I__12907\ : CascadeMux
    port map (
            O => \N__55078\,
            I => \N__54836\
        );

    \I__12906\ : CascadeMux
    port map (
            O => \N__55077\,
            I => \N__54833\
        );

    \I__12905\ : CascadeMux
    port map (
            O => \N__55076\,
            I => \N__54830\
        );

    \I__12904\ : InMux
    port map (
            O => \N__55073\,
            I => \N__54823\
        );

    \I__12903\ : InMux
    port map (
            O => \N__55070\,
            I => \N__54823\
        );

    \I__12902\ : InMux
    port map (
            O => \N__55067\,
            I => \N__54823\
        );

    \I__12901\ : CascadeMux
    port map (
            O => \N__55066\,
            I => \N__54820\
        );

    \I__12900\ : CascadeMux
    port map (
            O => \N__55065\,
            I => \N__54817\
        );

    \I__12899\ : CascadeMux
    port map (
            O => \N__55064\,
            I => \N__54814\
        );

    \I__12898\ : CascadeMux
    port map (
            O => \N__55063\,
            I => \N__54810\
        );

    \I__12897\ : CascadeMux
    port map (
            O => \N__55062\,
            I => \N__54807\
        );

    \I__12896\ : CascadeMux
    port map (
            O => \N__55061\,
            I => \N__54804\
        );

    \I__12895\ : CascadeMux
    port map (
            O => \N__55060\,
            I => \N__54801\
        );

    \I__12894\ : CascadeMux
    port map (
            O => \N__55059\,
            I => \N__54798\
        );

    \I__12893\ : CascadeMux
    port map (
            O => \N__55058\,
            I => \N__54795\
        );

    \I__12892\ : CascadeMux
    port map (
            O => \N__55057\,
            I => \N__54789\
        );

    \I__12891\ : CascadeMux
    port map (
            O => \N__55056\,
            I => \N__54780\
        );

    \I__12890\ : CascadeMux
    port map (
            O => \N__55055\,
            I => \N__54777\
        );

    \I__12889\ : Span4Mux_v
    port map (
            O => \N__55046\,
            I => \N__54773\
        );

    \I__12888\ : InMux
    port map (
            O => \N__55045\,
            I => \N__54770\
        );

    \I__12887\ : InMux
    port map (
            O => \N__55042\,
            I => \N__54767\
        );

    \I__12886\ : CascadeMux
    port map (
            O => \N__55041\,
            I => \N__54764\
        );

    \I__12885\ : CascadeMux
    port map (
            O => \N__55040\,
            I => \N__54759\
        );

    \I__12884\ : CascadeMux
    port map (
            O => \N__55039\,
            I => \N__54753\
        );

    \I__12883\ : CascadeMux
    port map (
            O => \N__55038\,
            I => \N__54750\
        );

    \I__12882\ : CascadeMux
    port map (
            O => \N__55037\,
            I => \N__54747\
        );

    \I__12881\ : CascadeMux
    port map (
            O => \N__55036\,
            I => \N__54740\
        );

    \I__12880\ : CascadeMux
    port map (
            O => \N__55035\,
            I => \N__54737\
        );

    \I__12879\ : CascadeMux
    port map (
            O => \N__55034\,
            I => \N__54733\
        );

    \I__12878\ : InMux
    port map (
            O => \N__55033\,
            I => \N__54714\
        );

    \I__12877\ : InMux
    port map (
            O => \N__55032\,
            I => \N__54714\
        );

    \I__12876\ : InMux
    port map (
            O => \N__55031\,
            I => \N__54714\
        );

    \I__12875\ : CascadeMux
    port map (
            O => \N__55030\,
            I => \N__54710\
        );

    \I__12874\ : Span4Mux_v
    port map (
            O => \N__55023\,
            I => \N__54702\
        );

    \I__12873\ : LocalMux
    port map (
            O => \N__55020\,
            I => \N__54695\
        );

    \I__12872\ : LocalMux
    port map (
            O => \N__55011\,
            I => \N__54695\
        );

    \I__12871\ : LocalMux
    port map (
            O => \N__55004\,
            I => \N__54690\
        );

    \I__12870\ : LocalMux
    port map (
            O => \N__54995\,
            I => \N__54690\
        );

    \I__12869\ : Span4Mux_h
    port map (
            O => \N__54988\,
            I => \N__54677\
        );

    \I__12868\ : Span4Mux_v
    port map (
            O => \N__54985\,
            I => \N__54677\
        );

    \I__12867\ : LocalMux
    port map (
            O => \N__54974\,
            I => \N__54677\
        );

    \I__12866\ : LocalMux
    port map (
            O => \N__54967\,
            I => \N__54677\
        );

    \I__12865\ : Span4Mux_v
    port map (
            O => \N__54964\,
            I => \N__54677\
        );

    \I__12864\ : LocalMux
    port map (
            O => \N__54959\,
            I => \N__54677\
        );

    \I__12863\ : InMux
    port map (
            O => \N__54958\,
            I => \N__54668\
        );

    \I__12862\ : InMux
    port map (
            O => \N__54957\,
            I => \N__54668\
        );

    \I__12861\ : InMux
    port map (
            O => \N__54956\,
            I => \N__54668\
        );

    \I__12860\ : InMux
    port map (
            O => \N__54955\,
            I => \N__54668\
        );

    \I__12859\ : InMux
    port map (
            O => \N__54954\,
            I => \N__54663\
        );

    \I__12858\ : InMux
    port map (
            O => \N__54953\,
            I => \N__54663\
        );

    \I__12857\ : CascadeMux
    port map (
            O => \N__54952\,
            I => \N__54658\
        );

    \I__12856\ : Span4Mux_h
    port map (
            O => \N__54947\,
            I => \N__54640\
        );

    \I__12855\ : LocalMux
    port map (
            O => \N__54944\,
            I => \N__54627\
        );

    \I__12854\ : LocalMux
    port map (
            O => \N__54937\,
            I => \N__54627\
        );

    \I__12853\ : LocalMux
    port map (
            O => \N__54932\,
            I => \N__54627\
        );

    \I__12852\ : LocalMux
    port map (
            O => \N__54925\,
            I => \N__54627\
        );

    \I__12851\ : LocalMux
    port map (
            O => \N__54922\,
            I => \N__54627\
        );

    \I__12850\ : LocalMux
    port map (
            O => \N__54915\,
            I => \N__54627\
        );

    \I__12849\ : Span4Mux_v
    port map (
            O => \N__54908\,
            I => \N__54624\
        );

    \I__12848\ : LocalMux
    port map (
            O => \N__54903\,
            I => \N__54621\
        );

    \I__12847\ : LocalMux
    port map (
            O => \N__54894\,
            I => \N__54618\
        );

    \I__12846\ : InMux
    port map (
            O => \N__54893\,
            I => \N__54615\
        );

    \I__12845\ : InMux
    port map (
            O => \N__54892\,
            I => \N__54608\
        );

    \I__12844\ : InMux
    port map (
            O => \N__54891\,
            I => \N__54608\
        );

    \I__12843\ : InMux
    port map (
            O => \N__54890\,
            I => \N__54608\
        );

    \I__12842\ : LocalMux
    port map (
            O => \N__54887\,
            I => \N__54603\
        );

    \I__12841\ : LocalMux
    port map (
            O => \N__54884\,
            I => \N__54603\
        );

    \I__12840\ : InMux
    port map (
            O => \N__54883\,
            I => \N__54596\
        );

    \I__12839\ : InMux
    port map (
            O => \N__54882\,
            I => \N__54596\
        );

    \I__12838\ : InMux
    port map (
            O => \N__54881\,
            I => \N__54596\
        );

    \I__12837\ : CascadeMux
    port map (
            O => \N__54880\,
            I => \N__54593\
        );

    \I__12836\ : CascadeMux
    port map (
            O => \N__54879\,
            I => \N__54583\
        );

    \I__12835\ : CascadeMux
    port map (
            O => \N__54878\,
            I => \N__54569\
        );

    \I__12834\ : CascadeMux
    port map (
            O => \N__54877\,
            I => \N__54566\
        );

    \I__12833\ : CascadeMux
    port map (
            O => \N__54876\,
            I => \N__54561\
        );

    \I__12832\ : CascadeMux
    port map (
            O => \N__54875\,
            I => \N__54558\
        );

    \I__12831\ : CascadeMux
    port map (
            O => \N__54874\,
            I => \N__54553\
        );

    \I__12830\ : CascadeMux
    port map (
            O => \N__54873\,
            I => \N__54550\
        );

    \I__12829\ : CascadeMux
    port map (
            O => \N__54872\,
            I => \N__54547\
        );

    \I__12828\ : CascadeMux
    port map (
            O => \N__54871\,
            I => \N__54544\
        );

    \I__12827\ : CascadeMux
    port map (
            O => \N__54870\,
            I => \N__54541\
        );

    \I__12826\ : CascadeMux
    port map (
            O => \N__54869\,
            I => \N__54538\
        );

    \I__12825\ : CascadeMux
    port map (
            O => \N__54868\,
            I => \N__54535\
        );

    \I__12824\ : CascadeMux
    port map (
            O => \N__54867\,
            I => \N__54531\
        );

    \I__12823\ : CascadeMux
    port map (
            O => \N__54866\,
            I => \N__54528\
        );

    \I__12822\ : CascadeMux
    port map (
            O => \N__54865\,
            I => \N__54525\
        );

    \I__12821\ : CascadeMux
    port map (
            O => \N__54864\,
            I => \N__54522\
        );

    \I__12820\ : CascadeMux
    port map (
            O => \N__54863\,
            I => \N__54519\
        );

    \I__12819\ : CascadeMux
    port map (
            O => \N__54862\,
            I => \N__54516\
        );

    \I__12818\ : CascadeMux
    port map (
            O => \N__54861\,
            I => \N__54512\
        );

    \I__12817\ : CascadeMux
    port map (
            O => \N__54860\,
            I => \N__54509\
        );

    \I__12816\ : InMux
    port map (
            O => \N__54857\,
            I => \N__54499\
        );

    \I__12815\ : InMux
    port map (
            O => \N__54854\,
            I => \N__54499\
        );

    \I__12814\ : InMux
    port map (
            O => \N__54851\,
            I => \N__54499\
        );

    \I__12813\ : InMux
    port map (
            O => \N__54848\,
            I => \N__54492\
        );

    \I__12812\ : InMux
    port map (
            O => \N__54845\,
            I => \N__54492\
        );

    \I__12811\ : InMux
    port map (
            O => \N__54842\,
            I => \N__54492\
        );

    \I__12810\ : InMux
    port map (
            O => \N__54839\,
            I => \N__54483\
        );

    \I__12809\ : InMux
    port map (
            O => \N__54836\,
            I => \N__54483\
        );

    \I__12808\ : InMux
    port map (
            O => \N__54833\,
            I => \N__54483\
        );

    \I__12807\ : InMux
    port map (
            O => \N__54830\,
            I => \N__54483\
        );

    \I__12806\ : LocalMux
    port map (
            O => \N__54823\,
            I => \N__54480\
        );

    \I__12805\ : InMux
    port map (
            O => \N__54820\,
            I => \N__54477\
        );

    \I__12804\ : InMux
    port map (
            O => \N__54817\,
            I => \N__54466\
        );

    \I__12803\ : InMux
    port map (
            O => \N__54814\,
            I => \N__54466\
        );

    \I__12802\ : InMux
    port map (
            O => \N__54813\,
            I => \N__54466\
        );

    \I__12801\ : InMux
    port map (
            O => \N__54810\,
            I => \N__54466\
        );

    \I__12800\ : InMux
    port map (
            O => \N__54807\,
            I => \N__54466\
        );

    \I__12799\ : InMux
    port map (
            O => \N__54804\,
            I => \N__54457\
        );

    \I__12798\ : InMux
    port map (
            O => \N__54801\,
            I => \N__54457\
        );

    \I__12797\ : InMux
    port map (
            O => \N__54798\,
            I => \N__54457\
        );

    \I__12796\ : InMux
    port map (
            O => \N__54795\,
            I => \N__54457\
        );

    \I__12795\ : InMux
    port map (
            O => \N__54794\,
            I => \N__54452\
        );

    \I__12794\ : InMux
    port map (
            O => \N__54793\,
            I => \N__54452\
        );

    \I__12793\ : InMux
    port map (
            O => \N__54792\,
            I => \N__54447\
        );

    \I__12792\ : InMux
    port map (
            O => \N__54789\,
            I => \N__54447\
        );

    \I__12791\ : InMux
    port map (
            O => \N__54788\,
            I => \N__54438\
        );

    \I__12790\ : InMux
    port map (
            O => \N__54787\,
            I => \N__54438\
        );

    \I__12789\ : InMux
    port map (
            O => \N__54786\,
            I => \N__54431\
        );

    \I__12788\ : InMux
    port map (
            O => \N__54785\,
            I => \N__54431\
        );

    \I__12787\ : InMux
    port map (
            O => \N__54784\,
            I => \N__54431\
        );

    \I__12786\ : InMux
    port map (
            O => \N__54783\,
            I => \N__54424\
        );

    \I__12785\ : InMux
    port map (
            O => \N__54780\,
            I => \N__54424\
        );

    \I__12784\ : InMux
    port map (
            O => \N__54777\,
            I => \N__54424\
        );

    \I__12783\ : CascadeMux
    port map (
            O => \N__54776\,
            I => \N__54418\
        );

    \I__12782\ : Span4Mux_h
    port map (
            O => \N__54773\,
            I => \N__54407\
        );

    \I__12781\ : LocalMux
    port map (
            O => \N__54770\,
            I => \N__54407\
        );

    \I__12780\ : LocalMux
    port map (
            O => \N__54767\,
            I => \N__54407\
        );

    \I__12779\ : InMux
    port map (
            O => \N__54764\,
            I => \N__54402\
        );

    \I__12778\ : InMux
    port map (
            O => \N__54763\,
            I => \N__54402\
        );

    \I__12777\ : InMux
    port map (
            O => \N__54762\,
            I => \N__54391\
        );

    \I__12776\ : InMux
    port map (
            O => \N__54759\,
            I => \N__54391\
        );

    \I__12775\ : InMux
    port map (
            O => \N__54758\,
            I => \N__54391\
        );

    \I__12774\ : InMux
    port map (
            O => \N__54757\,
            I => \N__54391\
        );

    \I__12773\ : InMux
    port map (
            O => \N__54756\,
            I => \N__54391\
        );

    \I__12772\ : InMux
    port map (
            O => \N__54753\,
            I => \N__54382\
        );

    \I__12771\ : InMux
    port map (
            O => \N__54750\,
            I => \N__54382\
        );

    \I__12770\ : InMux
    port map (
            O => \N__54747\,
            I => \N__54382\
        );

    \I__12769\ : InMux
    port map (
            O => \N__54746\,
            I => \N__54382\
        );

    \I__12768\ : CascadeMux
    port map (
            O => \N__54745\,
            I => \N__54376\
        );

    \I__12767\ : CascadeMux
    port map (
            O => \N__54744\,
            I => \N__54370\
        );

    \I__12766\ : InMux
    port map (
            O => \N__54743\,
            I => \N__54364\
        );

    \I__12765\ : InMux
    port map (
            O => \N__54740\,
            I => \N__54357\
        );

    \I__12764\ : InMux
    port map (
            O => \N__54737\,
            I => \N__54357\
        );

    \I__12763\ : InMux
    port map (
            O => \N__54736\,
            I => \N__54357\
        );

    \I__12762\ : InMux
    port map (
            O => \N__54733\,
            I => \N__54352\
        );

    \I__12761\ : InMux
    port map (
            O => \N__54732\,
            I => \N__54352\
        );

    \I__12760\ : CascadeMux
    port map (
            O => \N__54731\,
            I => \N__54348\
        );

    \I__12759\ : CascadeMux
    port map (
            O => \N__54730\,
            I => \N__54342\
        );

    \I__12758\ : CascadeMux
    port map (
            O => \N__54729\,
            I => \N__54339\
        );

    \I__12757\ : CascadeMux
    port map (
            O => \N__54728\,
            I => \N__54336\
        );

    \I__12756\ : CascadeMux
    port map (
            O => \N__54727\,
            I => \N__54333\
        );

    \I__12755\ : CascadeMux
    port map (
            O => \N__54726\,
            I => \N__54330\
        );

    \I__12754\ : CascadeMux
    port map (
            O => \N__54725\,
            I => \N__54321\
        );

    \I__12753\ : CascadeMux
    port map (
            O => \N__54724\,
            I => \N__54318\
        );

    \I__12752\ : CascadeMux
    port map (
            O => \N__54723\,
            I => \N__54315\
        );

    \I__12751\ : CascadeMux
    port map (
            O => \N__54722\,
            I => \N__54312\
        );

    \I__12750\ : CascadeMux
    port map (
            O => \N__54721\,
            I => \N__54309\
        );

    \I__12749\ : LocalMux
    port map (
            O => \N__54714\,
            I => \N__54306\
        );

    \I__12748\ : InMux
    port map (
            O => \N__54713\,
            I => \N__54297\
        );

    \I__12747\ : InMux
    port map (
            O => \N__54710\,
            I => \N__54297\
        );

    \I__12746\ : InMux
    port map (
            O => \N__54709\,
            I => \N__54297\
        );

    \I__12745\ : InMux
    port map (
            O => \N__54708\,
            I => \N__54297\
        );

    \I__12744\ : CascadeMux
    port map (
            O => \N__54707\,
            I => \N__54294\
        );

    \I__12743\ : CascadeMux
    port map (
            O => \N__54706\,
            I => \N__54289\
        );

    \I__12742\ : CascadeMux
    port map (
            O => \N__54705\,
            I => \N__54284\
        );

    \I__12741\ : Span4Mux_h
    port map (
            O => \N__54702\,
            I => \N__54280\
        );

    \I__12740\ : InMux
    port map (
            O => \N__54701\,
            I => \N__54275\
        );

    \I__12739\ : InMux
    port map (
            O => \N__54700\,
            I => \N__54275\
        );

    \I__12738\ : Span4Mux_v
    port map (
            O => \N__54695\,
            I => \N__54270\
        );

    \I__12737\ : Span4Mux_v
    port map (
            O => \N__54690\,
            I => \N__54270\
        );

    \I__12736\ : Span4Mux_h
    port map (
            O => \N__54677\,
            I => \N__54263\
        );

    \I__12735\ : LocalMux
    port map (
            O => \N__54668\,
            I => \N__54263\
        );

    \I__12734\ : LocalMux
    port map (
            O => \N__54663\,
            I => \N__54263\
        );

    \I__12733\ : InMux
    port map (
            O => \N__54662\,
            I => \N__54258\
        );

    \I__12732\ : InMux
    port map (
            O => \N__54661\,
            I => \N__54258\
        );

    \I__12731\ : InMux
    port map (
            O => \N__54658\,
            I => \N__54253\
        );

    \I__12730\ : InMux
    port map (
            O => \N__54657\,
            I => \N__54253\
        );

    \I__12729\ : CascadeMux
    port map (
            O => \N__54656\,
            I => \N__54249\
        );

    \I__12728\ : CascadeMux
    port map (
            O => \N__54655\,
            I => \N__54237\
        );

    \I__12727\ : CascadeMux
    port map (
            O => \N__54654\,
            I => \N__54233\
        );

    \I__12726\ : InMux
    port map (
            O => \N__54653\,
            I => \N__54230\
        );

    \I__12725\ : InMux
    port map (
            O => \N__54652\,
            I => \N__54223\
        );

    \I__12724\ : InMux
    port map (
            O => \N__54651\,
            I => \N__54223\
        );

    \I__12723\ : InMux
    port map (
            O => \N__54650\,
            I => \N__54223\
        );

    \I__12722\ : InMux
    port map (
            O => \N__54649\,
            I => \N__54218\
        );

    \I__12721\ : InMux
    port map (
            O => \N__54648\,
            I => \N__54218\
        );

    \I__12720\ : InMux
    port map (
            O => \N__54647\,
            I => \N__54215\
        );

    \I__12719\ : InMux
    port map (
            O => \N__54646\,
            I => \N__54212\
        );

    \I__12718\ : InMux
    port map (
            O => \N__54645\,
            I => \N__54205\
        );

    \I__12717\ : InMux
    port map (
            O => \N__54644\,
            I => \N__54205\
        );

    \I__12716\ : InMux
    port map (
            O => \N__54643\,
            I => \N__54205\
        );

    \I__12715\ : Span4Mux_h
    port map (
            O => \N__54640\,
            I => \N__54186\
        );

    \I__12714\ : Span4Mux_v
    port map (
            O => \N__54627\,
            I => \N__54186\
        );

    \I__12713\ : Span4Mux_v
    port map (
            O => \N__54624\,
            I => \N__54186\
        );

    \I__12712\ : Span4Mux_h
    port map (
            O => \N__54621\,
            I => \N__54186\
        );

    \I__12711\ : Span4Mux_h
    port map (
            O => \N__54618\,
            I => \N__54186\
        );

    \I__12710\ : LocalMux
    port map (
            O => \N__54615\,
            I => \N__54186\
        );

    \I__12709\ : LocalMux
    port map (
            O => \N__54608\,
            I => \N__54186\
        );

    \I__12708\ : Span4Mux_v
    port map (
            O => \N__54603\,
            I => \N__54186\
        );

    \I__12707\ : LocalMux
    port map (
            O => \N__54596\,
            I => \N__54186\
        );

    \I__12706\ : InMux
    port map (
            O => \N__54593\,
            I => \N__54177\
        );

    \I__12705\ : InMux
    port map (
            O => \N__54592\,
            I => \N__54177\
        );

    \I__12704\ : InMux
    port map (
            O => \N__54591\,
            I => \N__54177\
        );

    \I__12703\ : InMux
    port map (
            O => \N__54590\,
            I => \N__54177\
        );

    \I__12702\ : InMux
    port map (
            O => \N__54589\,
            I => \N__54168\
        );

    \I__12701\ : InMux
    port map (
            O => \N__54588\,
            I => \N__54168\
        );

    \I__12700\ : InMux
    port map (
            O => \N__54587\,
            I => \N__54168\
        );

    \I__12699\ : InMux
    port map (
            O => \N__54586\,
            I => \N__54168\
        );

    \I__12698\ : InMux
    port map (
            O => \N__54583\,
            I => \N__54163\
        );

    \I__12697\ : InMux
    port map (
            O => \N__54582\,
            I => \N__54163\
        );

    \I__12696\ : InMux
    port map (
            O => \N__54581\,
            I => \N__54154\
        );

    \I__12695\ : InMux
    port map (
            O => \N__54580\,
            I => \N__54154\
        );

    \I__12694\ : InMux
    port map (
            O => \N__54579\,
            I => \N__54154\
        );

    \I__12693\ : InMux
    port map (
            O => \N__54578\,
            I => \N__54154\
        );

    \I__12692\ : InMux
    port map (
            O => \N__54577\,
            I => \N__54145\
        );

    \I__12691\ : InMux
    port map (
            O => \N__54576\,
            I => \N__54145\
        );

    \I__12690\ : InMux
    port map (
            O => \N__54575\,
            I => \N__54145\
        );

    \I__12689\ : InMux
    port map (
            O => \N__54574\,
            I => \N__54145\
        );

    \I__12688\ : InMux
    port map (
            O => \N__54573\,
            I => \N__54140\
        );

    \I__12687\ : InMux
    port map (
            O => \N__54572\,
            I => \N__54140\
        );

    \I__12686\ : InMux
    port map (
            O => \N__54569\,
            I => \N__54131\
        );

    \I__12685\ : InMux
    port map (
            O => \N__54566\,
            I => \N__54131\
        );

    \I__12684\ : InMux
    port map (
            O => \N__54565\,
            I => \N__54131\
        );

    \I__12683\ : InMux
    port map (
            O => \N__54564\,
            I => \N__54131\
        );

    \I__12682\ : InMux
    port map (
            O => \N__54561\,
            I => \N__54122\
        );

    \I__12681\ : InMux
    port map (
            O => \N__54558\,
            I => \N__54122\
        );

    \I__12680\ : InMux
    port map (
            O => \N__54557\,
            I => \N__54122\
        );

    \I__12679\ : InMux
    port map (
            O => \N__54556\,
            I => \N__54122\
        );

    \I__12678\ : InMux
    port map (
            O => \N__54553\,
            I => \N__54113\
        );

    \I__12677\ : InMux
    port map (
            O => \N__54550\,
            I => \N__54113\
        );

    \I__12676\ : InMux
    port map (
            O => \N__54547\,
            I => \N__54113\
        );

    \I__12675\ : InMux
    port map (
            O => \N__54544\,
            I => \N__54113\
        );

    \I__12674\ : InMux
    port map (
            O => \N__54541\,
            I => \N__54106\
        );

    \I__12673\ : InMux
    port map (
            O => \N__54538\,
            I => \N__54106\
        );

    \I__12672\ : InMux
    port map (
            O => \N__54535\,
            I => \N__54106\
        );

    \I__12671\ : InMux
    port map (
            O => \N__54534\,
            I => \N__54095\
        );

    \I__12670\ : InMux
    port map (
            O => \N__54531\,
            I => \N__54095\
        );

    \I__12669\ : InMux
    port map (
            O => \N__54528\,
            I => \N__54095\
        );

    \I__12668\ : InMux
    port map (
            O => \N__54525\,
            I => \N__54095\
        );

    \I__12667\ : InMux
    port map (
            O => \N__54522\,
            I => \N__54095\
        );

    \I__12666\ : InMux
    port map (
            O => \N__54519\,
            I => \N__54090\
        );

    \I__12665\ : InMux
    port map (
            O => \N__54516\,
            I => \N__54090\
        );

    \I__12664\ : InMux
    port map (
            O => \N__54515\,
            I => \N__54083\
        );

    \I__12663\ : InMux
    port map (
            O => \N__54512\,
            I => \N__54083\
        );

    \I__12662\ : InMux
    port map (
            O => \N__54509\,
            I => \N__54083\
        );

    \I__12661\ : InMux
    port map (
            O => \N__54508\,
            I => \N__54076\
        );

    \I__12660\ : InMux
    port map (
            O => \N__54507\,
            I => \N__54076\
        );

    \I__12659\ : InMux
    port map (
            O => \N__54506\,
            I => \N__54076\
        );

    \I__12658\ : LocalMux
    port map (
            O => \N__54499\,
            I => \N__54067\
        );

    \I__12657\ : LocalMux
    port map (
            O => \N__54492\,
            I => \N__54067\
        );

    \I__12656\ : LocalMux
    port map (
            O => \N__54483\,
            I => \N__54067\
        );

    \I__12655\ : Span4Mux_s2_h
    port map (
            O => \N__54480\,
            I => \N__54058\
        );

    \I__12654\ : LocalMux
    port map (
            O => \N__54477\,
            I => \N__54058\
        );

    \I__12653\ : LocalMux
    port map (
            O => \N__54466\,
            I => \N__54058\
        );

    \I__12652\ : LocalMux
    port map (
            O => \N__54457\,
            I => \N__54058\
        );

    \I__12651\ : LocalMux
    port map (
            O => \N__54452\,
            I => \N__54053\
        );

    \I__12650\ : LocalMux
    port map (
            O => \N__54447\,
            I => \N__54053\
        );

    \I__12649\ : InMux
    port map (
            O => \N__54446\,
            I => \N__54050\
        );

    \I__12648\ : InMux
    port map (
            O => \N__54445\,
            I => \N__54043\
        );

    \I__12647\ : InMux
    port map (
            O => \N__54444\,
            I => \N__54043\
        );

    \I__12646\ : InMux
    port map (
            O => \N__54443\,
            I => \N__54043\
        );

    \I__12645\ : LocalMux
    port map (
            O => \N__54438\,
            I => \N__54036\
        );

    \I__12644\ : LocalMux
    port map (
            O => \N__54431\,
            I => \N__54036\
        );

    \I__12643\ : LocalMux
    port map (
            O => \N__54424\,
            I => \N__54036\
        );

    \I__12642\ : InMux
    port map (
            O => \N__54423\,
            I => \N__54025\
        );

    \I__12641\ : InMux
    port map (
            O => \N__54422\,
            I => \N__54025\
        );

    \I__12640\ : InMux
    port map (
            O => \N__54421\,
            I => \N__54025\
        );

    \I__12639\ : InMux
    port map (
            O => \N__54418\,
            I => \N__54025\
        );

    \I__12638\ : InMux
    port map (
            O => \N__54417\,
            I => \N__54025\
        );

    \I__12637\ : CascadeMux
    port map (
            O => \N__54416\,
            I => \N__54017\
        );

    \I__12636\ : CascadeMux
    port map (
            O => \N__54415\,
            I => \N__54014\
        );

    \I__12635\ : CascadeMux
    port map (
            O => \N__54414\,
            I => \N__54011\
        );

    \I__12634\ : Span4Mux_v
    port map (
            O => \N__54407\,
            I => \N__54001\
        );

    \I__12633\ : LocalMux
    port map (
            O => \N__54402\,
            I => \N__54001\
        );

    \I__12632\ : LocalMux
    port map (
            O => \N__54391\,
            I => \N__54001\
        );

    \I__12631\ : LocalMux
    port map (
            O => \N__54382\,
            I => \N__54001\
        );

    \I__12630\ : InMux
    port map (
            O => \N__54381\,
            I => \N__53994\
        );

    \I__12629\ : InMux
    port map (
            O => \N__54380\,
            I => \N__53994\
        );

    \I__12628\ : InMux
    port map (
            O => \N__54379\,
            I => \N__53994\
        );

    \I__12627\ : InMux
    port map (
            O => \N__54376\,
            I => \N__53983\
        );

    \I__12626\ : InMux
    port map (
            O => \N__54375\,
            I => \N__53983\
        );

    \I__12625\ : InMux
    port map (
            O => \N__54374\,
            I => \N__53983\
        );

    \I__12624\ : InMux
    port map (
            O => \N__54373\,
            I => \N__53983\
        );

    \I__12623\ : InMux
    port map (
            O => \N__54370\,
            I => \N__53983\
        );

    \I__12622\ : CascadeMux
    port map (
            O => \N__54369\,
            I => \N__53979\
        );

    \I__12621\ : CascadeMux
    port map (
            O => \N__54368\,
            I => \N__53972\
        );

    \I__12620\ : CascadeMux
    port map (
            O => \N__54367\,
            I => \N__53969\
        );

    \I__12619\ : LocalMux
    port map (
            O => \N__54364\,
            I => \N__53960\
        );

    \I__12618\ : LocalMux
    port map (
            O => \N__54357\,
            I => \N__53960\
        );

    \I__12617\ : LocalMux
    port map (
            O => \N__54352\,
            I => \N__53960\
        );

    \I__12616\ : InMux
    port map (
            O => \N__54351\,
            I => \N__53957\
        );

    \I__12615\ : InMux
    port map (
            O => \N__54348\,
            I => \N__53950\
        );

    \I__12614\ : InMux
    port map (
            O => \N__54347\,
            I => \N__53950\
        );

    \I__12613\ : InMux
    port map (
            O => \N__54346\,
            I => \N__53950\
        );

    \I__12612\ : InMux
    port map (
            O => \N__54345\,
            I => \N__53945\
        );

    \I__12611\ : InMux
    port map (
            O => \N__54342\,
            I => \N__53945\
        );

    \I__12610\ : InMux
    port map (
            O => \N__54339\,
            I => \N__53936\
        );

    \I__12609\ : InMux
    port map (
            O => \N__54336\,
            I => \N__53936\
        );

    \I__12608\ : InMux
    port map (
            O => \N__54333\,
            I => \N__53936\
        );

    \I__12607\ : InMux
    port map (
            O => \N__54330\,
            I => \N__53936\
        );

    \I__12606\ : CascadeMux
    port map (
            O => \N__54329\,
            I => \N__53932\
        );

    \I__12605\ : CascadeMux
    port map (
            O => \N__54328\,
            I => \N__53929\
        );

    \I__12604\ : CascadeMux
    port map (
            O => \N__54327\,
            I => \N__53926\
        );

    \I__12603\ : CascadeMux
    port map (
            O => \N__54326\,
            I => \N__53923\
        );

    \I__12602\ : CascadeMux
    port map (
            O => \N__54325\,
            I => \N__53920\
        );

    \I__12601\ : InMux
    port map (
            O => \N__54324\,
            I => \N__53910\
        );

    \I__12600\ : InMux
    port map (
            O => \N__54321\,
            I => \N__53910\
        );

    \I__12599\ : InMux
    port map (
            O => \N__54318\,
            I => \N__53910\
        );

    \I__12598\ : InMux
    port map (
            O => \N__54315\,
            I => \N__53903\
        );

    \I__12597\ : InMux
    port map (
            O => \N__54312\,
            I => \N__53903\
        );

    \I__12596\ : InMux
    port map (
            O => \N__54309\,
            I => \N__53903\
        );

    \I__12595\ : Span4Mux_v
    port map (
            O => \N__54306\,
            I => \N__53898\
        );

    \I__12594\ : LocalMux
    port map (
            O => \N__54297\,
            I => \N__53898\
        );

    \I__12593\ : InMux
    port map (
            O => \N__54294\,
            I => \N__53891\
        );

    \I__12592\ : InMux
    port map (
            O => \N__54293\,
            I => \N__53891\
        );

    \I__12591\ : InMux
    port map (
            O => \N__54292\,
            I => \N__53891\
        );

    \I__12590\ : InMux
    port map (
            O => \N__54289\,
            I => \N__53880\
        );

    \I__12589\ : InMux
    port map (
            O => \N__54288\,
            I => \N__53880\
        );

    \I__12588\ : InMux
    port map (
            O => \N__54287\,
            I => \N__53880\
        );

    \I__12587\ : InMux
    port map (
            O => \N__54284\,
            I => \N__53880\
        );

    \I__12586\ : InMux
    port map (
            O => \N__54283\,
            I => \N__53880\
        );

    \I__12585\ : Span4Mux_h
    port map (
            O => \N__54280\,
            I => \N__53875\
        );

    \I__12584\ : LocalMux
    port map (
            O => \N__54275\,
            I => \N__53875\
        );

    \I__12583\ : Span4Mux_h
    port map (
            O => \N__54270\,
            I => \N__53868\
        );

    \I__12582\ : Span4Mux_h
    port map (
            O => \N__54263\,
            I => \N__53868\
        );

    \I__12581\ : LocalMux
    port map (
            O => \N__54258\,
            I => \N__53868\
        );

    \I__12580\ : LocalMux
    port map (
            O => \N__54253\,
            I => \N__53865\
        );

    \I__12579\ : InMux
    port map (
            O => \N__54252\,
            I => \N__53856\
        );

    \I__12578\ : InMux
    port map (
            O => \N__54249\,
            I => \N__53856\
        );

    \I__12577\ : InMux
    port map (
            O => \N__54248\,
            I => \N__53856\
        );

    \I__12576\ : InMux
    port map (
            O => \N__54247\,
            I => \N__53856\
        );

    \I__12575\ : CascadeMux
    port map (
            O => \N__54246\,
            I => \N__53852\
        );

    \I__12574\ : CascadeMux
    port map (
            O => \N__54245\,
            I => \N__53847\
        );

    \I__12573\ : CascadeMux
    port map (
            O => \N__54244\,
            I => \N__53843\
        );

    \I__12572\ : CascadeMux
    port map (
            O => \N__54243\,
            I => \N__53838\
        );

    \I__12571\ : CascadeMux
    port map (
            O => \N__54242\,
            I => \N__53835\
        );

    \I__12570\ : CascadeMux
    port map (
            O => \N__54241\,
            I => \N__53831\
        );

    \I__12569\ : CascadeMux
    port map (
            O => \N__54240\,
            I => \N__53828\
        );

    \I__12568\ : InMux
    port map (
            O => \N__54237\,
            I => \N__53825\
        );

    \I__12567\ : InMux
    port map (
            O => \N__54236\,
            I => \N__53820\
        );

    \I__12566\ : InMux
    port map (
            O => \N__54233\,
            I => \N__53820\
        );

    \I__12565\ : LocalMux
    port map (
            O => \N__54230\,
            I => \N__53810\
        );

    \I__12564\ : LocalMux
    port map (
            O => \N__54223\,
            I => \N__53799\
        );

    \I__12563\ : LocalMux
    port map (
            O => \N__54218\,
            I => \N__53799\
        );

    \I__12562\ : LocalMux
    port map (
            O => \N__54215\,
            I => \N__53799\
        );

    \I__12561\ : LocalMux
    port map (
            O => \N__54212\,
            I => \N__53799\
        );

    \I__12560\ : LocalMux
    port map (
            O => \N__54205\,
            I => \N__53799\
        );

    \I__12559\ : Span4Mux_h
    port map (
            O => \N__54186\,
            I => \N__53792\
        );

    \I__12558\ : LocalMux
    port map (
            O => \N__54177\,
            I => \N__53792\
        );

    \I__12557\ : LocalMux
    port map (
            O => \N__54168\,
            I => \N__53792\
        );

    \I__12556\ : LocalMux
    port map (
            O => \N__54163\,
            I => \N__53778\
        );

    \I__12555\ : LocalMux
    port map (
            O => \N__54154\,
            I => \N__53778\
        );

    \I__12554\ : LocalMux
    port map (
            O => \N__54145\,
            I => \N__53778\
        );

    \I__12553\ : LocalMux
    port map (
            O => \N__54140\,
            I => \N__53761\
        );

    \I__12552\ : LocalMux
    port map (
            O => \N__54131\,
            I => \N__53761\
        );

    \I__12551\ : LocalMux
    port map (
            O => \N__54122\,
            I => \N__53761\
        );

    \I__12550\ : LocalMux
    port map (
            O => \N__54113\,
            I => \N__53761\
        );

    \I__12549\ : LocalMux
    port map (
            O => \N__54106\,
            I => \N__53761\
        );

    \I__12548\ : LocalMux
    port map (
            O => \N__54095\,
            I => \N__53761\
        );

    \I__12547\ : LocalMux
    port map (
            O => \N__54090\,
            I => \N__53761\
        );

    \I__12546\ : LocalMux
    port map (
            O => \N__54083\,
            I => \N__53761\
        );

    \I__12545\ : LocalMux
    port map (
            O => \N__54076\,
            I => \N__53758\
        );

    \I__12544\ : InMux
    port map (
            O => \N__54075\,
            I => \N__53753\
        );

    \I__12543\ : InMux
    port map (
            O => \N__54074\,
            I => \N__53753\
        );

    \I__12542\ : Span4Mux_v
    port map (
            O => \N__54067\,
            I => \N__53742\
        );

    \I__12541\ : Span4Mux_v
    port map (
            O => \N__54058\,
            I => \N__53742\
        );

    \I__12540\ : Span4Mux_s2_h
    port map (
            O => \N__54053\,
            I => \N__53742\
        );

    \I__12539\ : LocalMux
    port map (
            O => \N__54050\,
            I => \N__53742\
        );

    \I__12538\ : LocalMux
    port map (
            O => \N__54043\,
            I => \N__53742\
        );

    \I__12537\ : Span4Mux_v
    port map (
            O => \N__54036\,
            I => \N__53737\
        );

    \I__12536\ : LocalMux
    port map (
            O => \N__54025\,
            I => \N__53737\
        );

    \I__12535\ : InMux
    port map (
            O => \N__54024\,
            I => \N__53728\
        );

    \I__12534\ : InMux
    port map (
            O => \N__54023\,
            I => \N__53728\
        );

    \I__12533\ : InMux
    port map (
            O => \N__54022\,
            I => \N__53728\
        );

    \I__12532\ : InMux
    port map (
            O => \N__54021\,
            I => \N__53728\
        );

    \I__12531\ : InMux
    port map (
            O => \N__54020\,
            I => \N__53717\
        );

    \I__12530\ : InMux
    port map (
            O => \N__54017\,
            I => \N__53717\
        );

    \I__12529\ : InMux
    port map (
            O => \N__54014\,
            I => \N__53717\
        );

    \I__12528\ : InMux
    port map (
            O => \N__54011\,
            I => \N__53717\
        );

    \I__12527\ : InMux
    port map (
            O => \N__54010\,
            I => \N__53717\
        );

    \I__12526\ : Span4Mux_v
    port map (
            O => \N__54001\,
            I => \N__53710\
        );

    \I__12525\ : LocalMux
    port map (
            O => \N__53994\,
            I => \N__53710\
        );

    \I__12524\ : LocalMux
    port map (
            O => \N__53983\,
            I => \N__53710\
        );

    \I__12523\ : InMux
    port map (
            O => \N__53982\,
            I => \N__53705\
        );

    \I__12522\ : InMux
    port map (
            O => \N__53979\,
            I => \N__53705\
        );

    \I__12521\ : InMux
    port map (
            O => \N__53978\,
            I => \N__53696\
        );

    \I__12520\ : InMux
    port map (
            O => \N__53977\,
            I => \N__53696\
        );

    \I__12519\ : InMux
    port map (
            O => \N__53976\,
            I => \N__53696\
        );

    \I__12518\ : InMux
    port map (
            O => \N__53975\,
            I => \N__53696\
        );

    \I__12517\ : InMux
    port map (
            O => \N__53972\,
            I => \N__53689\
        );

    \I__12516\ : InMux
    port map (
            O => \N__53969\,
            I => \N__53689\
        );

    \I__12515\ : InMux
    port map (
            O => \N__53968\,
            I => \N__53689\
        );

    \I__12514\ : InMux
    port map (
            O => \N__53967\,
            I => \N__53686\
        );

    \I__12513\ : Span4Mux_h
    port map (
            O => \N__53960\,
            I => \N__53677\
        );

    \I__12512\ : LocalMux
    port map (
            O => \N__53957\,
            I => \N__53677\
        );

    \I__12511\ : LocalMux
    port map (
            O => \N__53950\,
            I => \N__53677\
        );

    \I__12510\ : LocalMux
    port map (
            O => \N__53945\,
            I => \N__53677\
        );

    \I__12509\ : LocalMux
    port map (
            O => \N__53936\,
            I => \N__53674\
        );

    \I__12508\ : InMux
    port map (
            O => \N__53935\,
            I => \N__53667\
        );

    \I__12507\ : InMux
    port map (
            O => \N__53932\,
            I => \N__53667\
        );

    \I__12506\ : InMux
    port map (
            O => \N__53929\,
            I => \N__53667\
        );

    \I__12505\ : InMux
    port map (
            O => \N__53926\,
            I => \N__53660\
        );

    \I__12504\ : InMux
    port map (
            O => \N__53923\,
            I => \N__53660\
        );

    \I__12503\ : InMux
    port map (
            O => \N__53920\,
            I => \N__53660\
        );

    \I__12502\ : CascadeMux
    port map (
            O => \N__53919\,
            I => \N__53656\
        );

    \I__12501\ : CascadeMux
    port map (
            O => \N__53918\,
            I => \N__53653\
        );

    \I__12500\ : CascadeMux
    port map (
            O => \N__53917\,
            I => \N__53650\
        );

    \I__12499\ : LocalMux
    port map (
            O => \N__53910\,
            I => \N__53635\
        );

    \I__12498\ : LocalMux
    port map (
            O => \N__53903\,
            I => \N__53635\
        );

    \I__12497\ : Sp12to4
    port map (
            O => \N__53898\,
            I => \N__53635\
        );

    \I__12496\ : LocalMux
    port map (
            O => \N__53891\,
            I => \N__53635\
        );

    \I__12495\ : LocalMux
    port map (
            O => \N__53880\,
            I => \N__53635\
        );

    \I__12494\ : Span4Mux_h
    port map (
            O => \N__53875\,
            I => \N__53630\
        );

    \I__12493\ : Span4Mux_v
    port map (
            O => \N__53868\,
            I => \N__53630\
        );

    \I__12492\ : Span4Mux_v
    port map (
            O => \N__53865\,
            I => \N__53625\
        );

    \I__12491\ : LocalMux
    port map (
            O => \N__53856\,
            I => \N__53625\
        );

    \I__12490\ : InMux
    port map (
            O => \N__53855\,
            I => \N__53616\
        );

    \I__12489\ : InMux
    port map (
            O => \N__53852\,
            I => \N__53616\
        );

    \I__12488\ : InMux
    port map (
            O => \N__53851\,
            I => \N__53616\
        );

    \I__12487\ : InMux
    port map (
            O => \N__53850\,
            I => \N__53616\
        );

    \I__12486\ : InMux
    port map (
            O => \N__53847\,
            I => \N__53605\
        );

    \I__12485\ : InMux
    port map (
            O => \N__53846\,
            I => \N__53605\
        );

    \I__12484\ : InMux
    port map (
            O => \N__53843\,
            I => \N__53605\
        );

    \I__12483\ : InMux
    port map (
            O => \N__53842\,
            I => \N__53605\
        );

    \I__12482\ : InMux
    port map (
            O => \N__53841\,
            I => \N__53605\
        );

    \I__12481\ : InMux
    port map (
            O => \N__53838\,
            I => \N__53594\
        );

    \I__12480\ : InMux
    port map (
            O => \N__53835\,
            I => \N__53594\
        );

    \I__12479\ : InMux
    port map (
            O => \N__53834\,
            I => \N__53594\
        );

    \I__12478\ : InMux
    port map (
            O => \N__53831\,
            I => \N__53594\
        );

    \I__12477\ : InMux
    port map (
            O => \N__53828\,
            I => \N__53594\
        );

    \I__12476\ : LocalMux
    port map (
            O => \N__53825\,
            I => \N__53589\
        );

    \I__12475\ : LocalMux
    port map (
            O => \N__53820\,
            I => \N__53589\
        );

    \I__12474\ : InMux
    port map (
            O => \N__53819\,
            I => \N__53586\
        );

    \I__12473\ : InMux
    port map (
            O => \N__53818\,
            I => \N__53579\
        );

    \I__12472\ : InMux
    port map (
            O => \N__53817\,
            I => \N__53579\
        );

    \I__12471\ : InMux
    port map (
            O => \N__53816\,
            I => \N__53579\
        );

    \I__12470\ : InMux
    port map (
            O => \N__53815\,
            I => \N__53572\
        );

    \I__12469\ : InMux
    port map (
            O => \N__53814\,
            I => \N__53572\
        );

    \I__12468\ : InMux
    port map (
            O => \N__53813\,
            I => \N__53572\
        );

    \I__12467\ : Span4Mux_v
    port map (
            O => \N__53810\,
            I => \N__53565\
        );

    \I__12466\ : Span4Mux_v
    port map (
            O => \N__53799\,
            I => \N__53565\
        );

    \I__12465\ : Span4Mux_v
    port map (
            O => \N__53792\,
            I => \N__53565\
        );

    \I__12464\ : InMux
    port map (
            O => \N__53791\,
            I => \N__53562\
        );

    \I__12463\ : InMux
    port map (
            O => \N__53790\,
            I => \N__53557\
        );

    \I__12462\ : InMux
    port map (
            O => \N__53789\,
            I => \N__53557\
        );

    \I__12461\ : InMux
    port map (
            O => \N__53788\,
            I => \N__53552\
        );

    \I__12460\ : InMux
    port map (
            O => \N__53787\,
            I => \N__53552\
        );

    \I__12459\ : InMux
    port map (
            O => \N__53786\,
            I => \N__53547\
        );

    \I__12458\ : InMux
    port map (
            O => \N__53785\,
            I => \N__53547\
        );

    \I__12457\ : Span4Mux_v
    port map (
            O => \N__53778\,
            I => \N__53542\
        );

    \I__12456\ : Span4Mux_v
    port map (
            O => \N__53761\,
            I => \N__53542\
        );

    \I__12455\ : Span4Mux_v
    port map (
            O => \N__53758\,
            I => \N__53537\
        );

    \I__12454\ : LocalMux
    port map (
            O => \N__53753\,
            I => \N__53537\
        );

    \I__12453\ : Span4Mux_h
    port map (
            O => \N__53742\,
            I => \N__53528\
        );

    \I__12452\ : Span4Mux_v
    port map (
            O => \N__53737\,
            I => \N__53528\
        );

    \I__12451\ : LocalMux
    port map (
            O => \N__53728\,
            I => \N__53528\
        );

    \I__12450\ : LocalMux
    port map (
            O => \N__53717\,
            I => \N__53528\
        );

    \I__12449\ : Span4Mux_v
    port map (
            O => \N__53710\,
            I => \N__53519\
        );

    \I__12448\ : LocalMux
    port map (
            O => \N__53705\,
            I => \N__53519\
        );

    \I__12447\ : LocalMux
    port map (
            O => \N__53696\,
            I => \N__53519\
        );

    \I__12446\ : LocalMux
    port map (
            O => \N__53689\,
            I => \N__53519\
        );

    \I__12445\ : LocalMux
    port map (
            O => \N__53686\,
            I => \N__53516\
        );

    \I__12444\ : Span4Mux_v
    port map (
            O => \N__53677\,
            I => \N__53513\
        );

    \I__12443\ : Span4Mux_v
    port map (
            O => \N__53674\,
            I => \N__53506\
        );

    \I__12442\ : LocalMux
    port map (
            O => \N__53667\,
            I => \N__53506\
        );

    \I__12441\ : LocalMux
    port map (
            O => \N__53660\,
            I => \N__53506\
        );

    \I__12440\ : InMux
    port map (
            O => \N__53659\,
            I => \N__53497\
        );

    \I__12439\ : InMux
    port map (
            O => \N__53656\,
            I => \N__53497\
        );

    \I__12438\ : InMux
    port map (
            O => \N__53653\,
            I => \N__53497\
        );

    \I__12437\ : InMux
    port map (
            O => \N__53650\,
            I => \N__53497\
        );

    \I__12436\ : CascadeMux
    port map (
            O => \N__53649\,
            I => \N__53494\
        );

    \I__12435\ : CascadeMux
    port map (
            O => \N__53648\,
            I => \N__53491\
        );

    \I__12434\ : CascadeMux
    port map (
            O => \N__53647\,
            I => \N__53488\
        );

    \I__12433\ : CascadeMux
    port map (
            O => \N__53646\,
            I => \N__53485\
        );

    \I__12432\ : Span12Mux_v
    port map (
            O => \N__53635\,
            I => \N__53482\
        );

    \I__12431\ : Span4Mux_v
    port map (
            O => \N__53630\,
            I => \N__53477\
        );

    \I__12430\ : Span4Mux_v
    port map (
            O => \N__53625\,
            I => \N__53477\
        );

    \I__12429\ : LocalMux
    port map (
            O => \N__53616\,
            I => \N__53472\
        );

    \I__12428\ : LocalMux
    port map (
            O => \N__53605\,
            I => \N__53472\
        );

    \I__12427\ : LocalMux
    port map (
            O => \N__53594\,
            I => \N__53461\
        );

    \I__12426\ : Span12Mux_s8_v
    port map (
            O => \N__53589\,
            I => \N__53461\
        );

    \I__12425\ : LocalMux
    port map (
            O => \N__53586\,
            I => \N__53461\
        );

    \I__12424\ : LocalMux
    port map (
            O => \N__53579\,
            I => \N__53461\
        );

    \I__12423\ : LocalMux
    port map (
            O => \N__53572\,
            I => \N__53461\
        );

    \I__12422\ : Sp12to4
    port map (
            O => \N__53565\,
            I => \N__53450\
        );

    \I__12421\ : LocalMux
    port map (
            O => \N__53562\,
            I => \N__53450\
        );

    \I__12420\ : LocalMux
    port map (
            O => \N__53557\,
            I => \N__53450\
        );

    \I__12419\ : LocalMux
    port map (
            O => \N__53552\,
            I => \N__53450\
        );

    \I__12418\ : LocalMux
    port map (
            O => \N__53547\,
            I => \N__53450\
        );

    \I__12417\ : Span4Mux_h
    port map (
            O => \N__53542\,
            I => \N__53445\
        );

    \I__12416\ : Span4Mux_v
    port map (
            O => \N__53537\,
            I => \N__53445\
        );

    \I__12415\ : Span4Mux_v
    port map (
            O => \N__53528\,
            I => \N__53440\
        );

    \I__12414\ : Span4Mux_v
    port map (
            O => \N__53519\,
            I => \N__53440\
        );

    \I__12413\ : Span12Mux_s4_h
    port map (
            O => \N__53516\,
            I => \N__53435\
        );

    \I__12412\ : Sp12to4
    port map (
            O => \N__53513\,
            I => \N__53435\
        );

    \I__12411\ : Span4Mux_h
    port map (
            O => \N__53506\,
            I => \N__53430\
        );

    \I__12410\ : LocalMux
    port map (
            O => \N__53497\,
            I => \N__53430\
        );

    \I__12409\ : InMux
    port map (
            O => \N__53494\,
            I => \N__53421\
        );

    \I__12408\ : InMux
    port map (
            O => \N__53491\,
            I => \N__53421\
        );

    \I__12407\ : InMux
    port map (
            O => \N__53488\,
            I => \N__53421\
        );

    \I__12406\ : InMux
    port map (
            O => \N__53485\,
            I => \N__53421\
        );

    \I__12405\ : Span12Mux_h
    port map (
            O => \N__53482\,
            I => \N__53418\
        );

    \I__12404\ : Span4Mux_v
    port map (
            O => \N__53477\,
            I => \N__53415\
        );

    \I__12403\ : Span12Mux_v
    port map (
            O => \N__53472\,
            I => \N__53408\
        );

    \I__12402\ : Span12Mux_h
    port map (
            O => \N__53461\,
            I => \N__53408\
        );

    \I__12401\ : Span12Mux_h
    port map (
            O => \N__53450\,
            I => \N__53408\
        );

    \I__12400\ : Span4Mux_h
    port map (
            O => \N__53445\,
            I => \N__53403\
        );

    \I__12399\ : Span4Mux_h
    port map (
            O => \N__53440\,
            I => \N__53403\
        );

    \I__12398\ : Span12Mux_v
    port map (
            O => \N__53435\,
            I => \N__53396\
        );

    \I__12397\ : Sp12to4
    port map (
            O => \N__53430\,
            I => \N__53396\
        );

    \I__12396\ : LocalMux
    port map (
            O => \N__53421\,
            I => \N__53396\
        );

    \I__12395\ : Odrv12
    port map (
            O => \N__53418\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12394\ : Odrv4
    port map (
            O => \N__53415\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12393\ : Odrv12
    port map (
            O => \N__53408\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12392\ : Odrv4
    port map (
            O => \N__53403\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12391\ : Odrv12
    port map (
            O => \N__53396\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12390\ : CascadeMux
    port map (
            O => \N__53385\,
            I => \N__53381\
        );

    \I__12389\ : CascadeMux
    port map (
            O => \N__53384\,
            I => \N__53378\
        );

    \I__12388\ : InMux
    port map (
            O => \N__53381\,
            I => \N__53374\
        );

    \I__12387\ : InMux
    port map (
            O => \N__53378\,
            I => \N__53371\
        );

    \I__12386\ : InMux
    port map (
            O => \N__53377\,
            I => \N__53368\
        );

    \I__12385\ : LocalMux
    port map (
            O => \N__53374\,
            I => \N__53365\
        );

    \I__12384\ : LocalMux
    port map (
            O => \N__53371\,
            I => n1026
        );

    \I__12383\ : LocalMux
    port map (
            O => \N__53368\,
            I => n1026
        );

    \I__12382\ : Odrv12
    port map (
            O => \N__53365\,
            I => n1026
        );

    \I__12381\ : InMux
    port map (
            O => \N__53358\,
            I => \bfn_16_24_0_\
        );

    \I__12380\ : InMux
    port map (
            O => \N__53355\,
            I => \N__53352\
        );

    \I__12379\ : LocalMux
    port map (
            O => \N__53352\,
            I => \N__53349\
        );

    \I__12378\ : Odrv4
    port map (
            O => \N__53349\,
            I => n1093
        );

    \I__12377\ : InMux
    port map (
            O => \N__53346\,
            I => \N__53342\
        );

    \I__12376\ : InMux
    port map (
            O => \N__53345\,
            I => \N__53339\
        );

    \I__12375\ : LocalMux
    port map (
            O => \N__53342\,
            I => \N__53336\
        );

    \I__12374\ : LocalMux
    port map (
            O => \N__53339\,
            I => sweep_counter_0
        );

    \I__12373\ : Odrv4
    port map (
            O => \N__53336\,
            I => sweep_counter_0
        );

    \I__12372\ : InMux
    port map (
            O => \N__53331\,
            I => \bfn_16_25_0_\
        );

    \I__12371\ : InMux
    port map (
            O => \N__53328\,
            I => \N__53324\
        );

    \I__12370\ : InMux
    port map (
            O => \N__53327\,
            I => \N__53321\
        );

    \I__12369\ : LocalMux
    port map (
            O => \N__53324\,
            I => \N__53318\
        );

    \I__12368\ : LocalMux
    port map (
            O => \N__53321\,
            I => sweep_counter_1
        );

    \I__12367\ : Odrv4
    port map (
            O => \N__53318\,
            I => sweep_counter_1
        );

    \I__12366\ : InMux
    port map (
            O => \N__53313\,
            I => n13053
        );

    \I__12365\ : InMux
    port map (
            O => \N__53310\,
            I => \N__53306\
        );

    \I__12364\ : InMux
    port map (
            O => \N__53309\,
            I => \N__53303\
        );

    \I__12363\ : LocalMux
    port map (
            O => \N__53306\,
            I => \N__53300\
        );

    \I__12362\ : LocalMux
    port map (
            O => \N__53303\,
            I => \N__53295\
        );

    \I__12361\ : Span4Mux_v
    port map (
            O => \N__53300\,
            I => \N__53295\
        );

    \I__12360\ : Odrv4
    port map (
            O => \N__53295\,
            I => sweep_counter_2
        );

    \I__12359\ : InMux
    port map (
            O => \N__53292\,
            I => n13054
        );

    \I__12358\ : InMux
    port map (
            O => \N__53289\,
            I => \N__53286\
        );

    \I__12357\ : LocalMux
    port map (
            O => \N__53286\,
            I => \N__53282\
        );

    \I__12356\ : InMux
    port map (
            O => \N__53285\,
            I => \N__53279\
        );

    \I__12355\ : Span4Mux_v
    port map (
            O => \N__53282\,
            I => \N__53276\
        );

    \I__12354\ : LocalMux
    port map (
            O => \N__53279\,
            I => sweep_counter_3
        );

    \I__12353\ : Odrv4
    port map (
            O => \N__53276\,
            I => sweep_counter_3
        );

    \I__12352\ : InMux
    port map (
            O => \N__53271\,
            I => n13055
        );

    \I__12351\ : InMux
    port map (
            O => \N__53268\,
            I => \N__53265\
        );

    \I__12350\ : LocalMux
    port map (
            O => \N__53265\,
            I => \N__53261\
        );

    \I__12349\ : InMux
    port map (
            O => \N__53264\,
            I => \N__53258\
        );

    \I__12348\ : Span4Mux_h
    port map (
            O => \N__53261\,
            I => \N__53255\
        );

    \I__12347\ : LocalMux
    port map (
            O => \N__53258\,
            I => sweep_counter_4
        );

    \I__12346\ : Odrv4
    port map (
            O => \N__53255\,
            I => sweep_counter_4
        );

    \I__12345\ : InMux
    port map (
            O => \N__53250\,
            I => n13056
        );

    \I__12344\ : InMux
    port map (
            O => \N__53247\,
            I => \N__53243\
        );

    \I__12343\ : InMux
    port map (
            O => \N__53246\,
            I => \N__53240\
        );

    \I__12342\ : LocalMux
    port map (
            O => \N__53243\,
            I => \N__53237\
        );

    \I__12341\ : LocalMux
    port map (
            O => \N__53240\,
            I => sweep_counter_5
        );

    \I__12340\ : Odrv4
    port map (
            O => \N__53237\,
            I => sweep_counter_5
        );

    \I__12339\ : InMux
    port map (
            O => \N__53232\,
            I => n13057
        );

    \I__12338\ : InMux
    port map (
            O => \N__53229\,
            I => \N__53226\
        );

    \I__12337\ : LocalMux
    port map (
            O => \N__53226\,
            I => n1298
        );

    \I__12336\ : CascadeMux
    port map (
            O => \N__53223\,
            I => \N__53218\
        );

    \I__12335\ : CascadeMux
    port map (
            O => \N__53222\,
            I => \N__53215\
        );

    \I__12334\ : CascadeMux
    port map (
            O => \N__53221\,
            I => \N__53212\
        );

    \I__12333\ : InMux
    port map (
            O => \N__53218\,
            I => \N__53209\
        );

    \I__12332\ : InMux
    port map (
            O => \N__53215\,
            I => \N__53206\
        );

    \I__12331\ : InMux
    port map (
            O => \N__53212\,
            I => \N__53203\
        );

    \I__12330\ : LocalMux
    port map (
            O => \N__53209\,
            I => \N__53200\
        );

    \I__12329\ : LocalMux
    port map (
            O => \N__53206\,
            I => n1231
        );

    \I__12328\ : LocalMux
    port map (
            O => \N__53203\,
            I => n1231
        );

    \I__12327\ : Odrv4
    port map (
            O => \N__53200\,
            I => n1231
        );

    \I__12326\ : CascadeMux
    port map (
            O => \N__53193\,
            I => \N__53190\
        );

    \I__12325\ : InMux
    port map (
            O => \N__53190\,
            I => \N__53187\
        );

    \I__12324\ : LocalMux
    port map (
            O => \N__53187\,
            I => \N__53184\
        );

    \I__12323\ : Span4Mux_v
    port map (
            O => \N__53184\,
            I => \N__53181\
        );

    \I__12322\ : Span4Mux_h
    port map (
            O => \N__53181\,
            I => \N__53176\
        );

    \I__12321\ : CascadeMux
    port map (
            O => \N__53180\,
            I => \N__53168\
        );

    \I__12320\ : CascadeMux
    port map (
            O => \N__53179\,
            I => \N__53163\
        );

    \I__12319\ : Span4Mux_h
    port map (
            O => \N__53176\,
            I => \N__53159\
        );

    \I__12318\ : InMux
    port map (
            O => \N__53175\,
            I => \N__53156\
        );

    \I__12317\ : InMux
    port map (
            O => \N__53174\,
            I => \N__53153\
        );

    \I__12316\ : InMux
    port map (
            O => \N__53173\,
            I => \N__53150\
        );

    \I__12315\ : InMux
    port map (
            O => \N__53172\,
            I => \N__53145\
        );

    \I__12314\ : InMux
    port map (
            O => \N__53171\,
            I => \N__53145\
        );

    \I__12313\ : InMux
    port map (
            O => \N__53168\,
            I => \N__53134\
        );

    \I__12312\ : InMux
    port map (
            O => \N__53167\,
            I => \N__53134\
        );

    \I__12311\ : InMux
    port map (
            O => \N__53166\,
            I => \N__53134\
        );

    \I__12310\ : InMux
    port map (
            O => \N__53163\,
            I => \N__53134\
        );

    \I__12309\ : InMux
    port map (
            O => \N__53162\,
            I => \N__53134\
        );

    \I__12308\ : Odrv4
    port map (
            O => \N__53159\,
            I => n1257
        );

    \I__12307\ : LocalMux
    port map (
            O => \N__53156\,
            I => n1257
        );

    \I__12306\ : LocalMux
    port map (
            O => \N__53153\,
            I => n1257
        );

    \I__12305\ : LocalMux
    port map (
            O => \N__53150\,
            I => n1257
        );

    \I__12304\ : LocalMux
    port map (
            O => \N__53145\,
            I => n1257
        );

    \I__12303\ : LocalMux
    port map (
            O => \N__53134\,
            I => n1257
        );

    \I__12302\ : CascadeMux
    port map (
            O => \N__53121\,
            I => \N__53118\
        );

    \I__12301\ : InMux
    port map (
            O => \N__53118\,
            I => \N__53115\
        );

    \I__12300\ : LocalMux
    port map (
            O => \N__53115\,
            I => \N__53110\
        );

    \I__12299\ : InMux
    port map (
            O => \N__53114\,
            I => \N__53107\
        );

    \I__12298\ : InMux
    port map (
            O => \N__53113\,
            I => \N__53104\
        );

    \I__12297\ : Span4Mux_h
    port map (
            O => \N__53110\,
            I => \N__53101\
        );

    \I__12296\ : LocalMux
    port map (
            O => \N__53107\,
            I => \N__53096\
        );

    \I__12295\ : LocalMux
    port map (
            O => \N__53104\,
            I => \N__53096\
        );

    \I__12294\ : Odrv4
    port map (
            O => \N__53101\,
            I => n1330
        );

    \I__12293\ : Odrv4
    port map (
            O => \N__53096\,
            I => n1330
        );

    \I__12292\ : InMux
    port map (
            O => \N__53091\,
            I => \N__53088\
        );

    \I__12291\ : LocalMux
    port map (
            O => \N__53088\,
            I => \N__53085\
        );

    \I__12290\ : Span4Mux_v
    port map (
            O => \N__53085\,
            I => \N__53080\
        );

    \I__12289\ : InMux
    port map (
            O => \N__53084\,
            I => \N__53075\
        );

    \I__12288\ : InMux
    port map (
            O => \N__53083\,
            I => \N__53075\
        );

    \I__12287\ : Odrv4
    port map (
            O => \N__53080\,
            I => n296
        );

    \I__12286\ : LocalMux
    port map (
            O => \N__53075\,
            I => n296
        );

    \I__12285\ : InMux
    port map (
            O => \N__53070\,
            I => \N__53067\
        );

    \I__12284\ : LocalMux
    port map (
            O => \N__53067\,
            I => \N__53064\
        );

    \I__12283\ : Span4Mux_h
    port map (
            O => \N__53064\,
            I => \N__53061\
        );

    \I__12282\ : Odrv4
    port map (
            O => \N__53061\,
            I => n1101
        );

    \I__12281\ : InMux
    port map (
            O => \N__53058\,
            I => \bfn_16_23_0_\
        );

    \I__12280\ : CascadeMux
    port map (
            O => \N__53055\,
            I => \N__53052\
        );

    \I__12279\ : InMux
    port map (
            O => \N__53052\,
            I => \N__53047\
        );

    \I__12278\ : InMux
    port map (
            O => \N__53051\,
            I => \N__53042\
        );

    \I__12277\ : InMux
    port map (
            O => \N__53050\,
            I => \N__53042\
        );

    \I__12276\ : LocalMux
    port map (
            O => \N__53047\,
            I => \N__53039\
        );

    \I__12275\ : LocalMux
    port map (
            O => \N__53042\,
            I => n1033
        );

    \I__12274\ : Odrv12
    port map (
            O => \N__53039\,
            I => n1033
        );

    \I__12273\ : InMux
    port map (
            O => \N__53034\,
            I => \N__53031\
        );

    \I__12272\ : LocalMux
    port map (
            O => \N__53031\,
            I => \N__53028\
        );

    \I__12271\ : Odrv12
    port map (
            O => \N__53028\,
            I => n1100
        );

    \I__12270\ : InMux
    port map (
            O => \N__53025\,
            I => n12514
        );

    \I__12269\ : CascadeMux
    port map (
            O => \N__53022\,
            I => \N__53018\
        );

    \I__12268\ : CascadeMux
    port map (
            O => \N__53021\,
            I => \N__53014\
        );

    \I__12267\ : InMux
    port map (
            O => \N__53018\,
            I => \N__53011\
        );

    \I__12266\ : InMux
    port map (
            O => \N__53017\,
            I => \N__53008\
        );

    \I__12265\ : InMux
    port map (
            O => \N__53014\,
            I => \N__53005\
        );

    \I__12264\ : LocalMux
    port map (
            O => \N__53011\,
            I => \N__53002\
        );

    \I__12263\ : LocalMux
    port map (
            O => \N__53008\,
            I => n1032
        );

    \I__12262\ : LocalMux
    port map (
            O => \N__53005\,
            I => n1032
        );

    \I__12261\ : Odrv12
    port map (
            O => \N__53002\,
            I => n1032
        );

    \I__12260\ : InMux
    port map (
            O => \N__52995\,
            I => \N__52992\
        );

    \I__12259\ : LocalMux
    port map (
            O => \N__52992\,
            I => \N__52989\
        );

    \I__12258\ : Span4Mux_h
    port map (
            O => \N__52989\,
            I => \N__52986\
        );

    \I__12257\ : Odrv4
    port map (
            O => \N__52986\,
            I => n1099
        );

    \I__12256\ : InMux
    port map (
            O => \N__52983\,
            I => n12515
        );

    \I__12255\ : CascadeMux
    port map (
            O => \N__52980\,
            I => \N__52976\
        );

    \I__12254\ : CascadeMux
    port map (
            O => \N__52979\,
            I => \N__52973\
        );

    \I__12253\ : InMux
    port map (
            O => \N__52976\,
            I => \N__52969\
        );

    \I__12252\ : InMux
    port map (
            O => \N__52973\,
            I => \N__52966\
        );

    \I__12251\ : InMux
    port map (
            O => \N__52972\,
            I => \N__52963\
        );

    \I__12250\ : LocalMux
    port map (
            O => \N__52969\,
            I => \N__52960\
        );

    \I__12249\ : LocalMux
    port map (
            O => \N__52966\,
            I => n1031
        );

    \I__12248\ : LocalMux
    port map (
            O => \N__52963\,
            I => n1031
        );

    \I__12247\ : Odrv12
    port map (
            O => \N__52960\,
            I => n1031
        );

    \I__12246\ : InMux
    port map (
            O => \N__52953\,
            I => \N__52950\
        );

    \I__12245\ : LocalMux
    port map (
            O => \N__52950\,
            I => \N__52947\
        );

    \I__12244\ : Span4Mux_h
    port map (
            O => \N__52947\,
            I => \N__52944\
        );

    \I__12243\ : Odrv4
    port map (
            O => \N__52944\,
            I => n1098
        );

    \I__12242\ : InMux
    port map (
            O => \N__52941\,
            I => n12516
        );

    \I__12241\ : CascadeMux
    port map (
            O => \N__52938\,
            I => \N__52934\
        );

    \I__12240\ : CascadeMux
    port map (
            O => \N__52937\,
            I => \N__52931\
        );

    \I__12239\ : InMux
    port map (
            O => \N__52934\,
            I => \N__52927\
        );

    \I__12238\ : InMux
    port map (
            O => \N__52931\,
            I => \N__52924\
        );

    \I__12237\ : InMux
    port map (
            O => \N__52930\,
            I => \N__52921\
        );

    \I__12236\ : LocalMux
    port map (
            O => \N__52927\,
            I => \N__52918\
        );

    \I__12235\ : LocalMux
    port map (
            O => \N__52924\,
            I => n1030
        );

    \I__12234\ : LocalMux
    port map (
            O => \N__52921\,
            I => n1030
        );

    \I__12233\ : Odrv4
    port map (
            O => \N__52918\,
            I => n1030
        );

    \I__12232\ : InMux
    port map (
            O => \N__52911\,
            I => \N__52908\
        );

    \I__12231\ : LocalMux
    port map (
            O => \N__52908\,
            I => \N__52905\
        );

    \I__12230\ : Span4Mux_h
    port map (
            O => \N__52905\,
            I => \N__52902\
        );

    \I__12229\ : Odrv4
    port map (
            O => \N__52902\,
            I => n1097
        );

    \I__12228\ : InMux
    port map (
            O => \N__52899\,
            I => n12517
        );

    \I__12227\ : CascadeMux
    port map (
            O => \N__52896\,
            I => \N__52892\
        );

    \I__12226\ : InMux
    port map (
            O => \N__52895\,
            I => \N__52889\
        );

    \I__12225\ : InMux
    port map (
            O => \N__52892\,
            I => \N__52886\
        );

    \I__12224\ : LocalMux
    port map (
            O => \N__52889\,
            I => \N__52880\
        );

    \I__12223\ : LocalMux
    port map (
            O => \N__52886\,
            I => \N__52880\
        );

    \I__12222\ : InMux
    port map (
            O => \N__52885\,
            I => \N__52877\
        );

    \I__12221\ : Span4Mux_h
    port map (
            O => \N__52880\,
            I => \N__52874\
        );

    \I__12220\ : LocalMux
    port map (
            O => \N__52877\,
            I => n1029
        );

    \I__12219\ : Odrv4
    port map (
            O => \N__52874\,
            I => n1029
        );

    \I__12218\ : InMux
    port map (
            O => \N__52869\,
            I => \N__52866\
        );

    \I__12217\ : LocalMux
    port map (
            O => \N__52866\,
            I => n1096
        );

    \I__12216\ : InMux
    port map (
            O => \N__52863\,
            I => n12518
        );

    \I__12215\ : CascadeMux
    port map (
            O => \N__52860\,
            I => \N__52856\
        );

    \I__12214\ : InMux
    port map (
            O => \N__52859\,
            I => \N__52853\
        );

    \I__12213\ : InMux
    port map (
            O => \N__52856\,
            I => \N__52849\
        );

    \I__12212\ : LocalMux
    port map (
            O => \N__52853\,
            I => \N__52846\
        );

    \I__12211\ : InMux
    port map (
            O => \N__52852\,
            I => \N__52843\
        );

    \I__12210\ : LocalMux
    port map (
            O => \N__52849\,
            I => \N__52840\
        );

    \I__12209\ : Odrv4
    port map (
            O => \N__52846\,
            I => n1028
        );

    \I__12208\ : LocalMux
    port map (
            O => \N__52843\,
            I => n1028
        );

    \I__12207\ : Odrv12
    port map (
            O => \N__52840\,
            I => n1028
        );

    \I__12206\ : InMux
    port map (
            O => \N__52833\,
            I => \N__52830\
        );

    \I__12205\ : LocalMux
    port map (
            O => \N__52830\,
            I => n1095
        );

    \I__12204\ : InMux
    port map (
            O => \N__52827\,
            I => n12519
        );

    \I__12203\ : InMux
    port map (
            O => \N__52824\,
            I => n12533
        );

    \I__12202\ : CascadeMux
    port map (
            O => \N__52821\,
            I => \N__52817\
        );

    \I__12201\ : CascadeMux
    port map (
            O => \N__52820\,
            I => \N__52814\
        );

    \I__12200\ : InMux
    port map (
            O => \N__52817\,
            I => \N__52810\
        );

    \I__12199\ : InMux
    port map (
            O => \N__52814\,
            I => \N__52807\
        );

    \I__12198\ : InMux
    port map (
            O => \N__52813\,
            I => \N__52804\
        );

    \I__12197\ : LocalMux
    port map (
            O => \N__52810\,
            I => \N__52799\
        );

    \I__12196\ : LocalMux
    port map (
            O => \N__52807\,
            I => \N__52799\
        );

    \I__12195\ : LocalMux
    port map (
            O => \N__52804\,
            I => n1230
        );

    \I__12194\ : Odrv4
    port map (
            O => \N__52799\,
            I => n1230
        );

    \I__12193\ : InMux
    port map (
            O => \N__52794\,
            I => \N__52791\
        );

    \I__12192\ : LocalMux
    port map (
            O => \N__52791\,
            I => n1297
        );

    \I__12191\ : InMux
    port map (
            O => \N__52788\,
            I => n12534
        );

    \I__12190\ : CascadeMux
    port map (
            O => \N__52785\,
            I => \N__52782\
        );

    \I__12189\ : InMux
    port map (
            O => \N__52782\,
            I => \N__52778\
        );

    \I__12188\ : InMux
    port map (
            O => \N__52781\,
            I => \N__52775\
        );

    \I__12187\ : LocalMux
    port map (
            O => \N__52778\,
            I => \N__52771\
        );

    \I__12186\ : LocalMux
    port map (
            O => \N__52775\,
            I => \N__52768\
        );

    \I__12185\ : InMux
    port map (
            O => \N__52774\,
            I => \N__52765\
        );

    \I__12184\ : Span4Mux_h
    port map (
            O => \N__52771\,
            I => \N__52762\
        );

    \I__12183\ : Odrv4
    port map (
            O => \N__52768\,
            I => n1229
        );

    \I__12182\ : LocalMux
    port map (
            O => \N__52765\,
            I => n1229
        );

    \I__12181\ : Odrv4
    port map (
            O => \N__52762\,
            I => n1229
        );

    \I__12180\ : InMux
    port map (
            O => \N__52755\,
            I => \N__52752\
        );

    \I__12179\ : LocalMux
    port map (
            O => \N__52752\,
            I => n1296
        );

    \I__12178\ : InMux
    port map (
            O => \N__52749\,
            I => n12535
        );

    \I__12177\ : CascadeMux
    port map (
            O => \N__52746\,
            I => \N__52742\
        );

    \I__12176\ : CascadeMux
    port map (
            O => \N__52745\,
            I => \N__52739\
        );

    \I__12175\ : InMux
    port map (
            O => \N__52742\,
            I => \N__52736\
        );

    \I__12174\ : InMux
    port map (
            O => \N__52739\,
            I => \N__52733\
        );

    \I__12173\ : LocalMux
    port map (
            O => \N__52736\,
            I => \N__52727\
        );

    \I__12172\ : LocalMux
    port map (
            O => \N__52733\,
            I => \N__52727\
        );

    \I__12171\ : InMux
    port map (
            O => \N__52732\,
            I => \N__52724\
        );

    \I__12170\ : Odrv4
    port map (
            O => \N__52727\,
            I => n1228
        );

    \I__12169\ : LocalMux
    port map (
            O => \N__52724\,
            I => n1228
        );

    \I__12168\ : InMux
    port map (
            O => \N__52719\,
            I => \N__52716\
        );

    \I__12167\ : LocalMux
    port map (
            O => \N__52716\,
            I => n1295
        );

    \I__12166\ : InMux
    port map (
            O => \N__52713\,
            I => n12536
        );

    \I__12165\ : CascadeMux
    port map (
            O => \N__52710\,
            I => \N__52706\
        );

    \I__12164\ : CascadeMux
    port map (
            O => \N__52709\,
            I => \N__52703\
        );

    \I__12163\ : InMux
    port map (
            O => \N__52706\,
            I => \N__52700\
        );

    \I__12162\ : InMux
    port map (
            O => \N__52703\,
            I => \N__52697\
        );

    \I__12161\ : LocalMux
    port map (
            O => \N__52700\,
            I => n1227
        );

    \I__12160\ : LocalMux
    port map (
            O => \N__52697\,
            I => n1227
        );

    \I__12159\ : InMux
    port map (
            O => \N__52692\,
            I => \N__52689\
        );

    \I__12158\ : LocalMux
    port map (
            O => \N__52689\,
            I => n1294
        );

    \I__12157\ : InMux
    port map (
            O => \N__52686\,
            I => n12537
        );

    \I__12156\ : CascadeMux
    port map (
            O => \N__52683\,
            I => \N__52680\
        );

    \I__12155\ : InMux
    port map (
            O => \N__52680\,
            I => \N__52675\
        );

    \I__12154\ : InMux
    port map (
            O => \N__52679\,
            I => \N__52670\
        );

    \I__12153\ : InMux
    port map (
            O => \N__52678\,
            I => \N__52670\
        );

    \I__12152\ : LocalMux
    port map (
            O => \N__52675\,
            I => n1226
        );

    \I__12151\ : LocalMux
    port map (
            O => \N__52670\,
            I => n1226
        );

    \I__12150\ : InMux
    port map (
            O => \N__52665\,
            I => \N__52662\
        );

    \I__12149\ : LocalMux
    port map (
            O => \N__52662\,
            I => n1293
        );

    \I__12148\ : InMux
    port map (
            O => \N__52659\,
            I => \bfn_16_22_0_\
        );

    \I__12147\ : CascadeMux
    port map (
            O => \N__52656\,
            I => \N__52653\
        );

    \I__12146\ : InMux
    port map (
            O => \N__52653\,
            I => \N__52649\
        );

    \I__12145\ : InMux
    port map (
            O => \N__52652\,
            I => \N__52646\
        );

    \I__12144\ : LocalMux
    port map (
            O => \N__52649\,
            I => n1225
        );

    \I__12143\ : LocalMux
    port map (
            O => \N__52646\,
            I => n1225
        );

    \I__12142\ : InMux
    port map (
            O => \N__52641\,
            I => \N__52638\
        );

    \I__12141\ : LocalMux
    port map (
            O => \N__52638\,
            I => n1292
        );

    \I__12140\ : InMux
    port map (
            O => \N__52635\,
            I => n12539
        );

    \I__12139\ : InMux
    port map (
            O => \N__52632\,
            I => \N__52629\
        );

    \I__12138\ : LocalMux
    port map (
            O => \N__52629\,
            I => \N__52626\
        );

    \I__12137\ : Span4Mux_v
    port map (
            O => \N__52626\,
            I => \N__52623\
        );

    \I__12136\ : Span4Mux_h
    port map (
            O => \N__52623\,
            I => \N__52620\
        );

    \I__12135\ : Span4Mux_h
    port map (
            O => \N__52620\,
            I => \N__52616\
        );

    \I__12134\ : InMux
    port map (
            O => \N__52619\,
            I => \N__52613\
        );

    \I__12133\ : Odrv4
    port map (
            O => \N__52616\,
            I => n15537
        );

    \I__12132\ : LocalMux
    port map (
            O => \N__52613\,
            I => n15537
        );

    \I__12131\ : CascadeMux
    port map (
            O => \N__52608\,
            I => \N__52605\
        );

    \I__12130\ : InMux
    port map (
            O => \N__52605\,
            I => \N__52602\
        );

    \I__12129\ : LocalMux
    port map (
            O => \N__52602\,
            I => \N__52598\
        );

    \I__12128\ : InMux
    port map (
            O => \N__52601\,
            I => \N__52595\
        );

    \I__12127\ : Span4Mux_h
    port map (
            O => \N__52598\,
            I => \N__52592\
        );

    \I__12126\ : LocalMux
    port map (
            O => \N__52595\,
            I => \N__52589\
        );

    \I__12125\ : Odrv4
    port map (
            O => \N__52592\,
            I => n1224
        );

    \I__12124\ : Odrv4
    port map (
            O => \N__52589\,
            I => n1224
        );

    \I__12123\ : InMux
    port map (
            O => \N__52584\,
            I => n12540
        );

    \I__12122\ : CascadeMux
    port map (
            O => \N__52581\,
            I => \N__52578\
        );

    \I__12121\ : InMux
    port map (
            O => \N__52578\,
            I => \N__52574\
        );

    \I__12120\ : CascadeMux
    port map (
            O => \N__52577\,
            I => \N__52571\
        );

    \I__12119\ : LocalMux
    port map (
            O => \N__52574\,
            I => \N__52568\
        );

    \I__12118\ : InMux
    port map (
            O => \N__52571\,
            I => \N__52565\
        );

    \I__12117\ : Span4Mux_h
    port map (
            O => \N__52568\,
            I => \N__52562\
        );

    \I__12116\ : LocalMux
    port map (
            O => \N__52565\,
            I => \N__52559\
        );

    \I__12115\ : Odrv4
    port map (
            O => \N__52562\,
            I => n1323
        );

    \I__12114\ : Odrv4
    port map (
            O => \N__52559\,
            I => n1323
        );

    \I__12113\ : InMux
    port map (
            O => \N__52554\,
            I => \N__52551\
        );

    \I__12112\ : LocalMux
    port map (
            O => \N__52551\,
            I => \N__52548\
        );

    \I__12111\ : Span4Mux_v
    port map (
            O => \N__52548\,
            I => \N__52545\
        );

    \I__12110\ : Span4Mux_h
    port map (
            O => \N__52545\,
            I => \N__52542\
        );

    \I__12109\ : Odrv4
    port map (
            O => \N__52542\,
            I => n1590
        );

    \I__12108\ : InMux
    port map (
            O => \N__52539\,
            I => n12574
        );

    \I__12107\ : InMux
    port map (
            O => \N__52536\,
            I => \N__52533\
        );

    \I__12106\ : LocalMux
    port map (
            O => \N__52533\,
            I => \N__52529\
        );

    \I__12105\ : InMux
    port map (
            O => \N__52532\,
            I => \N__52526\
        );

    \I__12104\ : Span4Mux_v
    port map (
            O => \N__52529\,
            I => \N__52522\
        );

    \I__12103\ : LocalMux
    port map (
            O => \N__52526\,
            I => \N__52519\
        );

    \I__12102\ : InMux
    port map (
            O => \N__52525\,
            I => \N__52516\
        );

    \I__12101\ : Odrv4
    port map (
            O => \N__52522\,
            I => n1522
        );

    \I__12100\ : Odrv4
    port map (
            O => \N__52519\,
            I => n1522
        );

    \I__12099\ : LocalMux
    port map (
            O => \N__52516\,
            I => n1522
        );

    \I__12098\ : InMux
    port map (
            O => \N__52509\,
            I => \N__52506\
        );

    \I__12097\ : LocalMux
    port map (
            O => \N__52506\,
            I => \N__52503\
        );

    \I__12096\ : Odrv4
    port map (
            O => \N__52503\,
            I => n1589
        );

    \I__12095\ : InMux
    port map (
            O => \N__52500\,
            I => n12575
        );

    \I__12094\ : InMux
    port map (
            O => \N__52497\,
            I => \N__52493\
        );

    \I__12093\ : InMux
    port map (
            O => \N__52496\,
            I => \N__52490\
        );

    \I__12092\ : LocalMux
    port map (
            O => \N__52493\,
            I => \N__52487\
        );

    \I__12091\ : LocalMux
    port map (
            O => \N__52490\,
            I => \N__52484\
        );

    \I__12090\ : Odrv4
    port map (
            O => \N__52487\,
            I => n1521
        );

    \I__12089\ : Odrv4
    port map (
            O => \N__52484\,
            I => n1521
        );

    \I__12088\ : InMux
    port map (
            O => \N__52479\,
            I => \N__52476\
        );

    \I__12087\ : LocalMux
    port map (
            O => \N__52476\,
            I => \N__52472\
        );

    \I__12086\ : CascadeMux
    port map (
            O => \N__52475\,
            I => \N__52469\
        );

    \I__12085\ : Span4Mux_v
    port map (
            O => \N__52472\,
            I => \N__52466\
        );

    \I__12084\ : InMux
    port map (
            O => \N__52469\,
            I => \N__52463\
        );

    \I__12083\ : Sp12to4
    port map (
            O => \N__52466\,
            I => \N__52460\
        );

    \I__12082\ : LocalMux
    port map (
            O => \N__52463\,
            I => \N__52457\
        );

    \I__12081\ : Span12Mux_h
    port map (
            O => \N__52460\,
            I => \N__52454\
        );

    \I__12080\ : Span4Mux_h
    port map (
            O => \N__52457\,
            I => \N__52451\
        );

    \I__12079\ : Odrv12
    port map (
            O => \N__52454\,
            I => n15591
        );

    \I__12078\ : Odrv4
    port map (
            O => \N__52451\,
            I => n15591
        );

    \I__12077\ : InMux
    port map (
            O => \N__52446\,
            I => n12576
        );

    \I__12076\ : CascadeMux
    port map (
            O => \N__52443\,
            I => \N__52440\
        );

    \I__12075\ : InMux
    port map (
            O => \N__52440\,
            I => \N__52436\
        );

    \I__12074\ : InMux
    port map (
            O => \N__52439\,
            I => \N__52433\
        );

    \I__12073\ : LocalMux
    port map (
            O => \N__52436\,
            I => \N__52430\
        );

    \I__12072\ : LocalMux
    port map (
            O => \N__52433\,
            I => \N__52427\
        );

    \I__12071\ : Span4Mux_h
    port map (
            O => \N__52430\,
            I => \N__52424\
        );

    \I__12070\ : Span4Mux_h
    port map (
            O => \N__52427\,
            I => \N__52421\
        );

    \I__12069\ : Odrv4
    port map (
            O => \N__52424\,
            I => n1620_adj_600
        );

    \I__12068\ : Odrv4
    port map (
            O => \N__52421\,
            I => n1620_adj_600
        );

    \I__12067\ : InMux
    port map (
            O => \N__52416\,
            I => \N__52413\
        );

    \I__12066\ : LocalMux
    port map (
            O => \N__52413\,
            I => \N__52410\
        );

    \I__12065\ : Span4Mux_v
    port map (
            O => \N__52410\,
            I => \N__52405\
        );

    \I__12064\ : InMux
    port map (
            O => \N__52409\,
            I => \N__52402\
        );

    \I__12063\ : InMux
    port map (
            O => \N__52408\,
            I => \N__52399\
        );

    \I__12062\ : Sp12to4
    port map (
            O => \N__52405\,
            I => \N__52394\
        );

    \I__12061\ : LocalMux
    port map (
            O => \N__52402\,
            I => \N__52394\
        );

    \I__12060\ : LocalMux
    port map (
            O => \N__52399\,
            I => encoder0_position_21
        );

    \I__12059\ : Odrv12
    port map (
            O => \N__52394\,
            I => encoder0_position_21
        );

    \I__12058\ : CascadeMux
    port map (
            O => \N__52389\,
            I => \N__52386\
        );

    \I__12057\ : InMux
    port map (
            O => \N__52386\,
            I => \N__52383\
        );

    \I__12056\ : LocalMux
    port map (
            O => \N__52383\,
            I => \N__52380\
        );

    \I__12055\ : Span4Mux_v
    port map (
            O => \N__52380\,
            I => \N__52377\
        );

    \I__12054\ : Span4Mux_h
    port map (
            O => \N__52377\,
            I => \N__52374\
        );

    \I__12053\ : Odrv4
    port map (
            O => \N__52374\,
            I => n12_adj_630
        );

    \I__12052\ : CascadeMux
    port map (
            O => \N__52371\,
            I => \N__52368\
        );

    \I__12051\ : InMux
    port map (
            O => \N__52368\,
            I => \N__52365\
        );

    \I__12050\ : LocalMux
    port map (
            O => \N__52365\,
            I => \N__52362\
        );

    \I__12049\ : Odrv12
    port map (
            O => \N__52362\,
            I => n1397
        );

    \I__12048\ : InMux
    port map (
            O => \N__52359\,
            I => \N__52356\
        );

    \I__12047\ : LocalMux
    port map (
            O => \N__52356\,
            I => \N__52353\
        );

    \I__12046\ : Span4Mux_h
    port map (
            O => \N__52353\,
            I => \N__52350\
        );

    \I__12045\ : Span4Mux_h
    port map (
            O => \N__52350\,
            I => \N__52344\
        );

    \I__12044\ : CascadeMux
    port map (
            O => \N__52349\,
            I => \N__52339\
        );

    \I__12043\ : CascadeMux
    port map (
            O => \N__52348\,
            I => \N__52333\
        );

    \I__12042\ : CascadeMux
    port map (
            O => \N__52347\,
            I => \N__52328\
        );

    \I__12041\ : Span4Mux_v
    port map (
            O => \N__52344\,
            I => \N__52324\
        );

    \I__12040\ : InMux
    port map (
            O => \N__52343\,
            I => \N__52319\
        );

    \I__12039\ : InMux
    port map (
            O => \N__52342\,
            I => \N__52319\
        );

    \I__12038\ : InMux
    port map (
            O => \N__52339\,
            I => \N__52314\
        );

    \I__12037\ : InMux
    port map (
            O => \N__52338\,
            I => \N__52314\
        );

    \I__12036\ : InMux
    port map (
            O => \N__52337\,
            I => \N__52311\
        );

    \I__12035\ : InMux
    port map (
            O => \N__52336\,
            I => \N__52304\
        );

    \I__12034\ : InMux
    port map (
            O => \N__52333\,
            I => \N__52304\
        );

    \I__12033\ : InMux
    port map (
            O => \N__52332\,
            I => \N__52304\
        );

    \I__12032\ : InMux
    port map (
            O => \N__52331\,
            I => \N__52301\
        );

    \I__12031\ : InMux
    port map (
            O => \N__52328\,
            I => \N__52296\
        );

    \I__12030\ : InMux
    port map (
            O => \N__52327\,
            I => \N__52296\
        );

    \I__12029\ : Odrv4
    port map (
            O => \N__52324\,
            I => n1356
        );

    \I__12028\ : LocalMux
    port map (
            O => \N__52319\,
            I => n1356
        );

    \I__12027\ : LocalMux
    port map (
            O => \N__52314\,
            I => n1356
        );

    \I__12026\ : LocalMux
    port map (
            O => \N__52311\,
            I => n1356
        );

    \I__12025\ : LocalMux
    port map (
            O => \N__52304\,
            I => n1356
        );

    \I__12024\ : LocalMux
    port map (
            O => \N__52301\,
            I => n1356
        );

    \I__12023\ : LocalMux
    port map (
            O => \N__52296\,
            I => n1356
        );

    \I__12022\ : CascadeMux
    port map (
            O => \N__52281\,
            I => \N__52277\
        );

    \I__12021\ : CascadeMux
    port map (
            O => \N__52280\,
            I => \N__52273\
        );

    \I__12020\ : InMux
    port map (
            O => \N__52277\,
            I => \N__52270\
        );

    \I__12019\ : InMux
    port map (
            O => \N__52276\,
            I => \N__52267\
        );

    \I__12018\ : InMux
    port map (
            O => \N__52273\,
            I => \N__52264\
        );

    \I__12017\ : LocalMux
    port map (
            O => \N__52270\,
            I => \N__52261\
        );

    \I__12016\ : LocalMux
    port map (
            O => \N__52267\,
            I => \N__52258\
        );

    \I__12015\ : LocalMux
    port map (
            O => \N__52264\,
            I => \N__52255\
        );

    \I__12014\ : Odrv4
    port map (
            O => \N__52261\,
            I => n1429
        );

    \I__12013\ : Odrv4
    port map (
            O => \N__52258\,
            I => n1429
        );

    \I__12012\ : Odrv12
    port map (
            O => \N__52255\,
            I => n1429
        );

    \I__12011\ : InMux
    port map (
            O => \N__52248\,
            I => \N__52243\
        );

    \I__12010\ : InMux
    port map (
            O => \N__52247\,
            I => \N__52240\
        );

    \I__12009\ : InMux
    port map (
            O => \N__52246\,
            I => \N__52237\
        );

    \I__12008\ : LocalMux
    port map (
            O => \N__52243\,
            I => n298
        );

    \I__12007\ : LocalMux
    port map (
            O => \N__52240\,
            I => n298
        );

    \I__12006\ : LocalMux
    port map (
            O => \N__52237\,
            I => n298
        );

    \I__12005\ : InMux
    port map (
            O => \N__52230\,
            I => \N__52227\
        );

    \I__12004\ : LocalMux
    port map (
            O => \N__52227\,
            I => \N__52224\
        );

    \I__12003\ : Odrv4
    port map (
            O => \N__52224\,
            I => n1301
        );

    \I__12002\ : InMux
    port map (
            O => \N__52221\,
            I => \bfn_16_21_0_\
        );

    \I__12001\ : CascadeMux
    port map (
            O => \N__52218\,
            I => \N__52215\
        );

    \I__12000\ : InMux
    port map (
            O => \N__52215\,
            I => \N__52211\
        );

    \I__11999\ : CascadeMux
    port map (
            O => \N__52214\,
            I => \N__52208\
        );

    \I__11998\ : LocalMux
    port map (
            O => \N__52211\,
            I => \N__52205\
        );

    \I__11997\ : InMux
    port map (
            O => \N__52208\,
            I => \N__52202\
        );

    \I__11996\ : Span4Mux_h
    port map (
            O => \N__52205\,
            I => \N__52199\
        );

    \I__11995\ : LocalMux
    port map (
            O => \N__52202\,
            I => n1233
        );

    \I__11994\ : Odrv4
    port map (
            O => \N__52199\,
            I => n1233
        );

    \I__11993\ : InMux
    port map (
            O => \N__52194\,
            I => \N__52191\
        );

    \I__11992\ : LocalMux
    port map (
            O => \N__52191\,
            I => n1300
        );

    \I__11991\ : InMux
    port map (
            O => \N__52188\,
            I => n12531
        );

    \I__11990\ : CascadeMux
    port map (
            O => \N__52185\,
            I => \N__52182\
        );

    \I__11989\ : InMux
    port map (
            O => \N__52182\,
            I => \N__52179\
        );

    \I__11988\ : LocalMux
    port map (
            O => \N__52179\,
            I => \N__52174\
        );

    \I__11987\ : InMux
    port map (
            O => \N__52178\,
            I => \N__52171\
        );

    \I__11986\ : InMux
    port map (
            O => \N__52177\,
            I => \N__52168\
        );

    \I__11985\ : Span4Mux_h
    port map (
            O => \N__52174\,
            I => \N__52165\
        );

    \I__11984\ : LocalMux
    port map (
            O => \N__52171\,
            I => n1232
        );

    \I__11983\ : LocalMux
    port map (
            O => \N__52168\,
            I => n1232
        );

    \I__11982\ : Odrv4
    port map (
            O => \N__52165\,
            I => n1232
        );

    \I__11981\ : InMux
    port map (
            O => \N__52158\,
            I => \N__52155\
        );

    \I__11980\ : LocalMux
    port map (
            O => \N__52155\,
            I => n1299
        );

    \I__11979\ : InMux
    port map (
            O => \N__52152\,
            I => n12532
        );

    \I__11978\ : CascadeMux
    port map (
            O => \N__52149\,
            I => \N__52145\
        );

    \I__11977\ : CascadeMux
    port map (
            O => \N__52148\,
            I => \N__52142\
        );

    \I__11976\ : InMux
    port map (
            O => \N__52145\,
            I => \N__52138\
        );

    \I__11975\ : InMux
    port map (
            O => \N__52142\,
            I => \N__52135\
        );

    \I__11974\ : InMux
    port map (
            O => \N__52141\,
            I => \N__52132\
        );

    \I__11973\ : LocalMux
    port map (
            O => \N__52138\,
            I => n1530
        );

    \I__11972\ : LocalMux
    port map (
            O => \N__52135\,
            I => n1530
        );

    \I__11971\ : LocalMux
    port map (
            O => \N__52132\,
            I => n1530
        );

    \I__11970\ : InMux
    port map (
            O => \N__52125\,
            I => \N__52122\
        );

    \I__11969\ : LocalMux
    port map (
            O => \N__52122\,
            I => \N__52119\
        );

    \I__11968\ : Span4Mux_h
    port map (
            O => \N__52119\,
            I => \N__52116\
        );

    \I__11967\ : Odrv4
    port map (
            O => \N__52116\,
            I => n1597
        );

    \I__11966\ : InMux
    port map (
            O => \N__52113\,
            I => n12567
        );

    \I__11965\ : CascadeMux
    port map (
            O => \N__52110\,
            I => \N__52106\
        );

    \I__11964\ : InMux
    port map (
            O => \N__52109\,
            I => \N__52102\
        );

    \I__11963\ : InMux
    port map (
            O => \N__52106\,
            I => \N__52099\
        );

    \I__11962\ : InMux
    port map (
            O => \N__52105\,
            I => \N__52096\
        );

    \I__11961\ : LocalMux
    port map (
            O => \N__52102\,
            I => n1529
        );

    \I__11960\ : LocalMux
    port map (
            O => \N__52099\,
            I => n1529
        );

    \I__11959\ : LocalMux
    port map (
            O => \N__52096\,
            I => n1529
        );

    \I__11958\ : InMux
    port map (
            O => \N__52089\,
            I => \N__52086\
        );

    \I__11957\ : LocalMux
    port map (
            O => \N__52086\,
            I => \N__52083\
        );

    \I__11956\ : Odrv4
    port map (
            O => \N__52083\,
            I => n1596
        );

    \I__11955\ : InMux
    port map (
            O => \N__52080\,
            I => n12568
        );

    \I__11954\ : CascadeMux
    port map (
            O => \N__52077\,
            I => \N__52072\
        );

    \I__11953\ : CascadeMux
    port map (
            O => \N__52076\,
            I => \N__52069\
        );

    \I__11952\ : CascadeMux
    port map (
            O => \N__52075\,
            I => \N__52066\
        );

    \I__11951\ : InMux
    port map (
            O => \N__52072\,
            I => \N__52063\
        );

    \I__11950\ : InMux
    port map (
            O => \N__52069\,
            I => \N__52060\
        );

    \I__11949\ : InMux
    port map (
            O => \N__52066\,
            I => \N__52057\
        );

    \I__11948\ : LocalMux
    port map (
            O => \N__52063\,
            I => n1528
        );

    \I__11947\ : LocalMux
    port map (
            O => \N__52060\,
            I => n1528
        );

    \I__11946\ : LocalMux
    port map (
            O => \N__52057\,
            I => n1528
        );

    \I__11945\ : InMux
    port map (
            O => \N__52050\,
            I => \N__52047\
        );

    \I__11944\ : LocalMux
    port map (
            O => \N__52047\,
            I => \N__52044\
        );

    \I__11943\ : Span4Mux_h
    port map (
            O => \N__52044\,
            I => \N__52041\
        );

    \I__11942\ : Odrv4
    port map (
            O => \N__52041\,
            I => n1595
        );

    \I__11941\ : InMux
    port map (
            O => \N__52038\,
            I => n12569
        );

    \I__11940\ : CascadeMux
    port map (
            O => \N__52035\,
            I => \N__52031\
        );

    \I__11939\ : CascadeMux
    port map (
            O => \N__52034\,
            I => \N__52028\
        );

    \I__11938\ : InMux
    port map (
            O => \N__52031\,
            I => \N__52024\
        );

    \I__11937\ : InMux
    port map (
            O => \N__52028\,
            I => \N__52021\
        );

    \I__11936\ : InMux
    port map (
            O => \N__52027\,
            I => \N__52018\
        );

    \I__11935\ : LocalMux
    port map (
            O => \N__52024\,
            I => n1527
        );

    \I__11934\ : LocalMux
    port map (
            O => \N__52021\,
            I => n1527
        );

    \I__11933\ : LocalMux
    port map (
            O => \N__52018\,
            I => n1527
        );

    \I__11932\ : InMux
    port map (
            O => \N__52011\,
            I => \N__52008\
        );

    \I__11931\ : LocalMux
    port map (
            O => \N__52008\,
            I => \N__52005\
        );

    \I__11930\ : Odrv12
    port map (
            O => \N__52005\,
            I => n1594
        );

    \I__11929\ : InMux
    port map (
            O => \N__52002\,
            I => n12570
        );

    \I__11928\ : CascadeMux
    port map (
            O => \N__51999\,
            I => \N__51996\
        );

    \I__11927\ : InMux
    port map (
            O => \N__51996\,
            I => \N__51993\
        );

    \I__11926\ : LocalMux
    port map (
            O => \N__51993\,
            I => \N__51989\
        );

    \I__11925\ : InMux
    port map (
            O => \N__51992\,
            I => \N__51986\
        );

    \I__11924\ : Span4Mux_v
    port map (
            O => \N__51989\,
            I => \N__51982\
        );

    \I__11923\ : LocalMux
    port map (
            O => \N__51986\,
            I => \N__51979\
        );

    \I__11922\ : InMux
    port map (
            O => \N__51985\,
            I => \N__51976\
        );

    \I__11921\ : Odrv4
    port map (
            O => \N__51982\,
            I => n1526
        );

    \I__11920\ : Odrv4
    port map (
            O => \N__51979\,
            I => n1526
        );

    \I__11919\ : LocalMux
    port map (
            O => \N__51976\,
            I => n1526
        );

    \I__11918\ : InMux
    port map (
            O => \N__51969\,
            I => \N__51966\
        );

    \I__11917\ : LocalMux
    port map (
            O => \N__51966\,
            I => \N__51963\
        );

    \I__11916\ : Span4Mux_v
    port map (
            O => \N__51963\,
            I => \N__51960\
        );

    \I__11915\ : Odrv4
    port map (
            O => \N__51960\,
            I => n1593
        );

    \I__11914\ : InMux
    port map (
            O => \N__51957\,
            I => \bfn_16_20_0_\
        );

    \I__11913\ : CascadeMux
    port map (
            O => \N__51954\,
            I => \N__51950\
        );

    \I__11912\ : CascadeMux
    port map (
            O => \N__51953\,
            I => \N__51947\
        );

    \I__11911\ : InMux
    port map (
            O => \N__51950\,
            I => \N__51944\
        );

    \I__11910\ : InMux
    port map (
            O => \N__51947\,
            I => \N__51940\
        );

    \I__11909\ : LocalMux
    port map (
            O => \N__51944\,
            I => \N__51937\
        );

    \I__11908\ : InMux
    port map (
            O => \N__51943\,
            I => \N__51934\
        );

    \I__11907\ : LocalMux
    port map (
            O => \N__51940\,
            I => n1525
        );

    \I__11906\ : Odrv4
    port map (
            O => \N__51937\,
            I => n1525
        );

    \I__11905\ : LocalMux
    port map (
            O => \N__51934\,
            I => n1525
        );

    \I__11904\ : InMux
    port map (
            O => \N__51927\,
            I => \N__51924\
        );

    \I__11903\ : LocalMux
    port map (
            O => \N__51924\,
            I => \N__51921\
        );

    \I__11902\ : Span4Mux_h
    port map (
            O => \N__51921\,
            I => \N__51918\
        );

    \I__11901\ : Odrv4
    port map (
            O => \N__51918\,
            I => n1592
        );

    \I__11900\ : InMux
    port map (
            O => \N__51915\,
            I => n12572
        );

    \I__11899\ : CascadeMux
    port map (
            O => \N__51912\,
            I => \N__51909\
        );

    \I__11898\ : InMux
    port map (
            O => \N__51909\,
            I => \N__51906\
        );

    \I__11897\ : LocalMux
    port map (
            O => \N__51906\,
            I => \N__51901\
        );

    \I__11896\ : InMux
    port map (
            O => \N__51905\,
            I => \N__51896\
        );

    \I__11895\ : InMux
    port map (
            O => \N__51904\,
            I => \N__51896\
        );

    \I__11894\ : Odrv4
    port map (
            O => \N__51901\,
            I => n1524
        );

    \I__11893\ : LocalMux
    port map (
            O => \N__51896\,
            I => n1524
        );

    \I__11892\ : InMux
    port map (
            O => \N__51891\,
            I => \N__51888\
        );

    \I__11891\ : LocalMux
    port map (
            O => \N__51888\,
            I => \N__51885\
        );

    \I__11890\ : Span4Mux_h
    port map (
            O => \N__51885\,
            I => \N__51882\
        );

    \I__11889\ : Odrv4
    port map (
            O => \N__51882\,
            I => n1591
        );

    \I__11888\ : InMux
    port map (
            O => \N__51879\,
            I => n12573
        );

    \I__11887\ : CascadeMux
    port map (
            O => \N__51876\,
            I => \N__51873\
        );

    \I__11886\ : InMux
    port map (
            O => \N__51873\,
            I => \N__51870\
        );

    \I__11885\ : LocalMux
    port map (
            O => \N__51870\,
            I => \N__51867\
        );

    \I__11884\ : Span4Mux_v
    port map (
            O => \N__51867\,
            I => \N__51863\
        );

    \I__11883\ : InMux
    port map (
            O => \N__51866\,
            I => \N__51860\
        );

    \I__11882\ : Odrv4
    port map (
            O => \N__51863\,
            I => n1523
        );

    \I__11881\ : LocalMux
    port map (
            O => \N__51860\,
            I => n1523
        );

    \I__11880\ : InMux
    port map (
            O => \N__51855\,
            I => \N__51851\
        );

    \I__11879\ : InMux
    port map (
            O => \N__51854\,
            I => \N__51848\
        );

    \I__11878\ : LocalMux
    port map (
            O => \N__51851\,
            I => n1425
        );

    \I__11877\ : LocalMux
    port map (
            O => \N__51848\,
            I => n1425
        );

    \I__11876\ : InMux
    port map (
            O => \N__51843\,
            I => \N__51840\
        );

    \I__11875\ : LocalMux
    port map (
            O => \N__51840\,
            I => n1492
        );

    \I__11874\ : InMux
    port map (
            O => \N__51837\,
            I => n12560
        );

    \I__11873\ : CascadeMux
    port map (
            O => \N__51834\,
            I => \N__51830\
        );

    \I__11872\ : CascadeMux
    port map (
            O => \N__51833\,
            I => \N__51827\
        );

    \I__11871\ : InMux
    port map (
            O => \N__51830\,
            I => \N__51824\
        );

    \I__11870\ : InMux
    port map (
            O => \N__51827\,
            I => \N__51821\
        );

    \I__11869\ : LocalMux
    port map (
            O => \N__51824\,
            I => \N__51816\
        );

    \I__11868\ : LocalMux
    port map (
            O => \N__51821\,
            I => \N__51816\
        );

    \I__11867\ : Span4Mux_h
    port map (
            O => \N__51816\,
            I => \N__51812\
        );

    \I__11866\ : InMux
    port map (
            O => \N__51815\,
            I => \N__51809\
        );

    \I__11865\ : Odrv4
    port map (
            O => \N__51812\,
            I => n1424
        );

    \I__11864\ : LocalMux
    port map (
            O => \N__51809\,
            I => n1424
        );

    \I__11863\ : InMux
    port map (
            O => \N__51804\,
            I => \N__51801\
        );

    \I__11862\ : LocalMux
    port map (
            O => \N__51801\,
            I => \N__51798\
        );

    \I__11861\ : Odrv4
    port map (
            O => \N__51798\,
            I => n1491
        );

    \I__11860\ : InMux
    port map (
            O => \N__51795\,
            I => n12561
        );

    \I__11859\ : CascadeMux
    port map (
            O => \N__51792\,
            I => \N__51788\
        );

    \I__11858\ : InMux
    port map (
            O => \N__51791\,
            I => \N__51785\
        );

    \I__11857\ : InMux
    port map (
            O => \N__51788\,
            I => \N__51782\
        );

    \I__11856\ : LocalMux
    port map (
            O => \N__51785\,
            I => \N__51778\
        );

    \I__11855\ : LocalMux
    port map (
            O => \N__51782\,
            I => \N__51775\
        );

    \I__11854\ : InMux
    port map (
            O => \N__51781\,
            I => \N__51772\
        );

    \I__11853\ : Odrv4
    port map (
            O => \N__51778\,
            I => n1423
        );

    \I__11852\ : Odrv4
    port map (
            O => \N__51775\,
            I => n1423
        );

    \I__11851\ : LocalMux
    port map (
            O => \N__51772\,
            I => n1423
        );

    \I__11850\ : CascadeMux
    port map (
            O => \N__51765\,
            I => \N__51762\
        );

    \I__11849\ : InMux
    port map (
            O => \N__51762\,
            I => \N__51759\
        );

    \I__11848\ : LocalMux
    port map (
            O => \N__51759\,
            I => n1490
        );

    \I__11847\ : InMux
    port map (
            O => \N__51756\,
            I => n12562
        );

    \I__11846\ : InMux
    port map (
            O => \N__51753\,
            I => \N__51750\
        );

    \I__11845\ : LocalMux
    port map (
            O => \N__51750\,
            I => \N__51747\
        );

    \I__11844\ : Span12Mux_h
    port map (
            O => \N__51747\,
            I => \N__51743\
        );

    \I__11843\ : InMux
    port map (
            O => \N__51746\,
            I => \N__51740\
        );

    \I__11842\ : Odrv12
    port map (
            O => \N__51743\,
            I => n15572
        );

    \I__11841\ : LocalMux
    port map (
            O => \N__51740\,
            I => n15572
        );

    \I__11840\ : CascadeMux
    port map (
            O => \N__51735\,
            I => \N__51732\
        );

    \I__11839\ : InMux
    port map (
            O => \N__51732\,
            I => \N__51729\
        );

    \I__11838\ : LocalMux
    port map (
            O => \N__51729\,
            I => \N__51725\
        );

    \I__11837\ : InMux
    port map (
            O => \N__51728\,
            I => \N__51722\
        );

    \I__11836\ : Span4Mux_h
    port map (
            O => \N__51725\,
            I => \N__51717\
        );

    \I__11835\ : LocalMux
    port map (
            O => \N__51722\,
            I => \N__51717\
        );

    \I__11834\ : Odrv4
    port map (
            O => \N__51717\,
            I => n1422
        );

    \I__11833\ : InMux
    port map (
            O => \N__51714\,
            I => n12563
        );

    \I__11832\ : InMux
    port map (
            O => \N__51711\,
            I => \N__51707\
        );

    \I__11831\ : InMux
    port map (
            O => \N__51710\,
            I => \N__51703\
        );

    \I__11830\ : LocalMux
    port map (
            O => \N__51707\,
            I => \N__51700\
        );

    \I__11829\ : InMux
    port map (
            O => \N__51706\,
            I => \N__51697\
        );

    \I__11828\ : LocalMux
    port map (
            O => \N__51703\,
            I => \N__51694\
        );

    \I__11827\ : Span4Mux_h
    port map (
            O => \N__51700\,
            I => \N__51689\
        );

    \I__11826\ : LocalMux
    port map (
            O => \N__51697\,
            I => \N__51689\
        );

    \I__11825\ : Span12Mux_v
    port map (
            O => \N__51694\,
            I => \N__51686\
        );

    \I__11824\ : Span4Mux_h
    port map (
            O => \N__51689\,
            I => \N__51683\
        );

    \I__11823\ : Odrv12
    port map (
            O => \N__51686\,
            I => n301
        );

    \I__11822\ : Odrv4
    port map (
            O => \N__51683\,
            I => n301
        );

    \I__11821\ : InMux
    port map (
            O => \N__51678\,
            I => \N__51675\
        );

    \I__11820\ : LocalMux
    port map (
            O => \N__51675\,
            I => \N__51672\
        );

    \I__11819\ : Span4Mux_h
    port map (
            O => \N__51672\,
            I => \N__51669\
        );

    \I__11818\ : Odrv4
    port map (
            O => \N__51669\,
            I => n1601
        );

    \I__11817\ : InMux
    port map (
            O => \N__51666\,
            I => \bfn_16_19_0_\
        );

    \I__11816\ : CascadeMux
    port map (
            O => \N__51663\,
            I => \N__51659\
        );

    \I__11815\ : InMux
    port map (
            O => \N__51662\,
            I => \N__51655\
        );

    \I__11814\ : InMux
    port map (
            O => \N__51659\,
            I => \N__51652\
        );

    \I__11813\ : InMux
    port map (
            O => \N__51658\,
            I => \N__51649\
        );

    \I__11812\ : LocalMux
    port map (
            O => \N__51655\,
            I => n1533
        );

    \I__11811\ : LocalMux
    port map (
            O => \N__51652\,
            I => n1533
        );

    \I__11810\ : LocalMux
    port map (
            O => \N__51649\,
            I => n1533
        );

    \I__11809\ : CascadeMux
    port map (
            O => \N__51642\,
            I => \N__51639\
        );

    \I__11808\ : InMux
    port map (
            O => \N__51639\,
            I => \N__51636\
        );

    \I__11807\ : LocalMux
    port map (
            O => \N__51636\,
            I => \N__51633\
        );

    \I__11806\ : Odrv4
    port map (
            O => \N__51633\,
            I => n1600
        );

    \I__11805\ : InMux
    port map (
            O => \N__51630\,
            I => n12564
        );

    \I__11804\ : CascadeMux
    port map (
            O => \N__51627\,
            I => \N__51623\
        );

    \I__11803\ : InMux
    port map (
            O => \N__51626\,
            I => \N__51619\
        );

    \I__11802\ : InMux
    port map (
            O => \N__51623\,
            I => \N__51616\
        );

    \I__11801\ : InMux
    port map (
            O => \N__51622\,
            I => \N__51613\
        );

    \I__11800\ : LocalMux
    port map (
            O => \N__51619\,
            I => n1532
        );

    \I__11799\ : LocalMux
    port map (
            O => \N__51616\,
            I => n1532
        );

    \I__11798\ : LocalMux
    port map (
            O => \N__51613\,
            I => n1532
        );

    \I__11797\ : InMux
    port map (
            O => \N__51606\,
            I => \N__51603\
        );

    \I__11796\ : LocalMux
    port map (
            O => \N__51603\,
            I => \N__51600\
        );

    \I__11795\ : Odrv4
    port map (
            O => \N__51600\,
            I => n1599
        );

    \I__11794\ : InMux
    port map (
            O => \N__51597\,
            I => n12565
        );

    \I__11793\ : CascadeMux
    port map (
            O => \N__51594\,
            I => \N__51591\
        );

    \I__11792\ : InMux
    port map (
            O => \N__51591\,
            I => \N__51587\
        );

    \I__11791\ : CascadeMux
    port map (
            O => \N__51590\,
            I => \N__51584\
        );

    \I__11790\ : LocalMux
    port map (
            O => \N__51587\,
            I => \N__51581\
        );

    \I__11789\ : InMux
    port map (
            O => \N__51584\,
            I => \N__51578\
        );

    \I__11788\ : Odrv4
    port map (
            O => \N__51581\,
            I => n1531
        );

    \I__11787\ : LocalMux
    port map (
            O => \N__51578\,
            I => n1531
        );

    \I__11786\ : InMux
    port map (
            O => \N__51573\,
            I => \N__51570\
        );

    \I__11785\ : LocalMux
    port map (
            O => \N__51570\,
            I => \N__51567\
        );

    \I__11784\ : Span4Mux_v
    port map (
            O => \N__51567\,
            I => \N__51564\
        );

    \I__11783\ : Odrv4
    port map (
            O => \N__51564\,
            I => n1598
        );

    \I__11782\ : InMux
    port map (
            O => \N__51561\,
            I => n12566
        );

    \I__11781\ : CascadeMux
    port map (
            O => \N__51558\,
            I => \N__51554\
        );

    \I__11780\ : CascadeMux
    port map (
            O => \N__51557\,
            I => \N__51551\
        );

    \I__11779\ : InMux
    port map (
            O => \N__51554\,
            I => \N__51548\
        );

    \I__11778\ : InMux
    port map (
            O => \N__51551\,
            I => \N__51545\
        );

    \I__11777\ : LocalMux
    port map (
            O => \N__51548\,
            I => \N__51542\
        );

    \I__11776\ : LocalMux
    port map (
            O => \N__51545\,
            I => \N__51539\
        );

    \I__11775\ : Span4Mux_h
    port map (
            O => \N__51542\,
            I => \N__51535\
        );

    \I__11774\ : Span4Mux_h
    port map (
            O => \N__51539\,
            I => \N__51532\
        );

    \I__11773\ : InMux
    port map (
            O => \N__51538\,
            I => \N__51529\
        );

    \I__11772\ : Span4Mux_v
    port map (
            O => \N__51535\,
            I => \N__51526\
        );

    \I__11771\ : Odrv4
    port map (
            O => \N__51532\,
            I => n1433
        );

    \I__11770\ : LocalMux
    port map (
            O => \N__51529\,
            I => n1433
        );

    \I__11769\ : Odrv4
    port map (
            O => \N__51526\,
            I => n1433
        );

    \I__11768\ : InMux
    port map (
            O => \N__51519\,
            I => \N__51516\
        );

    \I__11767\ : LocalMux
    port map (
            O => \N__51516\,
            I => n1500
        );

    \I__11766\ : InMux
    port map (
            O => \N__51513\,
            I => n12552
        );

    \I__11765\ : CascadeMux
    port map (
            O => \N__51510\,
            I => \N__51507\
        );

    \I__11764\ : InMux
    port map (
            O => \N__51507\,
            I => \N__51504\
        );

    \I__11763\ : LocalMux
    port map (
            O => \N__51504\,
            I => \N__51500\
        );

    \I__11762\ : InMux
    port map (
            O => \N__51503\,
            I => \N__51497\
        );

    \I__11761\ : Span4Mux_v
    port map (
            O => \N__51500\,
            I => \N__51494\
        );

    \I__11760\ : LocalMux
    port map (
            O => \N__51497\,
            I => n1432
        );

    \I__11759\ : Odrv4
    port map (
            O => \N__51494\,
            I => n1432
        );

    \I__11758\ : InMux
    port map (
            O => \N__51489\,
            I => \N__51486\
        );

    \I__11757\ : LocalMux
    port map (
            O => \N__51486\,
            I => \N__51483\
        );

    \I__11756\ : Odrv4
    port map (
            O => \N__51483\,
            I => n1499
        );

    \I__11755\ : InMux
    port map (
            O => \N__51480\,
            I => n12553
        );

    \I__11754\ : CascadeMux
    port map (
            O => \N__51477\,
            I => \N__51473\
        );

    \I__11753\ : InMux
    port map (
            O => \N__51476\,
            I => \N__51470\
        );

    \I__11752\ : InMux
    port map (
            O => \N__51473\,
            I => \N__51467\
        );

    \I__11751\ : LocalMux
    port map (
            O => \N__51470\,
            I => \N__51461\
        );

    \I__11750\ : LocalMux
    port map (
            O => \N__51467\,
            I => \N__51461\
        );

    \I__11749\ : InMux
    port map (
            O => \N__51466\,
            I => \N__51458\
        );

    \I__11748\ : Span4Mux_v
    port map (
            O => \N__51461\,
            I => \N__51455\
        );

    \I__11747\ : LocalMux
    port map (
            O => \N__51458\,
            I => n1431
        );

    \I__11746\ : Odrv4
    port map (
            O => \N__51455\,
            I => n1431
        );

    \I__11745\ : InMux
    port map (
            O => \N__51450\,
            I => \N__51447\
        );

    \I__11744\ : LocalMux
    port map (
            O => \N__51447\,
            I => n1498
        );

    \I__11743\ : InMux
    port map (
            O => \N__51444\,
            I => n12554
        );

    \I__11742\ : CascadeMux
    port map (
            O => \N__51441\,
            I => \N__51437\
        );

    \I__11741\ : CascadeMux
    port map (
            O => \N__51440\,
            I => \N__51434\
        );

    \I__11740\ : InMux
    port map (
            O => \N__51437\,
            I => \N__51431\
        );

    \I__11739\ : InMux
    port map (
            O => \N__51434\,
            I => \N__51428\
        );

    \I__11738\ : LocalMux
    port map (
            O => \N__51431\,
            I => \N__51425\
        );

    \I__11737\ : LocalMux
    port map (
            O => \N__51428\,
            I => n1430
        );

    \I__11736\ : Odrv4
    port map (
            O => \N__51425\,
            I => n1430
        );

    \I__11735\ : InMux
    port map (
            O => \N__51420\,
            I => \N__51417\
        );

    \I__11734\ : LocalMux
    port map (
            O => \N__51417\,
            I => \N__51414\
        );

    \I__11733\ : Odrv4
    port map (
            O => \N__51414\,
            I => n1497
        );

    \I__11732\ : InMux
    port map (
            O => \N__51411\,
            I => n12555
        );

    \I__11731\ : InMux
    port map (
            O => \N__51408\,
            I => \N__51405\
        );

    \I__11730\ : LocalMux
    port map (
            O => \N__51405\,
            I => n1496
        );

    \I__11729\ : InMux
    port map (
            O => \N__51402\,
            I => n12556
        );

    \I__11728\ : CascadeMux
    port map (
            O => \N__51399\,
            I => \N__51396\
        );

    \I__11727\ : InMux
    port map (
            O => \N__51396\,
            I => \N__51393\
        );

    \I__11726\ : LocalMux
    port map (
            O => \N__51393\,
            I => \N__51389\
        );

    \I__11725\ : InMux
    port map (
            O => \N__51392\,
            I => \N__51385\
        );

    \I__11724\ : Span4Mux_h
    port map (
            O => \N__51389\,
            I => \N__51382\
        );

    \I__11723\ : InMux
    port map (
            O => \N__51388\,
            I => \N__51379\
        );

    \I__11722\ : LocalMux
    port map (
            O => \N__51385\,
            I => n1428
        );

    \I__11721\ : Odrv4
    port map (
            O => \N__51382\,
            I => n1428
        );

    \I__11720\ : LocalMux
    port map (
            O => \N__51379\,
            I => n1428
        );

    \I__11719\ : InMux
    port map (
            O => \N__51372\,
            I => \N__51369\
        );

    \I__11718\ : LocalMux
    port map (
            O => \N__51369\,
            I => n1495
        );

    \I__11717\ : InMux
    port map (
            O => \N__51366\,
            I => n12557
        );

    \I__11716\ : CascadeMux
    port map (
            O => \N__51363\,
            I => \N__51360\
        );

    \I__11715\ : InMux
    port map (
            O => \N__51360\,
            I => \N__51357\
        );

    \I__11714\ : LocalMux
    port map (
            O => \N__51357\,
            I => \N__51353\
        );

    \I__11713\ : InMux
    port map (
            O => \N__51356\,
            I => \N__51350\
        );

    \I__11712\ : Span4Mux_h
    port map (
            O => \N__51353\,
            I => \N__51347\
        );

    \I__11711\ : LocalMux
    port map (
            O => \N__51350\,
            I => n1427
        );

    \I__11710\ : Odrv4
    port map (
            O => \N__51347\,
            I => n1427
        );

    \I__11709\ : InMux
    port map (
            O => \N__51342\,
            I => \N__51339\
        );

    \I__11708\ : LocalMux
    port map (
            O => \N__51339\,
            I => n1494
        );

    \I__11707\ : InMux
    port map (
            O => \N__51336\,
            I => n12558
        );

    \I__11706\ : InMux
    port map (
            O => \N__51333\,
            I => \N__51329\
        );

    \I__11705\ : CascadeMux
    port map (
            O => \N__51332\,
            I => \N__51326\
        );

    \I__11704\ : LocalMux
    port map (
            O => \N__51329\,
            I => \N__51322\
        );

    \I__11703\ : InMux
    port map (
            O => \N__51326\,
            I => \N__51319\
        );

    \I__11702\ : InMux
    port map (
            O => \N__51325\,
            I => \N__51316\
        );

    \I__11701\ : Odrv4
    port map (
            O => \N__51322\,
            I => n1426
        );

    \I__11700\ : LocalMux
    port map (
            O => \N__51319\,
            I => n1426
        );

    \I__11699\ : LocalMux
    port map (
            O => \N__51316\,
            I => n1426
        );

    \I__11698\ : InMux
    port map (
            O => \N__51309\,
            I => \N__51306\
        );

    \I__11697\ : LocalMux
    port map (
            O => \N__51306\,
            I => n1493
        );

    \I__11696\ : InMux
    port map (
            O => \N__51303\,
            I => \bfn_16_18_0_\
        );

    \I__11695\ : CascadeMux
    port map (
            O => \N__51300\,
            I => \N__51297\
        );

    \I__11694\ : InMux
    port map (
            O => \N__51297\,
            I => \N__51293\
        );

    \I__11693\ : InMux
    port map (
            O => \N__51296\,
            I => \N__51288\
        );

    \I__11692\ : LocalMux
    port map (
            O => \N__51293\,
            I => \N__51285\
        );

    \I__11691\ : InMux
    port map (
            O => \N__51292\,
            I => \N__51280\
        );

    \I__11690\ : InMux
    port map (
            O => \N__51291\,
            I => \N__51280\
        );

    \I__11689\ : LocalMux
    port map (
            O => \N__51288\,
            I => encoder0_position_target_20
        );

    \I__11688\ : Odrv4
    port map (
            O => \N__51285\,
            I => encoder0_position_target_20
        );

    \I__11687\ : LocalMux
    port map (
            O => \N__51280\,
            I => encoder0_position_target_20
        );

    \I__11686\ : InMux
    port map (
            O => \N__51273\,
            I => n12469
        );

    \I__11685\ : CascadeMux
    port map (
            O => \N__51270\,
            I => \N__51267\
        );

    \I__11684\ : InMux
    port map (
            O => \N__51267\,
            I => \N__51261\
        );

    \I__11683\ : InMux
    port map (
            O => \N__51266\,
            I => \N__51256\
        );

    \I__11682\ : InMux
    port map (
            O => \N__51265\,
            I => \N__51256\
        );

    \I__11681\ : CascadeMux
    port map (
            O => \N__51264\,
            I => \N__51253\
        );

    \I__11680\ : LocalMux
    port map (
            O => \N__51261\,
            I => \N__51250\
        );

    \I__11679\ : LocalMux
    port map (
            O => \N__51256\,
            I => \N__51247\
        );

    \I__11678\ : InMux
    port map (
            O => \N__51253\,
            I => \N__51244\
        );

    \I__11677\ : Span4Mux_h
    port map (
            O => \N__51250\,
            I => \N__51241\
        );

    \I__11676\ : Span4Mux_h
    port map (
            O => \N__51247\,
            I => \N__51238\
        );

    \I__11675\ : LocalMux
    port map (
            O => \N__51244\,
            I => encoder0_position_target_21
        );

    \I__11674\ : Odrv4
    port map (
            O => \N__51241\,
            I => encoder0_position_target_21
        );

    \I__11673\ : Odrv4
    port map (
            O => \N__51238\,
            I => encoder0_position_target_21
        );

    \I__11672\ : InMux
    port map (
            O => \N__51231\,
            I => n12470
        );

    \I__11671\ : CascadeMux
    port map (
            O => \N__51228\,
            I => \N__51224\
        );

    \I__11670\ : InMux
    port map (
            O => \N__51227\,
            I => \N__51221\
        );

    \I__11669\ : InMux
    port map (
            O => \N__51224\,
            I => \N__51217\
        );

    \I__11668\ : LocalMux
    port map (
            O => \N__51221\,
            I => \N__51213\
        );

    \I__11667\ : InMux
    port map (
            O => \N__51220\,
            I => \N__51210\
        );

    \I__11666\ : LocalMux
    port map (
            O => \N__51217\,
            I => \N__51207\
        );

    \I__11665\ : InMux
    port map (
            O => \N__51216\,
            I => \N__51204\
        );

    \I__11664\ : Span4Mux_h
    port map (
            O => \N__51213\,
            I => \N__51201\
        );

    \I__11663\ : LocalMux
    port map (
            O => \N__51210\,
            I => encoder0_position_target_22
        );

    \I__11662\ : Odrv4
    port map (
            O => \N__51207\,
            I => encoder0_position_target_22
        );

    \I__11661\ : LocalMux
    port map (
            O => \N__51204\,
            I => encoder0_position_target_22
        );

    \I__11660\ : Odrv4
    port map (
            O => \N__51201\,
            I => encoder0_position_target_22
        );

    \I__11659\ : InMux
    port map (
            O => \N__51192\,
            I => n12471
        );

    \I__11658\ : CascadeMux
    port map (
            O => \N__51189\,
            I => \N__51182\
        );

    \I__11657\ : CascadeMux
    port map (
            O => \N__51188\,
            I => \N__51178\
        );

    \I__11656\ : CascadeMux
    port map (
            O => \N__51187\,
            I => \N__51174\
        );

    \I__11655\ : CascadeMux
    port map (
            O => \N__51186\,
            I => \N__51170\
        );

    \I__11654\ : InMux
    port map (
            O => \N__51185\,
            I => \N__51161\
        );

    \I__11653\ : InMux
    port map (
            O => \N__51182\,
            I => \N__51144\
        );

    \I__11652\ : InMux
    port map (
            O => \N__51181\,
            I => \N__51144\
        );

    \I__11651\ : InMux
    port map (
            O => \N__51178\,
            I => \N__51144\
        );

    \I__11650\ : InMux
    port map (
            O => \N__51177\,
            I => \N__51144\
        );

    \I__11649\ : InMux
    port map (
            O => \N__51174\,
            I => \N__51144\
        );

    \I__11648\ : InMux
    port map (
            O => \N__51173\,
            I => \N__51144\
        );

    \I__11647\ : InMux
    port map (
            O => \N__51170\,
            I => \N__51144\
        );

    \I__11646\ : InMux
    port map (
            O => \N__51169\,
            I => \N__51144\
        );

    \I__11645\ : CascadeMux
    port map (
            O => \N__51168\,
            I => \N__51140\
        );

    \I__11644\ : CascadeMux
    port map (
            O => \N__51167\,
            I => \N__51136\
        );

    \I__11643\ : CascadeMux
    port map (
            O => \N__51166\,
            I => \N__51132\
        );

    \I__11642\ : CascadeMux
    port map (
            O => \N__51165\,
            I => \N__51128\
        );

    \I__11641\ : CascadeMux
    port map (
            O => \N__51164\,
            I => \N__51122\
        );

    \I__11640\ : LocalMux
    port map (
            O => \N__51161\,
            I => \N__51110\
        );

    \I__11639\ : LocalMux
    port map (
            O => \N__51144\,
            I => \N__51110\
        );

    \I__11638\ : InMux
    port map (
            O => \N__51143\,
            I => \N__51093\
        );

    \I__11637\ : InMux
    port map (
            O => \N__51140\,
            I => \N__51093\
        );

    \I__11636\ : InMux
    port map (
            O => \N__51139\,
            I => \N__51093\
        );

    \I__11635\ : InMux
    port map (
            O => \N__51136\,
            I => \N__51093\
        );

    \I__11634\ : InMux
    port map (
            O => \N__51135\,
            I => \N__51093\
        );

    \I__11633\ : InMux
    port map (
            O => \N__51132\,
            I => \N__51093\
        );

    \I__11632\ : InMux
    port map (
            O => \N__51131\,
            I => \N__51093\
        );

    \I__11631\ : InMux
    port map (
            O => \N__51128\,
            I => \N__51093\
        );

    \I__11630\ : InMux
    port map (
            O => \N__51127\,
            I => \N__51084\
        );

    \I__11629\ : InMux
    port map (
            O => \N__51126\,
            I => \N__51084\
        );

    \I__11628\ : InMux
    port map (
            O => \N__51125\,
            I => \N__51084\
        );

    \I__11627\ : InMux
    port map (
            O => \N__51122\,
            I => \N__51084\
        );

    \I__11626\ : InMux
    port map (
            O => \N__51121\,
            I => \N__51075\
        );

    \I__11625\ : InMux
    port map (
            O => \N__51120\,
            I => \N__51075\
        );

    \I__11624\ : InMux
    port map (
            O => \N__51119\,
            I => \N__51075\
        );

    \I__11623\ : InMux
    port map (
            O => \N__51118\,
            I => \N__51075\
        );

    \I__11622\ : InMux
    port map (
            O => \N__51117\,
            I => \N__51068\
        );

    \I__11621\ : InMux
    port map (
            O => \N__51116\,
            I => \N__51068\
        );

    \I__11620\ : InMux
    port map (
            O => \N__51115\,
            I => \N__51068\
        );

    \I__11619\ : Odrv4
    port map (
            O => \N__51110\,
            I => direction_c
        );

    \I__11618\ : LocalMux
    port map (
            O => \N__51093\,
            I => direction_c
        );

    \I__11617\ : LocalMux
    port map (
            O => \N__51084\,
            I => direction_c
        );

    \I__11616\ : LocalMux
    port map (
            O => \N__51075\,
            I => direction_c
        );

    \I__11615\ : LocalMux
    port map (
            O => \N__51068\,
            I => direction_c
        );

    \I__11614\ : InMux
    port map (
            O => \N__51057\,
            I => \bfn_15_28_0_\
        );

    \I__11613\ : InMux
    port map (
            O => \N__51054\,
            I => \N__51051\
        );

    \I__11612\ : LocalMux
    port map (
            O => \N__51051\,
            I => \N__51046\
        );

    \I__11611\ : InMux
    port map (
            O => \N__51050\,
            I => \N__51043\
        );

    \I__11610\ : CascadeMux
    port map (
            O => \N__51049\,
            I => \N__51040\
        );

    \I__11609\ : Span4Mux_v
    port map (
            O => \N__51046\,
            I => \N__51034\
        );

    \I__11608\ : LocalMux
    port map (
            O => \N__51043\,
            I => \N__51031\
        );

    \I__11607\ : InMux
    port map (
            O => \N__51040\,
            I => \N__51028\
        );

    \I__11606\ : InMux
    port map (
            O => \N__51039\,
            I => \N__51025\
        );

    \I__11605\ : InMux
    port map (
            O => \N__51038\,
            I => \N__51022\
        );

    \I__11604\ : InMux
    port map (
            O => \N__51037\,
            I => \N__51019\
        );

    \I__11603\ : Span4Mux_h
    port map (
            O => \N__51034\,
            I => \N__51016\
        );

    \I__11602\ : Span4Mux_h
    port map (
            O => \N__51031\,
            I => \N__51013\
        );

    \I__11601\ : LocalMux
    port map (
            O => \N__51028\,
            I => \N__51006\
        );

    \I__11600\ : LocalMux
    port map (
            O => \N__51025\,
            I => \N__51006\
        );

    \I__11599\ : LocalMux
    port map (
            O => \N__51022\,
            I => \N__51006\
        );

    \I__11598\ : LocalMux
    port map (
            O => \N__51019\,
            I => encoder0_position_target_23
        );

    \I__11597\ : Odrv4
    port map (
            O => \N__51016\,
            I => encoder0_position_target_23
        );

    \I__11596\ : Odrv4
    port map (
            O => \N__51013\,
            I => encoder0_position_target_23
        );

    \I__11595\ : Odrv4
    port map (
            O => \N__51006\,
            I => encoder0_position_target_23
        );

    \I__11594\ : InMux
    port map (
            O => \N__50997\,
            I => \N__50994\
        );

    \I__11593\ : LocalMux
    port map (
            O => \N__50994\,
            I => \N__50991\
        );

    \I__11592\ : Span4Mux_h
    port map (
            O => \N__50991\,
            I => \N__50988\
        );

    \I__11591\ : Span4Mux_h
    port map (
            O => \N__50988\,
            I => \N__50985\
        );

    \I__11590\ : Odrv4
    port map (
            O => \N__50985\,
            I => pwm_setpoint_23
        );

    \I__11589\ : InMux
    port map (
            O => \N__50982\,
            I => \N__50977\
        );

    \I__11588\ : InMux
    port map (
            O => \N__50981\,
            I => \N__50974\
        );

    \I__11587\ : InMux
    port map (
            O => \N__50980\,
            I => \N__50971\
        );

    \I__11586\ : LocalMux
    port map (
            O => \N__50977\,
            I => pwm_counter_23
        );

    \I__11585\ : LocalMux
    port map (
            O => \N__50974\,
            I => pwm_counter_23
        );

    \I__11584\ : LocalMux
    port map (
            O => \N__50971\,
            I => pwm_counter_23
        );

    \I__11583\ : InMux
    port map (
            O => \N__50964\,
            I => \N__50961\
        );

    \I__11582\ : LocalMux
    port map (
            O => \N__50961\,
            I => \N__50958\
        );

    \I__11581\ : Span4Mux_h
    port map (
            O => \N__50958\,
            I => \N__50955\
        );

    \I__11580\ : Odrv4
    port map (
            O => \N__50955\,
            I => n15245
        );

    \I__11579\ : InMux
    port map (
            O => \N__50952\,
            I => \N__50947\
        );

    \I__11578\ : InMux
    port map (
            O => \N__50951\,
            I => \N__50944\
        );

    \I__11577\ : InMux
    port map (
            O => \N__50950\,
            I => \N__50941\
        );

    \I__11576\ : LocalMux
    port map (
            O => \N__50947\,
            I => pwm_counter_31
        );

    \I__11575\ : LocalMux
    port map (
            O => \N__50944\,
            I => pwm_counter_31
        );

    \I__11574\ : LocalMux
    port map (
            O => \N__50941\,
            I => pwm_counter_31
        );

    \I__11573\ : InMux
    port map (
            O => \N__50934\,
            I => \N__50930\
        );

    \I__11572\ : InMux
    port map (
            O => \N__50933\,
            I => \N__50927\
        );

    \I__11571\ : LocalMux
    port map (
            O => \N__50930\,
            I => \N__50924\
        );

    \I__11570\ : LocalMux
    port map (
            O => \N__50927\,
            I => n5180
        );

    \I__11569\ : Odrv4
    port map (
            O => \N__50924\,
            I => n5180
        );

    \I__11568\ : SRMux
    port map (
            O => \N__50919\,
            I => \N__50916\
        );

    \I__11567\ : LocalMux
    port map (
            O => \N__50916\,
            I => \N__50913\
        );

    \I__11566\ : Odrv12
    port map (
            O => \N__50913\,
            I => n5182
        );

    \I__11565\ : InMux
    port map (
            O => \N__50910\,
            I => \N__50902\
        );

    \I__11564\ : InMux
    port map (
            O => \N__50909\,
            I => \N__50896\
        );

    \I__11563\ : InMux
    port map (
            O => \N__50908\,
            I => \N__50885\
        );

    \I__11562\ : InMux
    port map (
            O => \N__50907\,
            I => \N__50885\
        );

    \I__11561\ : InMux
    port map (
            O => \N__50906\,
            I => \N__50885\
        );

    \I__11560\ : InMux
    port map (
            O => \N__50905\,
            I => \N__50882\
        );

    \I__11559\ : LocalMux
    port map (
            O => \N__50902\,
            I => \N__50879\
        );

    \I__11558\ : InMux
    port map (
            O => \N__50901\,
            I => \N__50874\
        );

    \I__11557\ : InMux
    port map (
            O => \N__50900\,
            I => \N__50874\
        );

    \I__11556\ : InMux
    port map (
            O => \N__50899\,
            I => \N__50870\
        );

    \I__11555\ : LocalMux
    port map (
            O => \N__50896\,
            I => \N__50864\
        );

    \I__11554\ : InMux
    port map (
            O => \N__50895\,
            I => \N__50858\
        );

    \I__11553\ : InMux
    port map (
            O => \N__50894\,
            I => \N__50858\
        );

    \I__11552\ : InMux
    port map (
            O => \N__50893\,
            I => \N__50853\
        );

    \I__11551\ : InMux
    port map (
            O => \N__50892\,
            I => \N__50853\
        );

    \I__11550\ : LocalMux
    port map (
            O => \N__50885\,
            I => \N__50850\
        );

    \I__11549\ : LocalMux
    port map (
            O => \N__50882\,
            I => \N__50847\
        );

    \I__11548\ : Span4Mux_s1_v
    port map (
            O => \N__50879\,
            I => \N__50842\
        );

    \I__11547\ : LocalMux
    port map (
            O => \N__50874\,
            I => \N__50842\
        );

    \I__11546\ : InMux
    port map (
            O => \N__50873\,
            I => \N__50839\
        );

    \I__11545\ : LocalMux
    port map (
            O => \N__50870\,
            I => \N__50829\
        );

    \I__11544\ : InMux
    port map (
            O => \N__50869\,
            I => \N__50822\
        );

    \I__11543\ : InMux
    port map (
            O => \N__50868\,
            I => \N__50822\
        );

    \I__11542\ : InMux
    port map (
            O => \N__50867\,
            I => \N__50822\
        );

    \I__11541\ : Span4Mux_v
    port map (
            O => \N__50864\,
            I => \N__50819\
        );

    \I__11540\ : InMux
    port map (
            O => \N__50863\,
            I => \N__50816\
        );

    \I__11539\ : LocalMux
    port map (
            O => \N__50858\,
            I => \N__50811\
        );

    \I__11538\ : LocalMux
    port map (
            O => \N__50853\,
            I => \N__50811\
        );

    \I__11537\ : Span4Mux_v
    port map (
            O => \N__50850\,
            I => \N__50806\
        );

    \I__11536\ : Span4Mux_v
    port map (
            O => \N__50847\,
            I => \N__50806\
        );

    \I__11535\ : Sp12to4
    port map (
            O => \N__50842\,
            I => \N__50801\
        );

    \I__11534\ : LocalMux
    port map (
            O => \N__50839\,
            I => \N__50801\
        );

    \I__11533\ : InMux
    port map (
            O => \N__50838\,
            I => \N__50798\
        );

    \I__11532\ : InMux
    port map (
            O => \N__50837\,
            I => \N__50795\
        );

    \I__11531\ : InMux
    port map (
            O => \N__50836\,
            I => \N__50792\
        );

    \I__11530\ : InMux
    port map (
            O => \N__50835\,
            I => \N__50789\
        );

    \I__11529\ : InMux
    port map (
            O => \N__50834\,
            I => \N__50782\
        );

    \I__11528\ : InMux
    port map (
            O => \N__50833\,
            I => \N__50782\
        );

    \I__11527\ : InMux
    port map (
            O => \N__50832\,
            I => \N__50782\
        );

    \I__11526\ : Span12Mux_s5_v
    port map (
            O => \N__50829\,
            I => \N__50773\
        );

    \I__11525\ : LocalMux
    port map (
            O => \N__50822\,
            I => \N__50773\
        );

    \I__11524\ : Sp12to4
    port map (
            O => \N__50819\,
            I => \N__50773\
        );

    \I__11523\ : LocalMux
    port map (
            O => \N__50816\,
            I => \N__50773\
        );

    \I__11522\ : Odrv4
    port map (
            O => \N__50811\,
            I => duty_23
        );

    \I__11521\ : Odrv4
    port map (
            O => \N__50806\,
            I => duty_23
        );

    \I__11520\ : Odrv12
    port map (
            O => \N__50801\,
            I => duty_23
        );

    \I__11519\ : LocalMux
    port map (
            O => \N__50798\,
            I => duty_23
        );

    \I__11518\ : LocalMux
    port map (
            O => \N__50795\,
            I => duty_23
        );

    \I__11517\ : LocalMux
    port map (
            O => \N__50792\,
            I => duty_23
        );

    \I__11516\ : LocalMux
    port map (
            O => \N__50789\,
            I => duty_23
        );

    \I__11515\ : LocalMux
    port map (
            O => \N__50782\,
            I => duty_23
        );

    \I__11514\ : Odrv12
    port map (
            O => \N__50773\,
            I => duty_23
        );

    \I__11513\ : InMux
    port map (
            O => \N__50754\,
            I => \N__50751\
        );

    \I__11512\ : LocalMux
    port map (
            O => \N__50751\,
            I => \N__50747\
        );

    \I__11511\ : InMux
    port map (
            O => \N__50750\,
            I => \N__50744\
        );

    \I__11510\ : Span4Mux_h
    port map (
            O => \N__50747\,
            I => \N__50740\
        );

    \I__11509\ : LocalMux
    port map (
            O => \N__50744\,
            I => \N__50737\
        );

    \I__11508\ : InMux
    port map (
            O => \N__50743\,
            I => \N__50734\
        );

    \I__11507\ : Span4Mux_h
    port map (
            O => \N__50740\,
            I => \N__50731\
        );

    \I__11506\ : Span12Mux_h
    port map (
            O => \N__50737\,
            I => \N__50728\
        );

    \I__11505\ : LocalMux
    port map (
            O => \N__50734\,
            I => \N__50725\
        );

    \I__11504\ : Odrv4
    port map (
            O => \N__50731\,
            I => n300
        );

    \I__11503\ : Odrv12
    port map (
            O => \N__50728\,
            I => n300
        );

    \I__11502\ : Odrv12
    port map (
            O => \N__50725\,
            I => n300
        );

    \I__11501\ : InMux
    port map (
            O => \N__50718\,
            I => \N__50715\
        );

    \I__11500\ : LocalMux
    port map (
            O => \N__50715\,
            I => n1501
        );

    \I__11499\ : InMux
    port map (
            O => \N__50712\,
            I => \bfn_16_17_0_\
        );

    \I__11498\ : CascadeMux
    port map (
            O => \N__50709\,
            I => \N__50706\
        );

    \I__11497\ : InMux
    port map (
            O => \N__50706\,
            I => \N__50701\
        );

    \I__11496\ : CascadeMux
    port map (
            O => \N__50705\,
            I => \N__50697\
        );

    \I__11495\ : InMux
    port map (
            O => \N__50704\,
            I => \N__50694\
        );

    \I__11494\ : LocalMux
    port map (
            O => \N__50701\,
            I => \N__50691\
        );

    \I__11493\ : InMux
    port map (
            O => \N__50700\,
            I => \N__50686\
        );

    \I__11492\ : InMux
    port map (
            O => \N__50697\,
            I => \N__50686\
        );

    \I__11491\ : LocalMux
    port map (
            O => \N__50694\,
            I => encoder0_position_target_11
        );

    \I__11490\ : Odrv4
    port map (
            O => \N__50691\,
            I => encoder0_position_target_11
        );

    \I__11489\ : LocalMux
    port map (
            O => \N__50686\,
            I => encoder0_position_target_11
        );

    \I__11488\ : InMux
    port map (
            O => \N__50679\,
            I => n12460
        );

    \I__11487\ : CascadeMux
    port map (
            O => \N__50676\,
            I => \N__50671\
        );

    \I__11486\ : CascadeMux
    port map (
            O => \N__50675\,
            I => \N__50667\
        );

    \I__11485\ : InMux
    port map (
            O => \N__50674\,
            I => \N__50664\
        );

    \I__11484\ : InMux
    port map (
            O => \N__50671\,
            I => \N__50661\
        );

    \I__11483\ : InMux
    port map (
            O => \N__50670\,
            I => \N__50658\
        );

    \I__11482\ : InMux
    port map (
            O => \N__50667\,
            I => \N__50655\
        );

    \I__11481\ : LocalMux
    port map (
            O => \N__50664\,
            I => \N__50652\
        );

    \I__11480\ : LocalMux
    port map (
            O => \N__50661\,
            I => \N__50647\
        );

    \I__11479\ : LocalMux
    port map (
            O => \N__50658\,
            I => \N__50647\
        );

    \I__11478\ : LocalMux
    port map (
            O => \N__50655\,
            I => encoder0_position_target_12
        );

    \I__11477\ : Odrv4
    port map (
            O => \N__50652\,
            I => encoder0_position_target_12
        );

    \I__11476\ : Odrv4
    port map (
            O => \N__50647\,
            I => encoder0_position_target_12
        );

    \I__11475\ : InMux
    port map (
            O => \N__50640\,
            I => n12461
        );

    \I__11474\ : CascadeMux
    port map (
            O => \N__50637\,
            I => \N__50634\
        );

    \I__11473\ : InMux
    port map (
            O => \N__50634\,
            I => \N__50631\
        );

    \I__11472\ : LocalMux
    port map (
            O => \N__50631\,
            I => \N__50626\
        );

    \I__11471\ : InMux
    port map (
            O => \N__50630\,
            I => \N__50622\
        );

    \I__11470\ : InMux
    port map (
            O => \N__50629\,
            I => \N__50619\
        );

    \I__11469\ : Span4Mux_h
    port map (
            O => \N__50626\,
            I => \N__50616\
        );

    \I__11468\ : InMux
    port map (
            O => \N__50625\,
            I => \N__50613\
        );

    \I__11467\ : LocalMux
    port map (
            O => \N__50622\,
            I => \N__50610\
        );

    \I__11466\ : LocalMux
    port map (
            O => \N__50619\,
            I => encoder0_position_target_13
        );

    \I__11465\ : Odrv4
    port map (
            O => \N__50616\,
            I => encoder0_position_target_13
        );

    \I__11464\ : LocalMux
    port map (
            O => \N__50613\,
            I => encoder0_position_target_13
        );

    \I__11463\ : Odrv12
    port map (
            O => \N__50610\,
            I => encoder0_position_target_13
        );

    \I__11462\ : InMux
    port map (
            O => \N__50601\,
            I => n12462
        );

    \I__11461\ : CascadeMux
    port map (
            O => \N__50598\,
            I => \N__50594\
        );

    \I__11460\ : CascadeMux
    port map (
            O => \N__50597\,
            I => \N__50591\
        );

    \I__11459\ : InMux
    port map (
            O => \N__50594\,
            I => \N__50588\
        );

    \I__11458\ : InMux
    port map (
            O => \N__50591\,
            I => \N__50583\
        );

    \I__11457\ : LocalMux
    port map (
            O => \N__50588\,
            I => \N__50580\
        );

    \I__11456\ : InMux
    port map (
            O => \N__50587\,
            I => \N__50575\
        );

    \I__11455\ : InMux
    port map (
            O => \N__50586\,
            I => \N__50575\
        );

    \I__11454\ : LocalMux
    port map (
            O => \N__50583\,
            I => encoder0_position_target_14
        );

    \I__11453\ : Odrv12
    port map (
            O => \N__50580\,
            I => encoder0_position_target_14
        );

    \I__11452\ : LocalMux
    port map (
            O => \N__50575\,
            I => encoder0_position_target_14
        );

    \I__11451\ : InMux
    port map (
            O => \N__50568\,
            I => n12463
        );

    \I__11450\ : CascadeMux
    port map (
            O => \N__50565\,
            I => \N__50562\
        );

    \I__11449\ : InMux
    port map (
            O => \N__50562\,
            I => \N__50559\
        );

    \I__11448\ : LocalMux
    port map (
            O => \N__50559\,
            I => \N__50554\
        );

    \I__11447\ : CascadeMux
    port map (
            O => \N__50558\,
            I => \N__50551\
        );

    \I__11446\ : InMux
    port map (
            O => \N__50557\,
            I => \N__50548\
        );

    \I__11445\ : Span4Mux_v
    port map (
            O => \N__50554\,
            I => \N__50545\
        );

    \I__11444\ : InMux
    port map (
            O => \N__50551\,
            I => \N__50541\
        );

    \I__11443\ : LocalMux
    port map (
            O => \N__50548\,
            I => \N__50538\
        );

    \I__11442\ : Span4Mux_h
    port map (
            O => \N__50545\,
            I => \N__50535\
        );

    \I__11441\ : InMux
    port map (
            O => \N__50544\,
            I => \N__50532\
        );

    \I__11440\ : LocalMux
    port map (
            O => \N__50541\,
            I => \N__50527\
        );

    \I__11439\ : Span4Mux_v
    port map (
            O => \N__50538\,
            I => \N__50527\
        );

    \I__11438\ : Odrv4
    port map (
            O => \N__50535\,
            I => encoder0_position_target_15
        );

    \I__11437\ : LocalMux
    port map (
            O => \N__50532\,
            I => encoder0_position_target_15
        );

    \I__11436\ : Odrv4
    port map (
            O => \N__50527\,
            I => encoder0_position_target_15
        );

    \I__11435\ : InMux
    port map (
            O => \N__50520\,
            I => \bfn_15_27_0_\
        );

    \I__11434\ : CascadeMux
    port map (
            O => \N__50517\,
            I => \N__50514\
        );

    \I__11433\ : InMux
    port map (
            O => \N__50514\,
            I => \N__50511\
        );

    \I__11432\ : LocalMux
    port map (
            O => \N__50511\,
            I => \N__50506\
        );

    \I__11431\ : CascadeMux
    port map (
            O => \N__50510\,
            I => \N__50502\
        );

    \I__11430\ : InMux
    port map (
            O => \N__50509\,
            I => \N__50499\
        );

    \I__11429\ : Span4Mux_h
    port map (
            O => \N__50506\,
            I => \N__50496\
        );

    \I__11428\ : InMux
    port map (
            O => \N__50505\,
            I => \N__50491\
        );

    \I__11427\ : InMux
    port map (
            O => \N__50502\,
            I => \N__50491\
        );

    \I__11426\ : LocalMux
    port map (
            O => \N__50499\,
            I => encoder0_position_target_16
        );

    \I__11425\ : Odrv4
    port map (
            O => \N__50496\,
            I => encoder0_position_target_16
        );

    \I__11424\ : LocalMux
    port map (
            O => \N__50491\,
            I => encoder0_position_target_16
        );

    \I__11423\ : InMux
    port map (
            O => \N__50484\,
            I => n12465
        );

    \I__11422\ : CascadeMux
    port map (
            O => \N__50481\,
            I => \N__50478\
        );

    \I__11421\ : InMux
    port map (
            O => \N__50478\,
            I => \N__50473\
        );

    \I__11420\ : CascadeMux
    port map (
            O => \N__50477\,
            I => \N__50470\
        );

    \I__11419\ : InMux
    port map (
            O => \N__50476\,
            I => \N__50467\
        );

    \I__11418\ : LocalMux
    port map (
            O => \N__50473\,
            I => \N__50464\
        );

    \I__11417\ : InMux
    port map (
            O => \N__50470\,
            I => \N__50460\
        );

    \I__11416\ : LocalMux
    port map (
            O => \N__50467\,
            I => \N__50457\
        );

    \I__11415\ : Span4Mux_h
    port map (
            O => \N__50464\,
            I => \N__50454\
        );

    \I__11414\ : InMux
    port map (
            O => \N__50463\,
            I => \N__50451\
        );

    \I__11413\ : LocalMux
    port map (
            O => \N__50460\,
            I => \N__50446\
        );

    \I__11412\ : Span4Mux_v
    port map (
            O => \N__50457\,
            I => \N__50446\
        );

    \I__11411\ : Odrv4
    port map (
            O => \N__50454\,
            I => encoder0_position_target_17
        );

    \I__11410\ : LocalMux
    port map (
            O => \N__50451\,
            I => encoder0_position_target_17
        );

    \I__11409\ : Odrv4
    port map (
            O => \N__50446\,
            I => encoder0_position_target_17
        );

    \I__11408\ : InMux
    port map (
            O => \N__50439\,
            I => n12466
        );

    \I__11407\ : CascadeMux
    port map (
            O => \N__50436\,
            I => \N__50433\
        );

    \I__11406\ : InMux
    port map (
            O => \N__50433\,
            I => \N__50430\
        );

    \I__11405\ : LocalMux
    port map (
            O => \N__50430\,
            I => \N__50426\
        );

    \I__11404\ : InMux
    port map (
            O => \N__50429\,
            I => \N__50423\
        );

    \I__11403\ : Span4Mux_h
    port map (
            O => \N__50426\,
            I => \N__50420\
        );

    \I__11402\ : LocalMux
    port map (
            O => \N__50423\,
            I => \N__50413\
        );

    \I__11401\ : Span4Mux_v
    port map (
            O => \N__50420\,
            I => \N__50413\
        );

    \I__11400\ : InMux
    port map (
            O => \N__50419\,
            I => \N__50410\
        );

    \I__11399\ : InMux
    port map (
            O => \N__50418\,
            I => \N__50407\
        );

    \I__11398\ : Odrv4
    port map (
            O => \N__50413\,
            I => encoder0_position_target_18
        );

    \I__11397\ : LocalMux
    port map (
            O => \N__50410\,
            I => encoder0_position_target_18
        );

    \I__11396\ : LocalMux
    port map (
            O => \N__50407\,
            I => encoder0_position_target_18
        );

    \I__11395\ : InMux
    port map (
            O => \N__50400\,
            I => n12467
        );

    \I__11394\ : CascadeMux
    port map (
            O => \N__50397\,
            I => \N__50393\
        );

    \I__11393\ : CascadeMux
    port map (
            O => \N__50396\,
            I => \N__50388\
        );

    \I__11392\ : InMux
    port map (
            O => \N__50393\,
            I => \N__50385\
        );

    \I__11391\ : InMux
    port map (
            O => \N__50392\,
            I => \N__50382\
        );

    \I__11390\ : CascadeMux
    port map (
            O => \N__50391\,
            I => \N__50379\
        );

    \I__11389\ : InMux
    port map (
            O => \N__50388\,
            I => \N__50376\
        );

    \I__11388\ : LocalMux
    port map (
            O => \N__50385\,
            I => \N__50371\
        );

    \I__11387\ : LocalMux
    port map (
            O => \N__50382\,
            I => \N__50371\
        );

    \I__11386\ : InMux
    port map (
            O => \N__50379\,
            I => \N__50368\
        );

    \I__11385\ : LocalMux
    port map (
            O => \N__50376\,
            I => \N__50365\
        );

    \I__11384\ : Span4Mux_h
    port map (
            O => \N__50371\,
            I => \N__50362\
        );

    \I__11383\ : LocalMux
    port map (
            O => \N__50368\,
            I => encoder0_position_target_19
        );

    \I__11382\ : Odrv4
    port map (
            O => \N__50365\,
            I => encoder0_position_target_19
        );

    \I__11381\ : Odrv4
    port map (
            O => \N__50362\,
            I => encoder0_position_target_19
        );

    \I__11380\ : InMux
    port map (
            O => \N__50355\,
            I => n12468
        );

    \I__11379\ : CascadeMux
    port map (
            O => \N__50352\,
            I => \N__50348\
        );

    \I__11378\ : CascadeMux
    port map (
            O => \N__50351\,
            I => \N__50344\
        );

    \I__11377\ : InMux
    port map (
            O => \N__50348\,
            I => \N__50341\
        );

    \I__11376\ : InMux
    port map (
            O => \N__50347\,
            I => \N__50338\
        );

    \I__11375\ : InMux
    port map (
            O => \N__50344\,
            I => \N__50335\
        );

    \I__11374\ : LocalMux
    port map (
            O => \N__50341\,
            I => \N__50332\
        );

    \I__11373\ : LocalMux
    port map (
            O => \N__50338\,
            I => \N__50329\
        );

    \I__11372\ : LocalMux
    port map (
            O => \N__50335\,
            I => encoder0_position_target_3
        );

    \I__11371\ : Odrv4
    port map (
            O => \N__50332\,
            I => encoder0_position_target_3
        );

    \I__11370\ : Odrv4
    port map (
            O => \N__50329\,
            I => encoder0_position_target_3
        );

    \I__11369\ : InMux
    port map (
            O => \N__50322\,
            I => n12452
        );

    \I__11368\ : CascadeMux
    port map (
            O => \N__50319\,
            I => \N__50314\
        );

    \I__11367\ : InMux
    port map (
            O => \N__50318\,
            I => \N__50311\
        );

    \I__11366\ : CascadeMux
    port map (
            O => \N__50317\,
            I => \N__50307\
        );

    \I__11365\ : InMux
    port map (
            O => \N__50314\,
            I => \N__50304\
        );

    \I__11364\ : LocalMux
    port map (
            O => \N__50311\,
            I => \N__50301\
        );

    \I__11363\ : InMux
    port map (
            O => \N__50310\,
            I => \N__50298\
        );

    \I__11362\ : InMux
    port map (
            O => \N__50307\,
            I => \N__50295\
        );

    \I__11361\ : LocalMux
    port map (
            O => \N__50304\,
            I => \N__50292\
        );

    \I__11360\ : Span4Mux_h
    port map (
            O => \N__50301\,
            I => \N__50289\
        );

    \I__11359\ : LocalMux
    port map (
            O => \N__50298\,
            I => \N__50286\
        );

    \I__11358\ : LocalMux
    port map (
            O => \N__50295\,
            I => encoder0_position_target_4
        );

    \I__11357\ : Odrv12
    port map (
            O => \N__50292\,
            I => encoder0_position_target_4
        );

    \I__11356\ : Odrv4
    port map (
            O => \N__50289\,
            I => encoder0_position_target_4
        );

    \I__11355\ : Odrv4
    port map (
            O => \N__50286\,
            I => encoder0_position_target_4
        );

    \I__11354\ : InMux
    port map (
            O => \N__50277\,
            I => n12453
        );

    \I__11353\ : CascadeMux
    port map (
            O => \N__50274\,
            I => \N__50271\
        );

    \I__11352\ : InMux
    port map (
            O => \N__50271\,
            I => \N__50267\
        );

    \I__11351\ : CascadeMux
    port map (
            O => \N__50270\,
            I => \N__50262\
        );

    \I__11350\ : LocalMux
    port map (
            O => \N__50267\,
            I => \N__50259\
        );

    \I__11349\ : InMux
    port map (
            O => \N__50266\,
            I => \N__50254\
        );

    \I__11348\ : InMux
    port map (
            O => \N__50265\,
            I => \N__50254\
        );

    \I__11347\ : InMux
    port map (
            O => \N__50262\,
            I => \N__50251\
        );

    \I__11346\ : Span4Mux_h
    port map (
            O => \N__50259\,
            I => \N__50246\
        );

    \I__11345\ : LocalMux
    port map (
            O => \N__50254\,
            I => \N__50246\
        );

    \I__11344\ : LocalMux
    port map (
            O => \N__50251\,
            I => encoder0_position_target_5
        );

    \I__11343\ : Odrv4
    port map (
            O => \N__50246\,
            I => encoder0_position_target_5
        );

    \I__11342\ : InMux
    port map (
            O => \N__50241\,
            I => n12454
        );

    \I__11341\ : CascadeMux
    port map (
            O => \N__50238\,
            I => \N__50234\
        );

    \I__11340\ : CascadeMux
    port map (
            O => \N__50237\,
            I => \N__50229\
        );

    \I__11339\ : InMux
    port map (
            O => \N__50234\,
            I => \N__50226\
        );

    \I__11338\ : InMux
    port map (
            O => \N__50233\,
            I => \N__50221\
        );

    \I__11337\ : InMux
    port map (
            O => \N__50232\,
            I => \N__50221\
        );

    \I__11336\ : InMux
    port map (
            O => \N__50229\,
            I => \N__50218\
        );

    \I__11335\ : LocalMux
    port map (
            O => \N__50226\,
            I => \N__50215\
        );

    \I__11334\ : LocalMux
    port map (
            O => \N__50221\,
            I => \N__50212\
        );

    \I__11333\ : LocalMux
    port map (
            O => \N__50218\,
            I => encoder0_position_target_6
        );

    \I__11332\ : Odrv4
    port map (
            O => \N__50215\,
            I => encoder0_position_target_6
        );

    \I__11331\ : Odrv4
    port map (
            O => \N__50212\,
            I => encoder0_position_target_6
        );

    \I__11330\ : InMux
    port map (
            O => \N__50205\,
            I => n12455
        );

    \I__11329\ : CascadeMux
    port map (
            O => \N__50202\,
            I => \N__50199\
        );

    \I__11328\ : InMux
    port map (
            O => \N__50199\,
            I => \N__50195\
        );

    \I__11327\ : CascadeMux
    port map (
            O => \N__50198\,
            I => \N__50192\
        );

    \I__11326\ : LocalMux
    port map (
            O => \N__50195\,
            I => \N__50188\
        );

    \I__11325\ : InMux
    port map (
            O => \N__50192\,
            I => \N__50185\
        );

    \I__11324\ : InMux
    port map (
            O => \N__50191\,
            I => \N__50182\
        );

    \I__11323\ : Span4Mux_v
    port map (
            O => \N__50188\,
            I => \N__50178\
        );

    \I__11322\ : LocalMux
    port map (
            O => \N__50185\,
            I => \N__50173\
        );

    \I__11321\ : LocalMux
    port map (
            O => \N__50182\,
            I => \N__50173\
        );

    \I__11320\ : InMux
    port map (
            O => \N__50181\,
            I => \N__50170\
        );

    \I__11319\ : Span4Mux_v
    port map (
            O => \N__50178\,
            I => \N__50165\
        );

    \I__11318\ : Span4Mux_v
    port map (
            O => \N__50173\,
            I => \N__50165\
        );

    \I__11317\ : LocalMux
    port map (
            O => \N__50170\,
            I => encoder0_position_target_7
        );

    \I__11316\ : Odrv4
    port map (
            O => \N__50165\,
            I => encoder0_position_target_7
        );

    \I__11315\ : InMux
    port map (
            O => \N__50160\,
            I => \bfn_15_26_0_\
        );

    \I__11314\ : CascadeMux
    port map (
            O => \N__50157\,
            I => \N__50154\
        );

    \I__11313\ : InMux
    port map (
            O => \N__50154\,
            I => \N__50148\
        );

    \I__11312\ : InMux
    port map (
            O => \N__50153\,
            I => \N__50145\
        );

    \I__11311\ : CascadeMux
    port map (
            O => \N__50152\,
            I => \N__50142\
        );

    \I__11310\ : InMux
    port map (
            O => \N__50151\,
            I => \N__50139\
        );

    \I__11309\ : LocalMux
    port map (
            O => \N__50148\,
            I => \N__50134\
        );

    \I__11308\ : LocalMux
    port map (
            O => \N__50145\,
            I => \N__50134\
        );

    \I__11307\ : InMux
    port map (
            O => \N__50142\,
            I => \N__50131\
        );

    \I__11306\ : LocalMux
    port map (
            O => \N__50139\,
            I => \N__50126\
        );

    \I__11305\ : Span4Mux_v
    port map (
            O => \N__50134\,
            I => \N__50126\
        );

    \I__11304\ : LocalMux
    port map (
            O => \N__50131\,
            I => encoder0_position_target_8
        );

    \I__11303\ : Odrv4
    port map (
            O => \N__50126\,
            I => encoder0_position_target_8
        );

    \I__11302\ : InMux
    port map (
            O => \N__50121\,
            I => n12457
        );

    \I__11301\ : CascadeMux
    port map (
            O => \N__50118\,
            I => \N__50114\
        );

    \I__11300\ : InMux
    port map (
            O => \N__50117\,
            I => \N__50111\
        );

    \I__11299\ : InMux
    port map (
            O => \N__50114\,
            I => \N__50108\
        );

    \I__11298\ : LocalMux
    port map (
            O => \N__50111\,
            I => \N__50103\
        );

    \I__11297\ : LocalMux
    port map (
            O => \N__50108\,
            I => \N__50100\
        );

    \I__11296\ : InMux
    port map (
            O => \N__50107\,
            I => \N__50097\
        );

    \I__11295\ : InMux
    port map (
            O => \N__50106\,
            I => \N__50094\
        );

    \I__11294\ : Span4Mux_h
    port map (
            O => \N__50103\,
            I => \N__50091\
        );

    \I__11293\ : Span4Mux_v
    port map (
            O => \N__50100\,
            I => \N__50086\
        );

    \I__11292\ : LocalMux
    port map (
            O => \N__50097\,
            I => \N__50086\
        );

    \I__11291\ : LocalMux
    port map (
            O => \N__50094\,
            I => encoder0_position_target_9
        );

    \I__11290\ : Odrv4
    port map (
            O => \N__50091\,
            I => encoder0_position_target_9
        );

    \I__11289\ : Odrv4
    port map (
            O => \N__50086\,
            I => encoder0_position_target_9
        );

    \I__11288\ : InMux
    port map (
            O => \N__50079\,
            I => n12458
        );

    \I__11287\ : CascadeMux
    port map (
            O => \N__50076\,
            I => \N__50073\
        );

    \I__11286\ : InMux
    port map (
            O => \N__50073\,
            I => \N__50067\
        );

    \I__11285\ : InMux
    port map (
            O => \N__50072\,
            I => \N__50062\
        );

    \I__11284\ : InMux
    port map (
            O => \N__50071\,
            I => \N__50062\
        );

    \I__11283\ : CascadeMux
    port map (
            O => \N__50070\,
            I => \N__50059\
        );

    \I__11282\ : LocalMux
    port map (
            O => \N__50067\,
            I => \N__50056\
        );

    \I__11281\ : LocalMux
    port map (
            O => \N__50062\,
            I => \N__50053\
        );

    \I__11280\ : InMux
    port map (
            O => \N__50059\,
            I => \N__50050\
        );

    \I__11279\ : Span4Mux_h
    port map (
            O => \N__50056\,
            I => \N__50047\
        );

    \I__11278\ : Span4Mux_h
    port map (
            O => \N__50053\,
            I => \N__50044\
        );

    \I__11277\ : LocalMux
    port map (
            O => \N__50050\,
            I => encoder0_position_target_10
        );

    \I__11276\ : Odrv4
    port map (
            O => \N__50047\,
            I => encoder0_position_target_10
        );

    \I__11275\ : Odrv4
    port map (
            O => \N__50044\,
            I => encoder0_position_target_10
        );

    \I__11274\ : InMux
    port map (
            O => \N__50037\,
            I => n12459
        );

    \I__11273\ : InMux
    port map (
            O => \N__50034\,
            I => \N__50030\
        );

    \I__11272\ : CascadeMux
    port map (
            O => \N__50033\,
            I => \N__50027\
        );

    \I__11271\ : LocalMux
    port map (
            O => \N__50030\,
            I => \N__50023\
        );

    \I__11270\ : InMux
    port map (
            O => \N__50027\,
            I => \N__50020\
        );

    \I__11269\ : InMux
    port map (
            O => \N__50026\,
            I => \N__50017\
        );

    \I__11268\ : Odrv12
    port map (
            O => \N__50023\,
            I => n1126
        );

    \I__11267\ : LocalMux
    port map (
            O => \N__50020\,
            I => n1126
        );

    \I__11266\ : LocalMux
    port map (
            O => \N__50017\,
            I => n1126
        );

    \I__11265\ : InMux
    port map (
            O => \N__50010\,
            I => \N__50007\
        );

    \I__11264\ : LocalMux
    port map (
            O => \N__50007\,
            I => n1193
        );

    \I__11263\ : CascadeMux
    port map (
            O => \N__50004\,
            I => \n1225_cascade_\
        );

    \I__11262\ : InMux
    port map (
            O => \N__50001\,
            I => \N__49996\
        );

    \I__11261\ : InMux
    port map (
            O => \N__50000\,
            I => \N__49991\
        );

    \I__11260\ : InMux
    port map (
            O => \N__49999\,
            I => \N__49991\
        );

    \I__11259\ : LocalMux
    port map (
            O => \N__49996\,
            I => \N__49986\
        );

    \I__11258\ : LocalMux
    port map (
            O => \N__49991\,
            I => \N__49986\
        );

    \I__11257\ : Odrv4
    port map (
            O => \N__49986\,
            I => n1324
        );

    \I__11256\ : InMux
    port map (
            O => \N__49983\,
            I => \N__49980\
        );

    \I__11255\ : LocalMux
    port map (
            O => \N__49980\,
            I => \N__49976\
        );

    \I__11254\ : CascadeMux
    port map (
            O => \N__49979\,
            I => \N__49973\
        );

    \I__11253\ : Span4Mux_v
    port map (
            O => \N__49976\,
            I => \N__49970\
        );

    \I__11252\ : InMux
    port map (
            O => \N__49973\,
            I => \N__49967\
        );

    \I__11251\ : Odrv4
    port map (
            O => \N__49970\,
            I => n1129
        );

    \I__11250\ : LocalMux
    port map (
            O => \N__49967\,
            I => n1129
        );

    \I__11249\ : CascadeMux
    port map (
            O => \N__49962\,
            I => \N__49959\
        );

    \I__11248\ : InMux
    port map (
            O => \N__49959\,
            I => \N__49956\
        );

    \I__11247\ : LocalMux
    port map (
            O => \N__49956\,
            I => n1196
        );

    \I__11246\ : InMux
    port map (
            O => \N__49953\,
            I => \N__49950\
        );

    \I__11245\ : LocalMux
    port map (
            O => \N__49950\,
            I => \N__49947\
        );

    \I__11244\ : Span4Mux_h
    port map (
            O => \N__49947\,
            I => \N__49944\
        );

    \I__11243\ : Span4Mux_h
    port map (
            O => \N__49944\,
            I => \N__49938\
        );

    \I__11242\ : CascadeMux
    port map (
            O => \N__49943\,
            I => \N__49935\
        );

    \I__11241\ : CascadeMux
    port map (
            O => \N__49942\,
            I => \N__49931\
        );

    \I__11240\ : InMux
    port map (
            O => \N__49941\,
            I => \N__49925\
        );

    \I__11239\ : Span4Mux_v
    port map (
            O => \N__49938\,
            I => \N__49919\
        );

    \I__11238\ : InMux
    port map (
            O => \N__49935\,
            I => \N__49916\
        );

    \I__11237\ : InMux
    port map (
            O => \N__49934\,
            I => \N__49913\
        );

    \I__11236\ : InMux
    port map (
            O => \N__49931\,
            I => \N__49904\
        );

    \I__11235\ : InMux
    port map (
            O => \N__49930\,
            I => \N__49904\
        );

    \I__11234\ : InMux
    port map (
            O => \N__49929\,
            I => \N__49904\
        );

    \I__11233\ : InMux
    port map (
            O => \N__49928\,
            I => \N__49904\
        );

    \I__11232\ : LocalMux
    port map (
            O => \N__49925\,
            I => \N__49901\
        );

    \I__11231\ : InMux
    port map (
            O => \N__49924\,
            I => \N__49894\
        );

    \I__11230\ : InMux
    port map (
            O => \N__49923\,
            I => \N__49894\
        );

    \I__11229\ : InMux
    port map (
            O => \N__49922\,
            I => \N__49894\
        );

    \I__11228\ : Odrv4
    port map (
            O => \N__49919\,
            I => n1158
        );

    \I__11227\ : LocalMux
    port map (
            O => \N__49916\,
            I => n1158
        );

    \I__11226\ : LocalMux
    port map (
            O => \N__49913\,
            I => n1158
        );

    \I__11225\ : LocalMux
    port map (
            O => \N__49904\,
            I => n1158
        );

    \I__11224\ : Odrv4
    port map (
            O => \N__49901\,
            I => n1158
        );

    \I__11223\ : LocalMux
    port map (
            O => \N__49894\,
            I => n1158
        );

    \I__11222\ : InMux
    port map (
            O => \N__49881\,
            I => \N__49878\
        );

    \I__11221\ : LocalMux
    port map (
            O => \N__49878\,
            I => \N__49872\
        );

    \I__11220\ : InMux
    port map (
            O => \N__49877\,
            I => \N__49869\
        );

    \I__11219\ : CascadeMux
    port map (
            O => \N__49876\,
            I => \N__49864\
        );

    \I__11218\ : CascadeMux
    port map (
            O => \N__49875\,
            I => \N__49861\
        );

    \I__11217\ : Span4Mux_h
    port map (
            O => \N__49872\,
            I => \N__49855\
        );

    \I__11216\ : LocalMux
    port map (
            O => \N__49869\,
            I => \N__49855\
        );

    \I__11215\ : CascadeMux
    port map (
            O => \N__49868\,
            I => \N__49851\
        );

    \I__11214\ : CascadeMux
    port map (
            O => \N__49867\,
            I => \N__49848\
        );

    \I__11213\ : InMux
    port map (
            O => \N__49864\,
            I => \N__49843\
        );

    \I__11212\ : InMux
    port map (
            O => \N__49861\,
            I => \N__49843\
        );

    \I__11211\ : CascadeMux
    port map (
            O => \N__49860\,
            I => \N__49838\
        );

    \I__11210\ : Span4Mux_v
    port map (
            O => \N__49855\,
            I => \N__49835\
        );

    \I__11209\ : InMux
    port map (
            O => \N__49854\,
            I => \N__49832\
        );

    \I__11208\ : InMux
    port map (
            O => \N__49851\,
            I => \N__49827\
        );

    \I__11207\ : InMux
    port map (
            O => \N__49848\,
            I => \N__49827\
        );

    \I__11206\ : LocalMux
    port map (
            O => \N__49843\,
            I => \N__49824\
        );

    \I__11205\ : InMux
    port map (
            O => \N__49842\,
            I => \N__49817\
        );

    \I__11204\ : InMux
    port map (
            O => \N__49841\,
            I => \N__49817\
        );

    \I__11203\ : InMux
    port map (
            O => \N__49838\,
            I => \N__49817\
        );

    \I__11202\ : Odrv4
    port map (
            O => \N__49835\,
            I => n1059
        );

    \I__11201\ : LocalMux
    port map (
            O => \N__49832\,
            I => n1059
        );

    \I__11200\ : LocalMux
    port map (
            O => \N__49827\,
            I => n1059
        );

    \I__11199\ : Odrv4
    port map (
            O => \N__49824\,
            I => n1059
        );

    \I__11198\ : LocalMux
    port map (
            O => \N__49817\,
            I => n1059
        );

    \I__11197\ : InMux
    port map (
            O => \N__49806\,
            I => \N__49802\
        );

    \I__11196\ : CascadeMux
    port map (
            O => \N__49805\,
            I => \N__49798\
        );

    \I__11195\ : LocalMux
    port map (
            O => \N__49802\,
            I => \N__49795\
        );

    \I__11194\ : InMux
    port map (
            O => \N__49801\,
            I => \N__49792\
        );

    \I__11193\ : InMux
    port map (
            O => \N__49798\,
            I => \N__49789\
        );

    \I__11192\ : Odrv4
    port map (
            O => \N__49795\,
            I => n1128
        );

    \I__11191\ : LocalMux
    port map (
            O => \N__49792\,
            I => n1128
        );

    \I__11190\ : LocalMux
    port map (
            O => \N__49789\,
            I => n1128
        );

    \I__11189\ : CascadeMux
    port map (
            O => \N__49782\,
            I => \N__49779\
        );

    \I__11188\ : InMux
    port map (
            O => \N__49779\,
            I => \N__49776\
        );

    \I__11187\ : LocalMux
    port map (
            O => \N__49776\,
            I => \N__49773\
        );

    \I__11186\ : Odrv4
    port map (
            O => \N__49773\,
            I => n1693
        );

    \I__11185\ : CascadeMux
    port map (
            O => \N__49770\,
            I => \N__49767\
        );

    \I__11184\ : InMux
    port map (
            O => \N__49767\,
            I => \N__49764\
        );

    \I__11183\ : LocalMux
    port map (
            O => \N__49764\,
            I => \N__49759\
        );

    \I__11182\ : InMux
    port map (
            O => \N__49763\,
            I => \N__49756\
        );

    \I__11181\ : InMux
    port map (
            O => \N__49762\,
            I => \N__49753\
        );

    \I__11180\ : Span4Mux_h
    port map (
            O => \N__49759\,
            I => \N__49748\
        );

    \I__11179\ : LocalMux
    port map (
            O => \N__49756\,
            I => \N__49748\
        );

    \I__11178\ : LocalMux
    port map (
            O => \N__49753\,
            I => encoder0_position_target_0
        );

    \I__11177\ : Odrv4
    port map (
            O => \N__49748\,
            I => encoder0_position_target_0
        );

    \I__11176\ : InMux
    port map (
            O => \N__49743\,
            I => n12449
        );

    \I__11175\ : CascadeMux
    port map (
            O => \N__49740\,
            I => \N__49737\
        );

    \I__11174\ : InMux
    port map (
            O => \N__49737\,
            I => \N__49732\
        );

    \I__11173\ : CascadeMux
    port map (
            O => \N__49736\,
            I => \N__49729\
        );

    \I__11172\ : CascadeMux
    port map (
            O => \N__49735\,
            I => \N__49726\
        );

    \I__11171\ : LocalMux
    port map (
            O => \N__49732\,
            I => \N__49723\
        );

    \I__11170\ : InMux
    port map (
            O => \N__49729\,
            I => \N__49720\
        );

    \I__11169\ : InMux
    port map (
            O => \N__49726\,
            I => \N__49717\
        );

    \I__11168\ : Sp12to4
    port map (
            O => \N__49723\,
            I => \N__49712\
        );

    \I__11167\ : LocalMux
    port map (
            O => \N__49720\,
            I => \N__49712\
        );

    \I__11166\ : LocalMux
    port map (
            O => \N__49717\,
            I => encoder0_position_target_1
        );

    \I__11165\ : Odrv12
    port map (
            O => \N__49712\,
            I => encoder0_position_target_1
        );

    \I__11164\ : InMux
    port map (
            O => \N__49707\,
            I => n12450
        );

    \I__11163\ : CascadeMux
    port map (
            O => \N__49704\,
            I => \N__49700\
        );

    \I__11162\ : CascadeMux
    port map (
            O => \N__49703\,
            I => \N__49696\
        );

    \I__11161\ : InMux
    port map (
            O => \N__49700\,
            I => \N__49693\
        );

    \I__11160\ : InMux
    port map (
            O => \N__49699\,
            I => \N__49690\
        );

    \I__11159\ : InMux
    port map (
            O => \N__49696\,
            I => \N__49687\
        );

    \I__11158\ : LocalMux
    port map (
            O => \N__49693\,
            I => \N__49684\
        );

    \I__11157\ : LocalMux
    port map (
            O => \N__49690\,
            I => \N__49681\
        );

    \I__11156\ : LocalMux
    port map (
            O => \N__49687\,
            I => encoder0_position_target_2
        );

    \I__11155\ : Odrv12
    port map (
            O => \N__49684\,
            I => encoder0_position_target_2
        );

    \I__11154\ : Odrv4
    port map (
            O => \N__49681\,
            I => encoder0_position_target_2
        );

    \I__11153\ : InMux
    port map (
            O => \N__49674\,
            I => n12451
        );

    \I__11152\ : CascadeMux
    port map (
            O => \N__49671\,
            I => \n1257_cascade_\
        );

    \I__11151\ : CascadeMux
    port map (
            O => \N__49668\,
            I => \N__49665\
        );

    \I__11150\ : InMux
    port map (
            O => \N__49665\,
            I => \N__49661\
        );

    \I__11149\ : CascadeMux
    port map (
            O => \N__49664\,
            I => \N__49658\
        );

    \I__11148\ : LocalMux
    port map (
            O => \N__49661\,
            I => \N__49654\
        );

    \I__11147\ : InMux
    port map (
            O => \N__49658\,
            I => \N__49651\
        );

    \I__11146\ : InMux
    port map (
            O => \N__49657\,
            I => \N__49648\
        );

    \I__11145\ : Odrv4
    port map (
            O => \N__49654\,
            I => n1325
        );

    \I__11144\ : LocalMux
    port map (
            O => \N__49651\,
            I => n1325
        );

    \I__11143\ : LocalMux
    port map (
            O => \N__49648\,
            I => n1325
        );

    \I__11142\ : InMux
    port map (
            O => \N__49641\,
            I => \N__49638\
        );

    \I__11141\ : LocalMux
    port map (
            O => \N__49638\,
            I => \N__49635\
        );

    \I__11140\ : Span4Mux_h
    port map (
            O => \N__49635\,
            I => \N__49632\
        );

    \I__11139\ : Span4Mux_h
    port map (
            O => \N__49632\,
            I => \N__49629\
        );

    \I__11138\ : Odrv4
    port map (
            O => \N__49629\,
            I => n12
        );

    \I__11137\ : InMux
    port map (
            O => \N__49626\,
            I => \N__49612\
        );

    \I__11136\ : InMux
    port map (
            O => \N__49625\,
            I => \N__49612\
        );

    \I__11135\ : InMux
    port map (
            O => \N__49624\,
            I => \N__49612\
        );

    \I__11134\ : InMux
    port map (
            O => \N__49623\,
            I => \N__49612\
        );

    \I__11133\ : InMux
    port map (
            O => \N__49622\,
            I => \N__49607\
        );

    \I__11132\ : InMux
    port map (
            O => \N__49621\,
            I => \N__49594\
        );

    \I__11131\ : LocalMux
    port map (
            O => \N__49612\,
            I => \N__49586\
        );

    \I__11130\ : InMux
    port map (
            O => \N__49611\,
            I => \N__49581\
        );

    \I__11129\ : InMux
    port map (
            O => \N__49610\,
            I => \N__49581\
        );

    \I__11128\ : LocalMux
    port map (
            O => \N__49607\,
            I => \N__49577\
        );

    \I__11127\ : InMux
    port map (
            O => \N__49606\,
            I => \N__49574\
        );

    \I__11126\ : InMux
    port map (
            O => \N__49605\,
            I => \N__49569\
        );

    \I__11125\ : InMux
    port map (
            O => \N__49604\,
            I => \N__49569\
        );

    \I__11124\ : InMux
    port map (
            O => \N__49603\,
            I => \N__49566\
        );

    \I__11123\ : InMux
    port map (
            O => \N__49602\,
            I => \N__49561\
        );

    \I__11122\ : InMux
    port map (
            O => \N__49601\,
            I => \N__49561\
        );

    \I__11121\ : InMux
    port map (
            O => \N__49600\,
            I => \N__49557\
        );

    \I__11120\ : InMux
    port map (
            O => \N__49599\,
            I => \N__49554\
        );

    \I__11119\ : CascadeMux
    port map (
            O => \N__49598\,
            I => \N__49549\
        );

    \I__11118\ : CascadeMux
    port map (
            O => \N__49597\,
            I => \N__49543\
        );

    \I__11117\ : LocalMux
    port map (
            O => \N__49594\,
            I => \N__49535\
        );

    \I__11116\ : InMux
    port map (
            O => \N__49593\,
            I => \N__49528\
        );

    \I__11115\ : InMux
    port map (
            O => \N__49592\,
            I => \N__49528\
        );

    \I__11114\ : InMux
    port map (
            O => \N__49591\,
            I => \N__49528\
        );

    \I__11113\ : InMux
    port map (
            O => \N__49590\,
            I => \N__49523\
        );

    \I__11112\ : InMux
    port map (
            O => \N__49589\,
            I => \N__49523\
        );

    \I__11111\ : Span4Mux_h
    port map (
            O => \N__49586\,
            I => \N__49518\
        );

    \I__11110\ : LocalMux
    port map (
            O => \N__49581\,
            I => \N__49518\
        );

    \I__11109\ : CascadeMux
    port map (
            O => \N__49580\,
            I => \N__49514\
        );

    \I__11108\ : Span4Mux_v
    port map (
            O => \N__49577\,
            I => \N__49508\
        );

    \I__11107\ : LocalMux
    port map (
            O => \N__49574\,
            I => \N__49508\
        );

    \I__11106\ : LocalMux
    port map (
            O => \N__49569\,
            I => \N__49505\
        );

    \I__11105\ : LocalMux
    port map (
            O => \N__49566\,
            I => \N__49500\
        );

    \I__11104\ : LocalMux
    port map (
            O => \N__49561\,
            I => \N__49500\
        );

    \I__11103\ : InMux
    port map (
            O => \N__49560\,
            I => \N__49497\
        );

    \I__11102\ : LocalMux
    port map (
            O => \N__49557\,
            I => \N__49488\
        );

    \I__11101\ : LocalMux
    port map (
            O => \N__49554\,
            I => \N__49488\
        );

    \I__11100\ : CascadeMux
    port map (
            O => \N__49553\,
            I => \N__49485\
        );

    \I__11099\ : CascadeMux
    port map (
            O => \N__49552\,
            I => \N__49482\
        );

    \I__11098\ : InMux
    port map (
            O => \N__49549\,
            I => \N__49469\
        );

    \I__11097\ : InMux
    port map (
            O => \N__49548\,
            I => \N__49469\
        );

    \I__11096\ : InMux
    port map (
            O => \N__49547\,
            I => \N__49469\
        );

    \I__11095\ : InMux
    port map (
            O => \N__49546\,
            I => \N__49469\
        );

    \I__11094\ : InMux
    port map (
            O => \N__49543\,
            I => \N__49469\
        );

    \I__11093\ : InMux
    port map (
            O => \N__49542\,
            I => \N__49469\
        );

    \I__11092\ : InMux
    port map (
            O => \N__49541\,
            I => \N__49466\
        );

    \I__11091\ : InMux
    port map (
            O => \N__49540\,
            I => \N__49463\
        );

    \I__11090\ : InMux
    port map (
            O => \N__49539\,
            I => \N__49460\
        );

    \I__11089\ : InMux
    port map (
            O => \N__49538\,
            I => \N__49457\
        );

    \I__11088\ : Span4Mux_v
    port map (
            O => \N__49535\,
            I => \N__49452\
        );

    \I__11087\ : LocalMux
    port map (
            O => \N__49528\,
            I => \N__49452\
        );

    \I__11086\ : LocalMux
    port map (
            O => \N__49523\,
            I => \N__49447\
        );

    \I__11085\ : Span4Mux_h
    port map (
            O => \N__49518\,
            I => \N__49447\
        );

    \I__11084\ : InMux
    port map (
            O => \N__49517\,
            I => \N__49440\
        );

    \I__11083\ : InMux
    port map (
            O => \N__49514\,
            I => \N__49440\
        );

    \I__11082\ : InMux
    port map (
            O => \N__49513\,
            I => \N__49440\
        );

    \I__11081\ : Span4Mux_h
    port map (
            O => \N__49508\,
            I => \N__49437\
        );

    \I__11080\ : Span4Mux_h
    port map (
            O => \N__49505\,
            I => \N__49430\
        );

    \I__11079\ : Span4Mux_h
    port map (
            O => \N__49500\,
            I => \N__49430\
        );

    \I__11078\ : LocalMux
    port map (
            O => \N__49497\,
            I => \N__49430\
        );

    \I__11077\ : InMux
    port map (
            O => \N__49496\,
            I => \N__49427\
        );

    \I__11076\ : InMux
    port map (
            O => \N__49495\,
            I => \N__49420\
        );

    \I__11075\ : InMux
    port map (
            O => \N__49494\,
            I => \N__49420\
        );

    \I__11074\ : InMux
    port map (
            O => \N__49493\,
            I => \N__49420\
        );

    \I__11073\ : Span4Mux_h
    port map (
            O => \N__49488\,
            I => \N__49417\
        );

    \I__11072\ : InMux
    port map (
            O => \N__49485\,
            I => \N__49412\
        );

    \I__11071\ : InMux
    port map (
            O => \N__49482\,
            I => \N__49412\
        );

    \I__11070\ : LocalMux
    port map (
            O => \N__49469\,
            I => \N__49407\
        );

    \I__11069\ : LocalMux
    port map (
            O => \N__49466\,
            I => \N__49407\
        );

    \I__11068\ : LocalMux
    port map (
            O => \N__49463\,
            I => encoder0_position_31
        );

    \I__11067\ : LocalMux
    port map (
            O => \N__49460\,
            I => encoder0_position_31
        );

    \I__11066\ : LocalMux
    port map (
            O => \N__49457\,
            I => encoder0_position_31
        );

    \I__11065\ : Odrv4
    port map (
            O => \N__49452\,
            I => encoder0_position_31
        );

    \I__11064\ : Odrv4
    port map (
            O => \N__49447\,
            I => encoder0_position_31
        );

    \I__11063\ : LocalMux
    port map (
            O => \N__49440\,
            I => encoder0_position_31
        );

    \I__11062\ : Odrv4
    port map (
            O => \N__49437\,
            I => encoder0_position_31
        );

    \I__11061\ : Odrv4
    port map (
            O => \N__49430\,
            I => encoder0_position_31
        );

    \I__11060\ : LocalMux
    port map (
            O => \N__49427\,
            I => encoder0_position_31
        );

    \I__11059\ : LocalMux
    port map (
            O => \N__49420\,
            I => encoder0_position_31
        );

    \I__11058\ : Odrv4
    port map (
            O => \N__49417\,
            I => encoder0_position_31
        );

    \I__11057\ : LocalMux
    port map (
            O => \N__49412\,
            I => encoder0_position_31
        );

    \I__11056\ : Odrv12
    port map (
            O => \N__49407\,
            I => encoder0_position_31
        );

    \I__11055\ : CascadeMux
    port map (
            O => \N__49380\,
            I => \N__49377\
        );

    \I__11054\ : InMux
    port map (
            O => \N__49377\,
            I => \N__49373\
        );

    \I__11053\ : CascadeMux
    port map (
            O => \N__49376\,
            I => \N__49370\
        );

    \I__11052\ : LocalMux
    port map (
            O => \N__49373\,
            I => \N__49366\
        );

    \I__11051\ : InMux
    port map (
            O => \N__49370\,
            I => \N__49363\
        );

    \I__11050\ : InMux
    port map (
            O => \N__49369\,
            I => \N__49360\
        );

    \I__11049\ : Odrv4
    port map (
            O => \N__49366\,
            I => n1326
        );

    \I__11048\ : LocalMux
    port map (
            O => \N__49363\,
            I => n1326
        );

    \I__11047\ : LocalMux
    port map (
            O => \N__49360\,
            I => n1326
        );

    \I__11046\ : InMux
    port map (
            O => \N__49353\,
            I => \N__49350\
        );

    \I__11045\ : LocalMux
    port map (
            O => \N__49350\,
            I => n1195
        );

    \I__11044\ : CascadeMux
    port map (
            O => \N__49347\,
            I => \n1227_cascade_\
        );

    \I__11043\ : InMux
    port map (
            O => \N__49344\,
            I => \N__49341\
        );

    \I__11042\ : LocalMux
    port map (
            O => \N__49341\,
            I => n14476
        );

    \I__11041\ : InMux
    port map (
            O => \N__49338\,
            I => \N__49335\
        );

    \I__11040\ : LocalMux
    port map (
            O => \N__49335\,
            I => n1199
        );

    \I__11039\ : CascadeMux
    port map (
            O => \N__49332\,
            I => \N__49329\
        );

    \I__11038\ : InMux
    port map (
            O => \N__49329\,
            I => \N__49325\
        );

    \I__11037\ : CascadeMux
    port map (
            O => \N__49328\,
            I => \N__49322\
        );

    \I__11036\ : LocalMux
    port map (
            O => \N__49325\,
            I => \N__49319\
        );

    \I__11035\ : InMux
    port map (
            O => \N__49322\,
            I => \N__49316\
        );

    \I__11034\ : Odrv4
    port map (
            O => \N__49319\,
            I => n1132
        );

    \I__11033\ : LocalMux
    port map (
            O => \N__49316\,
            I => n1132
        );

    \I__11032\ : CascadeMux
    port map (
            O => \N__49311\,
            I => \N__49308\
        );

    \I__11031\ : InMux
    port map (
            O => \N__49308\,
            I => \N__49304\
        );

    \I__11030\ : InMux
    port map (
            O => \N__49307\,
            I => \N__49301\
        );

    \I__11029\ : LocalMux
    port map (
            O => \N__49304\,
            I => n1127
        );

    \I__11028\ : LocalMux
    port map (
            O => \N__49301\,
            I => n1127
        );

    \I__11027\ : InMux
    port map (
            O => \N__49296\,
            I => \N__49293\
        );

    \I__11026\ : LocalMux
    port map (
            O => \N__49293\,
            I => n1194
        );

    \I__11025\ : CascadeMux
    port map (
            O => \N__49290\,
            I => \n1127_cascade_\
        );

    \I__11024\ : InMux
    port map (
            O => \N__49287\,
            I => \N__49283\
        );

    \I__11023\ : CascadeMux
    port map (
            O => \N__49286\,
            I => \N__49280\
        );

    \I__11022\ : LocalMux
    port map (
            O => \N__49283\,
            I => \N__49277\
        );

    \I__11021\ : InMux
    port map (
            O => \N__49280\,
            I => \N__49274\
        );

    \I__11020\ : Odrv4
    port map (
            O => \N__49277\,
            I => n1328
        );

    \I__11019\ : LocalMux
    port map (
            O => \N__49274\,
            I => n1328
        );

    \I__11018\ : CascadeMux
    port map (
            O => \N__49269\,
            I => \n1328_cascade_\
        );

    \I__11017\ : InMux
    port map (
            O => \N__49266\,
            I => \N__49263\
        );

    \I__11016\ : LocalMux
    port map (
            O => \N__49263\,
            I => n14414
        );

    \I__11015\ : CascadeMux
    port map (
            O => \N__49260\,
            I => \N__49257\
        );

    \I__11014\ : InMux
    port map (
            O => \N__49257\,
            I => \N__49253\
        );

    \I__11013\ : CascadeMux
    port map (
            O => \N__49256\,
            I => \N__49250\
        );

    \I__11012\ : LocalMux
    port map (
            O => \N__49253\,
            I => \N__49246\
        );

    \I__11011\ : InMux
    port map (
            O => \N__49250\,
            I => \N__49243\
        );

    \I__11010\ : InMux
    port map (
            O => \N__49249\,
            I => \N__49240\
        );

    \I__11009\ : Odrv4
    port map (
            O => \N__49246\,
            I => n1327
        );

    \I__11008\ : LocalMux
    port map (
            O => \N__49243\,
            I => n1327
        );

    \I__11007\ : LocalMux
    port map (
            O => \N__49240\,
            I => n1327
        );

    \I__11006\ : CascadeMux
    port map (
            O => \N__49233\,
            I => \N__49229\
        );

    \I__11005\ : CascadeMux
    port map (
            O => \N__49232\,
            I => \N__49226\
        );

    \I__11004\ : InMux
    port map (
            O => \N__49229\,
            I => \N__49222\
        );

    \I__11003\ : InMux
    port map (
            O => \N__49226\,
            I => \N__49217\
        );

    \I__11002\ : InMux
    port map (
            O => \N__49225\,
            I => \N__49217\
        );

    \I__11001\ : LocalMux
    port map (
            O => \N__49222\,
            I => n1331
        );

    \I__11000\ : LocalMux
    port map (
            O => \N__49217\,
            I => n1331
        );

    \I__10999\ : CascadeMux
    port map (
            O => \N__49212\,
            I => \N__49209\
        );

    \I__10998\ : InMux
    port map (
            O => \N__49209\,
            I => \N__49205\
        );

    \I__10997\ : InMux
    port map (
            O => \N__49208\,
            I => \N__49202\
        );

    \I__10996\ : LocalMux
    port map (
            O => \N__49205\,
            I => n1332
        );

    \I__10995\ : LocalMux
    port map (
            O => \N__49202\,
            I => n1332
        );

    \I__10994\ : InMux
    port map (
            O => \N__49197\,
            I => \N__49194\
        );

    \I__10993\ : LocalMux
    port map (
            O => \N__49194\,
            I => n1399
        );

    \I__10992\ : CascadeMux
    port map (
            O => \N__49191\,
            I => \n1332_cascade_\
        );

    \I__10991\ : CascadeMux
    port map (
            O => \N__49188\,
            I => \N__49185\
        );

    \I__10990\ : InMux
    port map (
            O => \N__49185\,
            I => \N__49181\
        );

    \I__10989\ : CascadeMux
    port map (
            O => \N__49184\,
            I => \N__49178\
        );

    \I__10988\ : LocalMux
    port map (
            O => \N__49181\,
            I => \N__49174\
        );

    \I__10987\ : InMux
    port map (
            O => \N__49178\,
            I => \N__49171\
        );

    \I__10986\ : InMux
    port map (
            O => \N__49177\,
            I => \N__49168\
        );

    \I__10985\ : Odrv4
    port map (
            O => \N__49174\,
            I => n1329
        );

    \I__10984\ : LocalMux
    port map (
            O => \N__49171\,
            I => n1329
        );

    \I__10983\ : LocalMux
    port map (
            O => \N__49168\,
            I => n1329
        );

    \I__10982\ : InMux
    port map (
            O => \N__49161\,
            I => \N__49158\
        );

    \I__10981\ : LocalMux
    port map (
            O => \N__49158\,
            I => n11927
        );

    \I__10980\ : CascadeMux
    port map (
            O => \N__49155\,
            I => \n13723_cascade_\
        );

    \I__10979\ : InMux
    port map (
            O => \N__49152\,
            I => \N__49149\
        );

    \I__10978\ : LocalMux
    port map (
            O => \N__49149\,
            I => n1394
        );

    \I__10977\ : InMux
    port map (
            O => \N__49146\,
            I => \N__49143\
        );

    \I__10976\ : LocalMux
    port map (
            O => \N__49143\,
            I => n1391
        );

    \I__10975\ : InMux
    port map (
            O => \N__49140\,
            I => \N__49135\
        );

    \I__10974\ : InMux
    port map (
            O => \N__49139\,
            I => \N__49132\
        );

    \I__10973\ : InMux
    port map (
            O => \N__49138\,
            I => \N__49129\
        );

    \I__10972\ : LocalMux
    port map (
            O => \N__49135\,
            I => \N__49126\
        );

    \I__10971\ : LocalMux
    port map (
            O => \N__49132\,
            I => \N__49121\
        );

    \I__10970\ : LocalMux
    port map (
            O => \N__49129\,
            I => \N__49121\
        );

    \I__10969\ : Span4Mux_h
    port map (
            O => \N__49126\,
            I => \N__49118\
        );

    \I__10968\ : Odrv12
    port map (
            O => \N__49121\,
            I => n299
        );

    \I__10967\ : Odrv4
    port map (
            O => \N__49118\,
            I => n299
        );

    \I__10966\ : CascadeMux
    port map (
            O => \N__49113\,
            I => \n11925_cascade_\
        );

    \I__10965\ : InMux
    port map (
            O => \N__49110\,
            I => \N__49107\
        );

    \I__10964\ : LocalMux
    port map (
            O => \N__49107\,
            I => n1398
        );

    \I__10963\ : CascadeMux
    port map (
            O => \N__49104\,
            I => \n1430_cascade_\
        );

    \I__10962\ : InMux
    port map (
            O => \N__49101\,
            I => \N__49098\
        );

    \I__10961\ : LocalMux
    port map (
            O => \N__49098\,
            I => n13739
        );

    \I__10960\ : InMux
    port map (
            O => \N__49095\,
            I => \N__49092\
        );

    \I__10959\ : LocalMux
    port map (
            O => \N__49092\,
            I => n13720
        );

    \I__10958\ : InMux
    port map (
            O => \N__49089\,
            I => \N__49086\
        );

    \I__10957\ : LocalMux
    port map (
            O => \N__49086\,
            I => n1400
        );

    \I__10956\ : CascadeMux
    port map (
            O => \N__49083\,
            I => \n1356_cascade_\
        );

    \I__10955\ : CascadeMux
    port map (
            O => \N__49080\,
            I => \N__49076\
        );

    \I__10954\ : CascadeMux
    port map (
            O => \N__49079\,
            I => \N__49072\
        );

    \I__10953\ : InMux
    port map (
            O => \N__49076\,
            I => \N__49069\
        );

    \I__10952\ : InMux
    port map (
            O => \N__49075\,
            I => \N__49064\
        );

    \I__10951\ : InMux
    port map (
            O => \N__49072\,
            I => \N__49064\
        );

    \I__10950\ : LocalMux
    port map (
            O => \N__49069\,
            I => n1333
        );

    \I__10949\ : LocalMux
    port map (
            O => \N__49064\,
            I => n1333
        );

    \I__10948\ : CascadeMux
    port map (
            O => \N__49059\,
            I => \n1432_cascade_\
        );

    \I__10947\ : InMux
    port map (
            O => \N__49056\,
            I => \N__49053\
        );

    \I__10946\ : LocalMux
    port map (
            O => \N__49053\,
            I => n11923
        );

    \I__10945\ : InMux
    port map (
            O => \N__49050\,
            I => \N__49047\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__49047\,
            I => \N__49044\
        );

    \I__10943\ : Odrv4
    port map (
            O => \N__49044\,
            I => n1393
        );

    \I__10942\ : CascadeMux
    port map (
            O => \N__49041\,
            I => \n1425_cascade_\
        );

    \I__10941\ : InMux
    port map (
            O => \N__49038\,
            I => \N__49035\
        );

    \I__10940\ : LocalMux
    port map (
            O => \N__49035\,
            I => n14484
        );

    \I__10939\ : CascadeMux
    port map (
            O => \N__49032\,
            I => \n14490_cascade_\
        );

    \I__10938\ : CascadeMux
    port map (
            O => \N__49029\,
            I => \n1455_cascade_\
        );

    \I__10937\ : CascadeMux
    port map (
            O => \N__49026\,
            I => \n1531_cascade_\
        );

    \I__10936\ : CascadeMux
    port map (
            O => \N__49023\,
            I => \N__49020\
        );

    \I__10935\ : InMux
    port map (
            O => \N__49020\,
            I => \N__49017\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__49017\,
            I => n11997
        );

    \I__10933\ : CascadeMux
    port map (
            O => \N__49014\,
            I => \N__49011\
        );

    \I__10932\ : InMux
    port map (
            O => \N__49011\,
            I => \N__49008\
        );

    \I__10931\ : LocalMux
    port map (
            O => \N__49008\,
            I => \N__49004\
        );

    \I__10930\ : CascadeMux
    port map (
            O => \N__49007\,
            I => \N__49001\
        );

    \I__10929\ : Sp12to4
    port map (
            O => \N__49004\,
            I => \N__48994\
        );

    \I__10928\ : InMux
    port map (
            O => \N__49001\,
            I => \N__48988\
        );

    \I__10927\ : CascadeMux
    port map (
            O => \N__49000\,
            I => \N__48984\
        );

    \I__10926\ : CascadeMux
    port map (
            O => \N__48999\,
            I => \N__48981\
        );

    \I__10925\ : CascadeMux
    port map (
            O => \N__48998\,
            I => \N__48977\
        );

    \I__10924\ : CascadeMux
    port map (
            O => \N__48997\,
            I => \N__48973\
        );

    \I__10923\ : Span12Mux_v
    port map (
            O => \N__48994\,
            I => \N__48969\
        );

    \I__10922\ : InMux
    port map (
            O => \N__48993\,
            I => \N__48966\
        );

    \I__10921\ : InMux
    port map (
            O => \N__48992\,
            I => \N__48961\
        );

    \I__10920\ : InMux
    port map (
            O => \N__48991\,
            I => \N__48961\
        );

    \I__10919\ : LocalMux
    port map (
            O => \N__48988\,
            I => \N__48958\
        );

    \I__10918\ : InMux
    port map (
            O => \N__48987\,
            I => \N__48941\
        );

    \I__10917\ : InMux
    port map (
            O => \N__48984\,
            I => \N__48941\
        );

    \I__10916\ : InMux
    port map (
            O => \N__48981\,
            I => \N__48941\
        );

    \I__10915\ : InMux
    port map (
            O => \N__48980\,
            I => \N__48941\
        );

    \I__10914\ : InMux
    port map (
            O => \N__48977\,
            I => \N__48941\
        );

    \I__10913\ : InMux
    port map (
            O => \N__48976\,
            I => \N__48941\
        );

    \I__10912\ : InMux
    port map (
            O => \N__48973\,
            I => \N__48941\
        );

    \I__10911\ : InMux
    port map (
            O => \N__48972\,
            I => \N__48941\
        );

    \I__10910\ : Odrv12
    port map (
            O => \N__48969\,
            I => n1455
        );

    \I__10909\ : LocalMux
    port map (
            O => \N__48966\,
            I => n1455
        );

    \I__10908\ : LocalMux
    port map (
            O => \N__48961\,
            I => n1455
        );

    \I__10907\ : Odrv4
    port map (
            O => \N__48958\,
            I => n1455
        );

    \I__10906\ : LocalMux
    port map (
            O => \N__48941\,
            I => n1455
        );

    \I__10905\ : CascadeMux
    port map (
            O => \N__48930\,
            I => \N__48927\
        );

    \I__10904\ : InMux
    port map (
            O => \N__48927\,
            I => \N__48923\
        );

    \I__10903\ : CascadeMux
    port map (
            O => \N__48926\,
            I => \N__48920\
        );

    \I__10902\ : LocalMux
    port map (
            O => \N__48923\,
            I => \N__48917\
        );

    \I__10901\ : InMux
    port map (
            O => \N__48920\,
            I => \N__48914\
        );

    \I__10900\ : Span4Mux_v
    port map (
            O => \N__48917\,
            I => \N__48908\
        );

    \I__10899\ : LocalMux
    port map (
            O => \N__48914\,
            I => \N__48908\
        );

    \I__10898\ : InMux
    port map (
            O => \N__48913\,
            I => \N__48905\
        );

    \I__10897\ : Odrv4
    port map (
            O => \N__48908\,
            I => n1631_adj_611
        );

    \I__10896\ : LocalMux
    port map (
            O => \N__48905\,
            I => n1631_adj_611
        );

    \I__10895\ : InMux
    port map (
            O => \N__48900\,
            I => \N__48897\
        );

    \I__10894\ : LocalMux
    port map (
            O => \N__48897\,
            I => \N__48894\
        );

    \I__10893\ : Span4Mux_v
    port map (
            O => \N__48894\,
            I => \N__48890\
        );

    \I__10892\ : CascadeMux
    port map (
            O => \N__48893\,
            I => \N__48887\
        );

    \I__10891\ : Sp12to4
    port map (
            O => \N__48890\,
            I => \N__48881\
        );

    \I__10890\ : InMux
    port map (
            O => \N__48887\,
            I => \N__48878\
        );

    \I__10889\ : CascadeMux
    port map (
            O => \N__48886\,
            I => \N__48871\
        );

    \I__10888\ : CascadeMux
    port map (
            O => \N__48885\,
            I => \N__48867\
        );

    \I__10887\ : CascadeMux
    port map (
            O => \N__48884\,
            I => \N__48863\
        );

    \I__10886\ : Span12Mux_h
    port map (
            O => \N__48881\,
            I => \N__48857\
        );

    \I__10885\ : LocalMux
    port map (
            O => \N__48878\,
            I => \N__48854\
        );

    \I__10884\ : InMux
    port map (
            O => \N__48877\,
            I => \N__48851\
        );

    \I__10883\ : InMux
    port map (
            O => \N__48876\,
            I => \N__48844\
        );

    \I__10882\ : InMux
    port map (
            O => \N__48875\,
            I => \N__48844\
        );

    \I__10881\ : InMux
    port map (
            O => \N__48874\,
            I => \N__48844\
        );

    \I__10880\ : InMux
    port map (
            O => \N__48871\,
            I => \N__48839\
        );

    \I__10879\ : InMux
    port map (
            O => \N__48870\,
            I => \N__48839\
        );

    \I__10878\ : InMux
    port map (
            O => \N__48867\,
            I => \N__48834\
        );

    \I__10877\ : InMux
    port map (
            O => \N__48866\,
            I => \N__48834\
        );

    \I__10876\ : InMux
    port map (
            O => \N__48863\,
            I => \N__48825\
        );

    \I__10875\ : InMux
    port map (
            O => \N__48862\,
            I => \N__48825\
        );

    \I__10874\ : InMux
    port map (
            O => \N__48861\,
            I => \N__48825\
        );

    \I__10873\ : InMux
    port map (
            O => \N__48860\,
            I => \N__48825\
        );

    \I__10872\ : Odrv12
    port map (
            O => \N__48857\,
            I => n1554
        );

    \I__10871\ : Odrv4
    port map (
            O => \N__48854\,
            I => n1554
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__48851\,
            I => n1554
        );

    \I__10869\ : LocalMux
    port map (
            O => \N__48844\,
            I => n1554
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__48839\,
            I => n1554
        );

    \I__10867\ : LocalMux
    port map (
            O => \N__48834\,
            I => n1554
        );

    \I__10866\ : LocalMux
    port map (
            O => \N__48825\,
            I => n1554
        );

    \I__10865\ : InMux
    port map (
            O => \N__48810\,
            I => \N__48806\
        );

    \I__10864\ : CascadeMux
    port map (
            O => \N__48809\,
            I => \N__48803\
        );

    \I__10863\ : LocalMux
    port map (
            O => \N__48806\,
            I => \N__48800\
        );

    \I__10862\ : InMux
    port map (
            O => \N__48803\,
            I => \N__48797\
        );

    \I__10861\ : Span4Mux_v
    port map (
            O => \N__48800\,
            I => \N__48792\
        );

    \I__10860\ : LocalMux
    port map (
            O => \N__48797\,
            I => \N__48792\
        );

    \I__10859\ : Odrv4
    port map (
            O => \N__48792\,
            I => n1632_adj_612
        );

    \I__10858\ : InMux
    port map (
            O => \N__48789\,
            I => \N__48784\
        );

    \I__10857\ : InMux
    port map (
            O => \N__48788\,
            I => \N__48781\
        );

    \I__10856\ : InMux
    port map (
            O => \N__48787\,
            I => \N__48778\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__48784\,
            I => \N__48775\
        );

    \I__10854\ : LocalMux
    port map (
            O => \N__48781\,
            I => \N__48770\
        );

    \I__10853\ : LocalMux
    port map (
            O => \N__48778\,
            I => \N__48770\
        );

    \I__10852\ : Span4Mux_h
    port map (
            O => \N__48775\,
            I => \N__48767\
        );

    \I__10851\ : Span4Mux_h
    port map (
            O => \N__48770\,
            I => \N__48764\
        );

    \I__10850\ : Odrv4
    port map (
            O => \N__48767\,
            I => n302
        );

    \I__10849\ : Odrv4
    port map (
            O => \N__48764\,
            I => n302
        );

    \I__10848\ : CascadeMux
    port map (
            O => \N__48759\,
            I => \n1632_adj_612_cascade_\
        );

    \I__10847\ : CascadeMux
    port map (
            O => \N__48756\,
            I => \N__48753\
        );

    \I__10846\ : InMux
    port map (
            O => \N__48753\,
            I => \N__48750\
        );

    \I__10845\ : LocalMux
    port map (
            O => \N__48750\,
            I => \N__48746\
        );

    \I__10844\ : CascadeMux
    port map (
            O => \N__48749\,
            I => \N__48743\
        );

    \I__10843\ : Span4Mux_h
    port map (
            O => \N__48746\,
            I => \N__48739\
        );

    \I__10842\ : InMux
    port map (
            O => \N__48743\,
            I => \N__48736\
        );

    \I__10841\ : InMux
    port map (
            O => \N__48742\,
            I => \N__48733\
        );

    \I__10840\ : Odrv4
    port map (
            O => \N__48739\,
            I => n1633_adj_613
        );

    \I__10839\ : LocalMux
    port map (
            O => \N__48736\,
            I => n1633_adj_613
        );

    \I__10838\ : LocalMux
    port map (
            O => \N__48733\,
            I => n1633_adj_613
        );

    \I__10837\ : InMux
    port map (
            O => \N__48726\,
            I => \N__48723\
        );

    \I__10836\ : LocalMux
    port map (
            O => \N__48723\,
            I => n11919
        );

    \I__10835\ : InMux
    port map (
            O => \N__48720\,
            I => \PWM.n13047\
        );

    \I__10834\ : InMux
    port map (
            O => \N__48717\,
            I => \PWM.n13048\
        );

    \I__10833\ : InMux
    port map (
            O => \N__48714\,
            I => \PWM.n13049\
        );

    \I__10832\ : InMux
    port map (
            O => \N__48711\,
            I => \PWM.n13050\
        );

    \I__10831\ : InMux
    port map (
            O => \N__48708\,
            I => \PWM.n13051\
        );

    \I__10830\ : InMux
    port map (
            O => \N__48705\,
            I => \PWM.n13052\
        );

    \I__10829\ : SRMux
    port map (
            O => \N__48702\,
            I => \N__48699\
        );

    \I__10828\ : LocalMux
    port map (
            O => \N__48699\,
            I => \N__48696\
        );

    \I__10827\ : Span4Mux_h
    port map (
            O => \N__48696\,
            I => \N__48690\
        );

    \I__10826\ : SRMux
    port map (
            O => \N__48695\,
            I => \N__48687\
        );

    \I__10825\ : SRMux
    port map (
            O => \N__48694\,
            I => \N__48684\
        );

    \I__10824\ : SRMux
    port map (
            O => \N__48693\,
            I => \N__48681\
        );

    \I__10823\ : Odrv4
    port map (
            O => \N__48690\,
            I => \PWM.pwm_counter_31__N_407\
        );

    \I__10822\ : LocalMux
    port map (
            O => \N__48687\,
            I => \PWM.pwm_counter_31__N_407\
        );

    \I__10821\ : LocalMux
    port map (
            O => \N__48684\,
            I => \PWM.pwm_counter_31__N_407\
        );

    \I__10820\ : LocalMux
    port map (
            O => \N__48681\,
            I => \PWM.pwm_counter_31__N_407\
        );

    \I__10819\ : InMux
    port map (
            O => \N__48672\,
            I => \N__48668\
        );

    \I__10818\ : InMux
    port map (
            O => \N__48671\,
            I => \N__48665\
        );

    \I__10817\ : LocalMux
    port map (
            O => \N__48668\,
            I => pwm_counter_24
        );

    \I__10816\ : LocalMux
    port map (
            O => \N__48665\,
            I => pwm_counter_24
        );

    \I__10815\ : InMux
    port map (
            O => \N__48660\,
            I => \N__48656\
        );

    \I__10814\ : InMux
    port map (
            O => \N__48659\,
            I => \N__48653\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__48656\,
            I => pwm_counter_29
        );

    \I__10812\ : LocalMux
    port map (
            O => \N__48653\,
            I => pwm_counter_29
        );

    \I__10811\ : CascadeMux
    port map (
            O => \N__48648\,
            I => \N__48644\
        );

    \I__10810\ : InMux
    port map (
            O => \N__48647\,
            I => \N__48641\
        );

    \I__10809\ : InMux
    port map (
            O => \N__48644\,
            I => \N__48638\
        );

    \I__10808\ : LocalMux
    port map (
            O => \N__48641\,
            I => pwm_counter_27
        );

    \I__10807\ : LocalMux
    port map (
            O => \N__48638\,
            I => pwm_counter_27
        );

    \I__10806\ : InMux
    port map (
            O => \N__48633\,
            I => \N__48629\
        );

    \I__10805\ : InMux
    port map (
            O => \N__48632\,
            I => \N__48626\
        );

    \I__10804\ : LocalMux
    port map (
            O => \N__48629\,
            I => pwm_counter_26
        );

    \I__10803\ : LocalMux
    port map (
            O => \N__48626\,
            I => pwm_counter_26
        );

    \I__10802\ : InMux
    port map (
            O => \N__48621\,
            I => \N__48617\
        );

    \I__10801\ : InMux
    port map (
            O => \N__48620\,
            I => \N__48614\
        );

    \I__10800\ : LocalMux
    port map (
            O => \N__48617\,
            I => pwm_counter_30
        );

    \I__10799\ : LocalMux
    port map (
            O => \N__48614\,
            I => pwm_counter_30
        );

    \I__10798\ : InMux
    port map (
            O => \N__48609\,
            I => \N__48605\
        );

    \I__10797\ : InMux
    port map (
            O => \N__48608\,
            I => \N__48602\
        );

    \I__10796\ : LocalMux
    port map (
            O => \N__48605\,
            I => pwm_counter_25
        );

    \I__10795\ : LocalMux
    port map (
            O => \N__48602\,
            I => pwm_counter_25
        );

    \I__10794\ : CascadeMux
    port map (
            O => \N__48597\,
            I => \n12_adj_615_cascade_\
        );

    \I__10793\ : InMux
    port map (
            O => \N__48594\,
            I => \N__48590\
        );

    \I__10792\ : InMux
    port map (
            O => \N__48593\,
            I => \N__48587\
        );

    \I__10791\ : LocalMux
    port map (
            O => \N__48590\,
            I => pwm_counter_28
        );

    \I__10790\ : LocalMux
    port map (
            O => \N__48587\,
            I => pwm_counter_28
        );

    \I__10789\ : InMux
    port map (
            O => \N__48582\,
            I => \N__48579\
        );

    \I__10788\ : LocalMux
    port map (
            O => \N__48579\,
            I => \N__48574\
        );

    \I__10787\ : InMux
    port map (
            O => \N__48578\,
            I => \N__48571\
        );

    \I__10786\ : InMux
    port map (
            O => \N__48577\,
            I => \N__48568\
        );

    \I__10785\ : Span4Mux_s2_v
    port map (
            O => \N__48574\,
            I => \N__48565\
        );

    \I__10784\ : LocalMux
    port map (
            O => \N__48571\,
            I => pwm_counter_17
        );

    \I__10783\ : LocalMux
    port map (
            O => \N__48568\,
            I => pwm_counter_17
        );

    \I__10782\ : Odrv4
    port map (
            O => \N__48565\,
            I => pwm_counter_17
        );

    \I__10781\ : InMux
    port map (
            O => \N__48558\,
            I => \PWM.n13038\
        );

    \I__10780\ : InMux
    port map (
            O => \N__48555\,
            I => \N__48551\
        );

    \I__10779\ : InMux
    port map (
            O => \N__48554\,
            I => \N__48547\
        );

    \I__10778\ : LocalMux
    port map (
            O => \N__48551\,
            I => \N__48544\
        );

    \I__10777\ : InMux
    port map (
            O => \N__48550\,
            I => \N__48541\
        );

    \I__10776\ : LocalMux
    port map (
            O => \N__48547\,
            I => \N__48536\
        );

    \I__10775\ : Span4Mux_s2_v
    port map (
            O => \N__48544\,
            I => \N__48536\
        );

    \I__10774\ : LocalMux
    port map (
            O => \N__48541\,
            I => pwm_counter_18
        );

    \I__10773\ : Odrv4
    port map (
            O => \N__48536\,
            I => pwm_counter_18
        );

    \I__10772\ : InMux
    port map (
            O => \N__48531\,
            I => \PWM.n13039\
        );

    \I__10771\ : InMux
    port map (
            O => \N__48528\,
            I => \N__48523\
        );

    \I__10770\ : InMux
    port map (
            O => \N__48527\,
            I => \N__48520\
        );

    \I__10769\ : InMux
    port map (
            O => \N__48526\,
            I => \N__48517\
        );

    \I__10768\ : LocalMux
    port map (
            O => \N__48523\,
            I => \N__48514\
        );

    \I__10767\ : LocalMux
    port map (
            O => \N__48520\,
            I => pwm_counter_19
        );

    \I__10766\ : LocalMux
    port map (
            O => \N__48517\,
            I => pwm_counter_19
        );

    \I__10765\ : Odrv4
    port map (
            O => \N__48514\,
            I => pwm_counter_19
        );

    \I__10764\ : InMux
    port map (
            O => \N__48507\,
            I => \PWM.n13040\
        );

    \I__10763\ : InMux
    port map (
            O => \N__48504\,
            I => \N__48501\
        );

    \I__10762\ : LocalMux
    port map (
            O => \N__48501\,
            I => \N__48496\
        );

    \I__10761\ : InMux
    port map (
            O => \N__48500\,
            I => \N__48493\
        );

    \I__10760\ : InMux
    port map (
            O => \N__48499\,
            I => \N__48490\
        );

    \I__10759\ : Span4Mux_h
    port map (
            O => \N__48496\,
            I => \N__48487\
        );

    \I__10758\ : LocalMux
    port map (
            O => \N__48493\,
            I => pwm_counter_20
        );

    \I__10757\ : LocalMux
    port map (
            O => \N__48490\,
            I => pwm_counter_20
        );

    \I__10756\ : Odrv4
    port map (
            O => \N__48487\,
            I => pwm_counter_20
        );

    \I__10755\ : InMux
    port map (
            O => \N__48480\,
            I => \PWM.n13041\
        );

    \I__10754\ : CascadeMux
    port map (
            O => \N__48477\,
            I => \N__48472\
        );

    \I__10753\ : InMux
    port map (
            O => \N__48476\,
            I => \N__48469\
        );

    \I__10752\ : InMux
    port map (
            O => \N__48475\,
            I => \N__48464\
        );

    \I__10751\ : InMux
    port map (
            O => \N__48472\,
            I => \N__48464\
        );

    \I__10750\ : LocalMux
    port map (
            O => \N__48469\,
            I => \N__48459\
        );

    \I__10749\ : LocalMux
    port map (
            O => \N__48464\,
            I => \N__48456\
        );

    \I__10748\ : InMux
    port map (
            O => \N__48463\,
            I => \N__48453\
        );

    \I__10747\ : InMux
    port map (
            O => \N__48462\,
            I => \N__48450\
        );

    \I__10746\ : Span4Mux_h
    port map (
            O => \N__48459\,
            I => \N__48447\
        );

    \I__10745\ : Span4Mux_h
    port map (
            O => \N__48456\,
            I => \N__48444\
        );

    \I__10744\ : LocalMux
    port map (
            O => \N__48453\,
            I => pwm_counter_21
        );

    \I__10743\ : LocalMux
    port map (
            O => \N__48450\,
            I => pwm_counter_21
        );

    \I__10742\ : Odrv4
    port map (
            O => \N__48447\,
            I => pwm_counter_21
        );

    \I__10741\ : Odrv4
    port map (
            O => \N__48444\,
            I => pwm_counter_21
        );

    \I__10740\ : InMux
    port map (
            O => \N__48435\,
            I => \PWM.n13042\
        );

    \I__10739\ : InMux
    port map (
            O => \N__48432\,
            I => \N__48429\
        );

    \I__10738\ : LocalMux
    port map (
            O => \N__48429\,
            I => \N__48424\
        );

    \I__10737\ : InMux
    port map (
            O => \N__48428\,
            I => \N__48421\
        );

    \I__10736\ : InMux
    port map (
            O => \N__48427\,
            I => \N__48418\
        );

    \I__10735\ : Span4Mux_h
    port map (
            O => \N__48424\,
            I => \N__48415\
        );

    \I__10734\ : LocalMux
    port map (
            O => \N__48421\,
            I => pwm_counter_22
        );

    \I__10733\ : LocalMux
    port map (
            O => \N__48418\,
            I => pwm_counter_22
        );

    \I__10732\ : Odrv4
    port map (
            O => \N__48415\,
            I => pwm_counter_22
        );

    \I__10731\ : InMux
    port map (
            O => \N__48408\,
            I => \PWM.n13043\
        );

    \I__10730\ : InMux
    port map (
            O => \N__48405\,
            I => \PWM.n13044\
        );

    \I__10729\ : InMux
    port map (
            O => \N__48402\,
            I => \bfn_14_31_0_\
        );

    \I__10728\ : InMux
    port map (
            O => \N__48399\,
            I => \PWM.n13046\
        );

    \I__10727\ : InMux
    port map (
            O => \N__48396\,
            I => \N__48388\
        );

    \I__10726\ : InMux
    port map (
            O => \N__48395\,
            I => \N__48388\
        );

    \I__10725\ : InMux
    port map (
            O => \N__48394\,
            I => \N__48385\
        );

    \I__10724\ : InMux
    port map (
            O => \N__48393\,
            I => \N__48382\
        );

    \I__10723\ : LocalMux
    port map (
            O => \N__48388\,
            I => \N__48379\
        );

    \I__10722\ : LocalMux
    port map (
            O => \N__48385\,
            I => pwm_counter_9
        );

    \I__10721\ : LocalMux
    port map (
            O => \N__48382\,
            I => pwm_counter_9
        );

    \I__10720\ : Odrv12
    port map (
            O => \N__48379\,
            I => pwm_counter_9
        );

    \I__10719\ : InMux
    port map (
            O => \N__48372\,
            I => \PWM.n13030\
        );

    \I__10718\ : InMux
    port map (
            O => \N__48369\,
            I => \N__48364\
        );

    \I__10717\ : InMux
    port map (
            O => \N__48368\,
            I => \N__48361\
        );

    \I__10716\ : InMux
    port map (
            O => \N__48367\,
            I => \N__48358\
        );

    \I__10715\ : LocalMux
    port map (
            O => \N__48364\,
            I => \N__48355\
        );

    \I__10714\ : LocalMux
    port map (
            O => \N__48361\,
            I => pwm_counter_10
        );

    \I__10713\ : LocalMux
    port map (
            O => \N__48358\,
            I => pwm_counter_10
        );

    \I__10712\ : Odrv4
    port map (
            O => \N__48355\,
            I => pwm_counter_10
        );

    \I__10711\ : InMux
    port map (
            O => \N__48348\,
            I => \PWM.n13031\
        );

    \I__10710\ : InMux
    port map (
            O => \N__48345\,
            I => \N__48341\
        );

    \I__10709\ : InMux
    port map (
            O => \N__48344\,
            I => \N__48337\
        );

    \I__10708\ : LocalMux
    port map (
            O => \N__48341\,
            I => \N__48334\
        );

    \I__10707\ : InMux
    port map (
            O => \N__48340\,
            I => \N__48331\
        );

    \I__10706\ : LocalMux
    port map (
            O => \N__48337\,
            I => \N__48328\
        );

    \I__10705\ : Odrv4
    port map (
            O => \N__48334\,
            I => pwm_counter_11
        );

    \I__10704\ : LocalMux
    port map (
            O => \N__48331\,
            I => pwm_counter_11
        );

    \I__10703\ : Odrv4
    port map (
            O => \N__48328\,
            I => pwm_counter_11
        );

    \I__10702\ : InMux
    port map (
            O => \N__48321\,
            I => \PWM.n13032\
        );

    \I__10701\ : InMux
    port map (
            O => \N__48318\,
            I => \N__48315\
        );

    \I__10700\ : LocalMux
    port map (
            O => \N__48315\,
            I => \N__48310\
        );

    \I__10699\ : InMux
    port map (
            O => \N__48314\,
            I => \N__48307\
        );

    \I__10698\ : InMux
    port map (
            O => \N__48313\,
            I => \N__48304\
        );

    \I__10697\ : Span4Mux_s3_v
    port map (
            O => \N__48310\,
            I => \N__48301\
        );

    \I__10696\ : LocalMux
    port map (
            O => \N__48307\,
            I => pwm_counter_12
        );

    \I__10695\ : LocalMux
    port map (
            O => \N__48304\,
            I => pwm_counter_12
        );

    \I__10694\ : Odrv4
    port map (
            O => \N__48301\,
            I => pwm_counter_12
        );

    \I__10693\ : InMux
    port map (
            O => \N__48294\,
            I => \PWM.n13033\
        );

    \I__10692\ : InMux
    port map (
            O => \N__48291\,
            I => \N__48286\
        );

    \I__10691\ : InMux
    port map (
            O => \N__48290\,
            I => \N__48283\
        );

    \I__10690\ : InMux
    port map (
            O => \N__48289\,
            I => \N__48280\
        );

    \I__10689\ : LocalMux
    port map (
            O => \N__48286\,
            I => pwm_counter_13
        );

    \I__10688\ : LocalMux
    port map (
            O => \N__48283\,
            I => pwm_counter_13
        );

    \I__10687\ : LocalMux
    port map (
            O => \N__48280\,
            I => pwm_counter_13
        );

    \I__10686\ : InMux
    port map (
            O => \N__48273\,
            I => \PWM.n13034\
        );

    \I__10685\ : CascadeMux
    port map (
            O => \N__48270\,
            I => \N__48267\
        );

    \I__10684\ : InMux
    port map (
            O => \N__48267\,
            I => \N__48262\
        );

    \I__10683\ : InMux
    port map (
            O => \N__48266\,
            I => \N__48259\
        );

    \I__10682\ : InMux
    port map (
            O => \N__48265\,
            I => \N__48256\
        );

    \I__10681\ : LocalMux
    port map (
            O => \N__48262\,
            I => \N__48251\
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__48259\,
            I => \N__48251\
        );

    \I__10679\ : LocalMux
    port map (
            O => \N__48256\,
            I => pwm_counter_14
        );

    \I__10678\ : Odrv4
    port map (
            O => \N__48251\,
            I => pwm_counter_14
        );

    \I__10677\ : InMux
    port map (
            O => \N__48246\,
            I => \PWM.n13035\
        );

    \I__10676\ : CascadeMux
    port map (
            O => \N__48243\,
            I => \N__48239\
        );

    \I__10675\ : InMux
    port map (
            O => \N__48242\,
            I => \N__48236\
        );

    \I__10674\ : InMux
    port map (
            O => \N__48239\,
            I => \N__48232\
        );

    \I__10673\ : LocalMux
    port map (
            O => \N__48236\,
            I => \N__48229\
        );

    \I__10672\ : InMux
    port map (
            O => \N__48235\,
            I => \N__48226\
        );

    \I__10671\ : LocalMux
    port map (
            O => \N__48232\,
            I => \N__48221\
        );

    \I__10670\ : Span4Mux_h
    port map (
            O => \N__48229\,
            I => \N__48221\
        );

    \I__10669\ : LocalMux
    port map (
            O => \N__48226\,
            I => pwm_counter_15
        );

    \I__10668\ : Odrv4
    port map (
            O => \N__48221\,
            I => pwm_counter_15
        );

    \I__10667\ : InMux
    port map (
            O => \N__48216\,
            I => \PWM.n13036\
        );

    \I__10666\ : InMux
    port map (
            O => \N__48213\,
            I => \N__48203\
        );

    \I__10665\ : InMux
    port map (
            O => \N__48212\,
            I => \N__48203\
        );

    \I__10664\ : InMux
    port map (
            O => \N__48211\,
            I => \N__48203\
        );

    \I__10663\ : CascadeMux
    port map (
            O => \N__48210\,
            I => \N__48199\
        );

    \I__10662\ : LocalMux
    port map (
            O => \N__48203\,
            I => \N__48196\
        );

    \I__10661\ : InMux
    port map (
            O => \N__48202\,
            I => \N__48193\
        );

    \I__10660\ : InMux
    port map (
            O => \N__48199\,
            I => \N__48190\
        );

    \I__10659\ : Span4Mux_s2_v
    port map (
            O => \N__48196\,
            I => \N__48187\
        );

    \I__10658\ : LocalMux
    port map (
            O => \N__48193\,
            I => pwm_counter_16
        );

    \I__10657\ : LocalMux
    port map (
            O => \N__48190\,
            I => pwm_counter_16
        );

    \I__10656\ : Odrv4
    port map (
            O => \N__48187\,
            I => pwm_counter_16
        );

    \I__10655\ : InMux
    port map (
            O => \N__48180\,
            I => \bfn_14_30_0_\
        );

    \I__10654\ : CascadeMux
    port map (
            O => \N__48177\,
            I => \N__48174\
        );

    \I__10653\ : InMux
    port map (
            O => \N__48174\,
            I => \N__48170\
        );

    \I__10652\ : InMux
    port map (
            O => \N__48173\,
            I => \N__48167\
        );

    \I__10651\ : LocalMux
    port map (
            O => \N__48170\,
            I => \N__48164\
        );

    \I__10650\ : LocalMux
    port map (
            O => \N__48167\,
            I => pwm_counter_0
        );

    \I__10649\ : Odrv4
    port map (
            O => \N__48164\,
            I => pwm_counter_0
        );

    \I__10648\ : InMux
    port map (
            O => \N__48159\,
            I => \bfn_14_28_0_\
        );

    \I__10647\ : InMux
    port map (
            O => \N__48156\,
            I => \N__48152\
        );

    \I__10646\ : InMux
    port map (
            O => \N__48155\,
            I => \N__48149\
        );

    \I__10645\ : LocalMux
    port map (
            O => \N__48152\,
            I => \N__48146\
        );

    \I__10644\ : LocalMux
    port map (
            O => \N__48149\,
            I => pwm_counter_1
        );

    \I__10643\ : Odrv4
    port map (
            O => \N__48146\,
            I => pwm_counter_1
        );

    \I__10642\ : InMux
    port map (
            O => \N__48141\,
            I => \PWM.n13022\
        );

    \I__10641\ : CascadeMux
    port map (
            O => \N__48138\,
            I => \N__48134\
        );

    \I__10640\ : InMux
    port map (
            O => \N__48137\,
            I => \N__48131\
        );

    \I__10639\ : InMux
    port map (
            O => \N__48134\,
            I => \N__48128\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__48131\,
            I => pwm_counter_2
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__48128\,
            I => pwm_counter_2
        );

    \I__10636\ : InMux
    port map (
            O => \N__48123\,
            I => \PWM.n13023\
        );

    \I__10635\ : InMux
    port map (
            O => \N__48120\,
            I => \N__48115\
        );

    \I__10634\ : InMux
    port map (
            O => \N__48119\,
            I => \N__48110\
        );

    \I__10633\ : InMux
    port map (
            O => \N__48118\,
            I => \N__48110\
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__48115\,
            I => pwm_counter_3
        );

    \I__10631\ : LocalMux
    port map (
            O => \N__48110\,
            I => pwm_counter_3
        );

    \I__10630\ : InMux
    port map (
            O => \N__48105\,
            I => \PWM.n13024\
        );

    \I__10629\ : InMux
    port map (
            O => \N__48102\,
            I => \N__48099\
        );

    \I__10628\ : LocalMux
    port map (
            O => \N__48099\,
            I => \N__48095\
        );

    \I__10627\ : InMux
    port map (
            O => \N__48098\,
            I => \N__48092\
        );

    \I__10626\ : Span4Mux_h
    port map (
            O => \N__48095\,
            I => \N__48089\
        );

    \I__10625\ : LocalMux
    port map (
            O => \N__48092\,
            I => pwm_counter_4
        );

    \I__10624\ : Odrv4
    port map (
            O => \N__48089\,
            I => pwm_counter_4
        );

    \I__10623\ : InMux
    port map (
            O => \N__48084\,
            I => \PWM.n13025\
        );

    \I__10622\ : InMux
    port map (
            O => \N__48081\,
            I => \N__48076\
        );

    \I__10621\ : InMux
    port map (
            O => \N__48080\,
            I => \N__48073\
        );

    \I__10620\ : InMux
    port map (
            O => \N__48079\,
            I => \N__48070\
        );

    \I__10619\ : LocalMux
    port map (
            O => \N__48076\,
            I => \N__48067\
        );

    \I__10618\ : LocalMux
    port map (
            O => \N__48073\,
            I => pwm_counter_5
        );

    \I__10617\ : LocalMux
    port map (
            O => \N__48070\,
            I => pwm_counter_5
        );

    \I__10616\ : Odrv4
    port map (
            O => \N__48067\,
            I => pwm_counter_5
        );

    \I__10615\ : InMux
    port map (
            O => \N__48060\,
            I => \PWM.n13026\
        );

    \I__10614\ : InMux
    port map (
            O => \N__48057\,
            I => \N__48053\
        );

    \I__10613\ : InMux
    port map (
            O => \N__48056\,
            I => \N__48050\
        );

    \I__10612\ : LocalMux
    port map (
            O => \N__48053\,
            I => \N__48045\
        );

    \I__10611\ : LocalMux
    port map (
            O => \N__48050\,
            I => \N__48042\
        );

    \I__10610\ : InMux
    port map (
            O => \N__48049\,
            I => \N__48039\
        );

    \I__10609\ : InMux
    port map (
            O => \N__48048\,
            I => \N__48036\
        );

    \I__10608\ : Span4Mux_h
    port map (
            O => \N__48045\,
            I => \N__48033\
        );

    \I__10607\ : Span4Mux_h
    port map (
            O => \N__48042\,
            I => \N__48030\
        );

    \I__10606\ : LocalMux
    port map (
            O => \N__48039\,
            I => pwm_counter_6
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__48036\,
            I => pwm_counter_6
        );

    \I__10604\ : Odrv4
    port map (
            O => \N__48033\,
            I => pwm_counter_6
        );

    \I__10603\ : Odrv4
    port map (
            O => \N__48030\,
            I => pwm_counter_6
        );

    \I__10602\ : InMux
    port map (
            O => \N__48021\,
            I => \PWM.n13027\
        );

    \I__10601\ : InMux
    port map (
            O => \N__48018\,
            I => \N__48014\
        );

    \I__10600\ : InMux
    port map (
            O => \N__48017\,
            I => \N__48011\
        );

    \I__10599\ : LocalMux
    port map (
            O => \N__48014\,
            I => \N__48006\
        );

    \I__10598\ : LocalMux
    port map (
            O => \N__48011\,
            I => \N__48003\
        );

    \I__10597\ : InMux
    port map (
            O => \N__48010\,
            I => \N__48000\
        );

    \I__10596\ : InMux
    port map (
            O => \N__48009\,
            I => \N__47997\
        );

    \I__10595\ : Span4Mux_h
    port map (
            O => \N__48006\,
            I => \N__47994\
        );

    \I__10594\ : Span4Mux_h
    port map (
            O => \N__48003\,
            I => \N__47991\
        );

    \I__10593\ : LocalMux
    port map (
            O => \N__48000\,
            I => pwm_counter_7
        );

    \I__10592\ : LocalMux
    port map (
            O => \N__47997\,
            I => pwm_counter_7
        );

    \I__10591\ : Odrv4
    port map (
            O => \N__47994\,
            I => pwm_counter_7
        );

    \I__10590\ : Odrv4
    port map (
            O => \N__47991\,
            I => pwm_counter_7
        );

    \I__10589\ : InMux
    port map (
            O => \N__47982\,
            I => \PWM.n13028\
        );

    \I__10588\ : InMux
    port map (
            O => \N__47979\,
            I => \N__47974\
        );

    \I__10587\ : InMux
    port map (
            O => \N__47978\,
            I => \N__47971\
        );

    \I__10586\ : CascadeMux
    port map (
            O => \N__47977\,
            I => \N__47968\
        );

    \I__10585\ : LocalMux
    port map (
            O => \N__47974\,
            I => \N__47964\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__47971\,
            I => \N__47961\
        );

    \I__10583\ : InMux
    port map (
            O => \N__47968\,
            I => \N__47958\
        );

    \I__10582\ : InMux
    port map (
            O => \N__47967\,
            I => \N__47955\
        );

    \I__10581\ : Span4Mux_h
    port map (
            O => \N__47964\,
            I => \N__47950\
        );

    \I__10580\ : Span4Mux_h
    port map (
            O => \N__47961\,
            I => \N__47950\
        );

    \I__10579\ : LocalMux
    port map (
            O => \N__47958\,
            I => pwm_counter_8
        );

    \I__10578\ : LocalMux
    port map (
            O => \N__47955\,
            I => pwm_counter_8
        );

    \I__10577\ : Odrv4
    port map (
            O => \N__47950\,
            I => pwm_counter_8
        );

    \I__10576\ : InMux
    port map (
            O => \N__47943\,
            I => \bfn_14_29_0_\
        );

    \I__10575\ : InMux
    port map (
            O => \N__47940\,
            I => \N__47937\
        );

    \I__10574\ : LocalMux
    port map (
            O => \N__47937\,
            I => \N__47934\
        );

    \I__10573\ : Span4Mux_h
    port map (
            O => \N__47934\,
            I => \N__47931\
        );

    \I__10572\ : Odrv4
    port map (
            O => \N__47931\,
            I => pwm_setpoint_1
        );

    \I__10571\ : CascadeMux
    port map (
            O => \N__47928\,
            I => \n16_adj_679_cascade_\
        );

    \I__10570\ : InMux
    port map (
            O => \N__47925\,
            I => \N__47922\
        );

    \I__10569\ : LocalMux
    port map (
            O => \N__47922\,
            I => n15_adj_680
        );

    \I__10568\ : InMux
    port map (
            O => \N__47919\,
            I => \N__47916\
        );

    \I__10567\ : LocalMux
    port map (
            O => \N__47916\,
            I => n25_adj_652
        );

    \I__10566\ : CascadeMux
    port map (
            O => \N__47913\,
            I => \n16_adj_619_cascade_\
        );

    \I__10565\ : InMux
    port map (
            O => \N__47910\,
            I => \N__47907\
        );

    \I__10564\ : LocalMux
    port map (
            O => \N__47907\,
            I => n22_adj_617
        );

    \I__10563\ : InMux
    port map (
            O => \N__47904\,
            I => \N__47901\
        );

    \I__10562\ : LocalMux
    port map (
            O => \N__47901\,
            I => \N__47898\
        );

    \I__10561\ : Odrv4
    port map (
            O => \N__47898\,
            I => n24_adj_616
        );

    \I__10560\ : InMux
    port map (
            O => \N__47895\,
            I => \N__47892\
        );

    \I__10559\ : LocalMux
    port map (
            O => \N__47892\,
            I => \N__47889\
        );

    \I__10558\ : Span4Mux_h
    port map (
            O => \N__47889\,
            I => \N__47886\
        );

    \I__10557\ : Odrv4
    port map (
            O => \N__47886\,
            I => encoder0_position_scaled_16
        );

    \I__10556\ : InMux
    port map (
            O => \N__47883\,
            I => \N__47880\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__47880\,
            I => \N__47877\
        );

    \I__10554\ : Odrv4
    port map (
            O => \N__47877\,
            I => n9_adj_567
        );

    \I__10553\ : InMux
    port map (
            O => \N__47874\,
            I => \N__47870\
        );

    \I__10552\ : InMux
    port map (
            O => \N__47873\,
            I => \N__47867\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__47870\,
            I => \N__47864\
        );

    \I__10550\ : LocalMux
    port map (
            O => \N__47867\,
            I => \N__47861\
        );

    \I__10549\ : Span4Mux_h
    port map (
            O => \N__47864\,
            I => \N__47858\
        );

    \I__10548\ : Span4Mux_h
    port map (
            O => \N__47861\,
            I => \N__47855\
        );

    \I__10547\ : Odrv4
    port map (
            O => \N__47858\,
            I => duty_1
        );

    \I__10546\ : Odrv4
    port map (
            O => \N__47855\,
            I => duty_1
        );

    \I__10545\ : InMux
    port map (
            O => \N__47850\,
            I => \N__47847\
        );

    \I__10544\ : LocalMux
    port map (
            O => \N__47847\,
            I => \N__47844\
        );

    \I__10543\ : Span4Mux_h
    port map (
            O => \N__47844\,
            I => \N__47841\
        );

    \I__10542\ : Odrv4
    port map (
            O => \N__47841\,
            I => n24_adj_596
        );

    \I__10541\ : SRMux
    port map (
            O => \N__47838\,
            I => \N__47832\
        );

    \I__10540\ : InMux
    port map (
            O => \N__47837\,
            I => \N__47832\
        );

    \I__10539\ : LocalMux
    port map (
            O => \N__47832\,
            I => \N__47829\
        );

    \I__10538\ : Span4Mux_h
    port map (
            O => \N__47829\,
            I => \N__47826\
        );

    \I__10537\ : Odrv4
    port map (
            O => \N__47826\,
            I => \pwm_setpoint_23__N_195\
        );

    \I__10536\ : CascadeMux
    port map (
            O => \N__47823\,
            I => \n13197_cascade_\
        );

    \I__10535\ : InMux
    port map (
            O => \N__47820\,
            I => \N__47817\
        );

    \I__10534\ : LocalMux
    port map (
            O => \N__47817\,
            I => n24_adj_653
        );

    \I__10533\ : CascadeMux
    port map (
            O => \N__47814\,
            I => \direction_N_342_cascade_\
        );

    \I__10532\ : InMux
    port map (
            O => \N__47811\,
            I => \N__47808\
        );

    \I__10531\ : LocalMux
    port map (
            O => \N__47808\,
            I => \direction_N_342\
        );

    \I__10530\ : InMux
    port map (
            O => \N__47805\,
            I => \N__47802\
        );

    \I__10529\ : LocalMux
    port map (
            O => \N__47802\,
            I => n13675
        );

    \I__10528\ : CascadeMux
    port map (
            O => \N__47799\,
            I => \n23_adj_709_cascade_\
        );

    \I__10527\ : InMux
    port map (
            O => \N__47796\,
            I => \N__47793\
        );

    \I__10526\ : LocalMux
    port map (
            O => \N__47793\,
            I => n25_adj_707
        );

    \I__10525\ : InMux
    port map (
            O => \N__47790\,
            I => \N__47786\
        );

    \I__10524\ : InMux
    port map (
            O => \N__47789\,
            I => \N__47783\
        );

    \I__10523\ : LocalMux
    port map (
            O => \N__47786\,
            I => \direction_N_340\
        );

    \I__10522\ : LocalMux
    port map (
            O => \N__47783\,
            I => \direction_N_340\
        );

    \I__10521\ : InMux
    port map (
            O => \N__47778\,
            I => \N__47775\
        );

    \I__10520\ : LocalMux
    port map (
            O => \N__47775\,
            I => n24_adj_708
        );

    \I__10519\ : InMux
    port map (
            O => \N__47772\,
            I => \N__47769\
        );

    \I__10518\ : LocalMux
    port map (
            O => \N__47769\,
            I => n23_adj_654
        );

    \I__10517\ : InMux
    port map (
            O => \N__47766\,
            I => \N__47763\
        );

    \I__10516\ : LocalMux
    port map (
            O => \N__47763\,
            I => \N__47760\
        );

    \I__10515\ : Odrv12
    port map (
            O => \N__47760\,
            I => \pwm_setpoint_23_N_171_1\
        );

    \I__10514\ : InMux
    port map (
            O => \N__47757\,
            I => n12527
        );

    \I__10513\ : InMux
    port map (
            O => \N__47754\,
            I => n12528
        );

    \I__10512\ : InMux
    port map (
            O => \N__47751\,
            I => \bfn_14_24_0_\
        );

    \I__10511\ : InMux
    port map (
            O => \N__47748\,
            I => n12530
        );

    \I__10510\ : InMux
    port map (
            O => \N__47745\,
            I => \N__47742\
        );

    \I__10509\ : LocalMux
    port map (
            O => \N__47742\,
            I => \N__47739\
        );

    \I__10508\ : Span12Mux_s8_v
    port map (
            O => \N__47739\,
            I => \N__47735\
        );

    \I__10507\ : InMux
    port map (
            O => \N__47738\,
            I => \N__47732\
        );

    \I__10506\ : Odrv12
    port map (
            O => \N__47735\,
            I => n15522
        );

    \I__10505\ : LocalMux
    port map (
            O => \N__47732\,
            I => n15522
        );

    \I__10504\ : InMux
    port map (
            O => \N__47727\,
            I => \N__47724\
        );

    \I__10503\ : LocalMux
    port map (
            O => \N__47724\,
            I => \N__47721\
        );

    \I__10502\ : Span4Mux_h
    port map (
            O => \N__47721\,
            I => \N__47718\
        );

    \I__10501\ : Odrv4
    port map (
            O => \N__47718\,
            I => n13
        );

    \I__10500\ : CascadeMux
    port map (
            O => \N__47715\,
            I => \N__47712\
        );

    \I__10499\ : InMux
    port map (
            O => \N__47712\,
            I => \N__47708\
        );

    \I__10498\ : CascadeMux
    port map (
            O => \N__47711\,
            I => \N__47704\
        );

    \I__10497\ : LocalMux
    port map (
            O => \N__47708\,
            I => \N__47701\
        );

    \I__10496\ : InMux
    port map (
            O => \N__47707\,
            I => \N__47698\
        );

    \I__10495\ : InMux
    port map (
            O => \N__47704\,
            I => \N__47695\
        );

    \I__10494\ : Span4Mux_v
    port map (
            O => \N__47701\,
            I => \N__47692\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__47698\,
            I => \N__47689\
        );

    \I__10492\ : LocalMux
    port map (
            O => \N__47695\,
            I => encoder0_position_20
        );

    \I__10491\ : Odrv4
    port map (
            O => \N__47692\,
            I => encoder0_position_20
        );

    \I__10490\ : Odrv4
    port map (
            O => \N__47689\,
            I => encoder0_position_20
        );

    \I__10489\ : CascadeMux
    port map (
            O => \N__47682\,
            I => \N__47678\
        );

    \I__10488\ : InMux
    port map (
            O => \N__47681\,
            I => \N__47675\
        );

    \I__10487\ : InMux
    port map (
            O => \N__47678\,
            I => \N__47672\
        );

    \I__10486\ : LocalMux
    port map (
            O => \N__47675\,
            I => \N__47669\
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__47672\,
            I => n1125
        );

    \I__10484\ : Odrv4
    port map (
            O => \N__47669\,
            I => n1125
        );

    \I__10483\ : CascadeMux
    port map (
            O => \N__47664\,
            I => \n20_adj_618_cascade_\
        );

    \I__10482\ : InMux
    port map (
            O => \N__47661\,
            I => \N__47658\
        );

    \I__10481\ : LocalMux
    port map (
            O => \N__47658\,
            I => \N__47655\
        );

    \I__10480\ : Odrv4
    port map (
            O => \N__47655\,
            I => n13197
        );

    \I__10479\ : CascadeMux
    port map (
            O => \N__47652\,
            I => \n1233_cascade_\
        );

    \I__10478\ : InMux
    port map (
            O => \N__47649\,
            I => \N__47644\
        );

    \I__10477\ : InMux
    port map (
            O => \N__47648\,
            I => \N__47641\
        );

    \I__10476\ : InMux
    port map (
            O => \N__47647\,
            I => \N__47638\
        );

    \I__10475\ : LocalMux
    port map (
            O => \N__47644\,
            I => \N__47631\
        );

    \I__10474\ : LocalMux
    port map (
            O => \N__47641\,
            I => \N__47631\
        );

    \I__10473\ : LocalMux
    port map (
            O => \N__47638\,
            I => \N__47631\
        );

    \I__10472\ : Span4Mux_v
    port map (
            O => \N__47631\,
            I => \N__47628\
        );

    \I__10471\ : Odrv4
    port map (
            O => \N__47628\,
            I => n297
        );

    \I__10470\ : InMux
    port map (
            O => \N__47625\,
            I => \N__47622\
        );

    \I__10469\ : LocalMux
    port map (
            O => \N__47622\,
            I => n1201
        );

    \I__10468\ : InMux
    port map (
            O => \N__47619\,
            I => \bfn_14_23_0_\
        );

    \I__10467\ : CascadeMux
    port map (
            O => \N__47616\,
            I => \N__47612\
        );

    \I__10466\ : InMux
    port map (
            O => \N__47615\,
            I => \N__47608\
        );

    \I__10465\ : InMux
    port map (
            O => \N__47612\,
            I => \N__47605\
        );

    \I__10464\ : InMux
    port map (
            O => \N__47611\,
            I => \N__47602\
        );

    \I__10463\ : LocalMux
    port map (
            O => \N__47608\,
            I => n1133
        );

    \I__10462\ : LocalMux
    port map (
            O => \N__47605\,
            I => n1133
        );

    \I__10461\ : LocalMux
    port map (
            O => \N__47602\,
            I => n1133
        );

    \I__10460\ : CascadeMux
    port map (
            O => \N__47595\,
            I => \N__47592\
        );

    \I__10459\ : InMux
    port map (
            O => \N__47592\,
            I => \N__47589\
        );

    \I__10458\ : LocalMux
    port map (
            O => \N__47589\,
            I => n1200
        );

    \I__10457\ : InMux
    port map (
            O => \N__47586\,
            I => n12522
        );

    \I__10456\ : InMux
    port map (
            O => \N__47583\,
            I => n12523
        );

    \I__10455\ : CascadeMux
    port map (
            O => \N__47580\,
            I => \N__47576\
        );

    \I__10454\ : CascadeMux
    port map (
            O => \N__47579\,
            I => \N__47573\
        );

    \I__10453\ : InMux
    port map (
            O => \N__47576\,
            I => \N__47569\
        );

    \I__10452\ : InMux
    port map (
            O => \N__47573\,
            I => \N__47566\
        );

    \I__10451\ : InMux
    port map (
            O => \N__47572\,
            I => \N__47563\
        );

    \I__10450\ : LocalMux
    port map (
            O => \N__47569\,
            I => n1131
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__47566\,
            I => n1131
        );

    \I__10448\ : LocalMux
    port map (
            O => \N__47563\,
            I => n1131
        );

    \I__10447\ : InMux
    port map (
            O => \N__47556\,
            I => \N__47553\
        );

    \I__10446\ : LocalMux
    port map (
            O => \N__47553\,
            I => \N__47550\
        );

    \I__10445\ : Odrv4
    port map (
            O => \N__47550\,
            I => n1198
        );

    \I__10444\ : InMux
    port map (
            O => \N__47547\,
            I => n12524
        );

    \I__10443\ : CascadeMux
    port map (
            O => \N__47544\,
            I => \N__47540\
        );

    \I__10442\ : CascadeMux
    port map (
            O => \N__47543\,
            I => \N__47537\
        );

    \I__10441\ : InMux
    port map (
            O => \N__47540\,
            I => \N__47533\
        );

    \I__10440\ : InMux
    port map (
            O => \N__47537\,
            I => \N__47530\
        );

    \I__10439\ : InMux
    port map (
            O => \N__47536\,
            I => \N__47527\
        );

    \I__10438\ : LocalMux
    port map (
            O => \N__47533\,
            I => n1130
        );

    \I__10437\ : LocalMux
    port map (
            O => \N__47530\,
            I => n1130
        );

    \I__10436\ : LocalMux
    port map (
            O => \N__47527\,
            I => n1130
        );

    \I__10435\ : InMux
    port map (
            O => \N__47520\,
            I => \N__47517\
        );

    \I__10434\ : LocalMux
    port map (
            O => \N__47517\,
            I => n1197
        );

    \I__10433\ : InMux
    port map (
            O => \N__47514\,
            I => n12525
        );

    \I__10432\ : InMux
    port map (
            O => \N__47511\,
            I => n12526
        );

    \I__10431\ : InMux
    port map (
            O => \N__47508\,
            I => n12550
        );

    \I__10430\ : InMux
    port map (
            O => \N__47505\,
            I => n12551
        );

    \I__10429\ : InMux
    port map (
            O => \N__47502\,
            I => \N__47499\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__47499\,
            I => \N__47496\
        );

    \I__10427\ : Span4Mux_h
    port map (
            O => \N__47496\,
            I => \N__47493\
        );

    \I__10426\ : Span4Mux_h
    port map (
            O => \N__47493\,
            I => \N__47490\
        );

    \I__10425\ : Span4Mux_v
    port map (
            O => \N__47490\,
            I => \N__47486\
        );

    \I__10424\ : InMux
    port map (
            O => \N__47489\,
            I => \N__47483\
        );

    \I__10423\ : Odrv4
    port map (
            O => \N__47486\,
            I => n15553
        );

    \I__10422\ : LocalMux
    port map (
            O => \N__47483\,
            I => n15553
        );

    \I__10421\ : CascadeMux
    port map (
            O => \N__47478\,
            I => \N__47475\
        );

    \I__10420\ : InMux
    port map (
            O => \N__47475\,
            I => \N__47472\
        );

    \I__10419\ : LocalMux
    port map (
            O => \N__47472\,
            I => n1401
        );

    \I__10418\ : InMux
    port map (
            O => \N__47469\,
            I => \N__47466\
        );

    \I__10417\ : LocalMux
    port map (
            O => \N__47466\,
            I => n12019
        );

    \I__10416\ : CascadeMux
    port map (
            O => \N__47463\,
            I => \n14406_cascade_\
        );

    \I__10415\ : InMux
    port map (
            O => \N__47460\,
            I => \N__47457\
        );

    \I__10414\ : LocalMux
    port map (
            O => \N__47457\,
            I => n14464
        );

    \I__10413\ : InMux
    port map (
            O => \N__47454\,
            I => n12542
        );

    \I__10412\ : InMux
    port map (
            O => \N__47451\,
            I => n12543
        );

    \I__10411\ : InMux
    port map (
            O => \N__47448\,
            I => n12544
        );

    \I__10410\ : InMux
    port map (
            O => \N__47445\,
            I => \N__47442\
        );

    \I__10409\ : LocalMux
    port map (
            O => \N__47442\,
            I => n1396
        );

    \I__10408\ : InMux
    port map (
            O => \N__47439\,
            I => n12545
        );

    \I__10407\ : InMux
    port map (
            O => \N__47436\,
            I => \N__47433\
        );

    \I__10406\ : LocalMux
    port map (
            O => \N__47433\,
            I => n1395
        );

    \I__10405\ : InMux
    port map (
            O => \N__47430\,
            I => n12546
        );

    \I__10404\ : InMux
    port map (
            O => \N__47427\,
            I => n12547
        );

    \I__10403\ : InMux
    port map (
            O => \N__47424\,
            I => \bfn_14_21_0_\
        );

    \I__10402\ : InMux
    port map (
            O => \N__47421\,
            I => \N__47418\
        );

    \I__10401\ : LocalMux
    port map (
            O => \N__47418\,
            I => \N__47415\
        );

    \I__10400\ : Odrv4
    port map (
            O => \N__47415\,
            I => n1392
        );

    \I__10399\ : InMux
    port map (
            O => \N__47412\,
            I => n12549
        );

    \I__10398\ : CascadeMux
    port map (
            O => \N__47409\,
            I => \n1427_cascade_\
        );

    \I__10397\ : InMux
    port map (
            O => \N__47406\,
            I => \N__47402\
        );

    \I__10396\ : InMux
    port map (
            O => \N__47405\,
            I => \N__47398\
        );

    \I__10395\ : LocalMux
    port map (
            O => \N__47402\,
            I => \N__47395\
        );

    \I__10394\ : InMux
    port map (
            O => \N__47401\,
            I => \N__47392\
        );

    \I__10393\ : LocalMux
    port map (
            O => \N__47398\,
            I => n1628_adj_608
        );

    \I__10392\ : Odrv4
    port map (
            O => \N__47395\,
            I => n1628_adj_608
        );

    \I__10391\ : LocalMux
    port map (
            O => \N__47392\,
            I => n1628_adj_608
        );

    \I__10390\ : InMux
    port map (
            O => \N__47385\,
            I => \N__47382\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__47382\,
            I => \N__47379\
        );

    \I__10388\ : Span4Mux_v
    port map (
            O => \N__47379\,
            I => \N__47376\
        );

    \I__10387\ : Span4Mux_h
    port map (
            O => \N__47376\,
            I => \N__47373\
        );

    \I__10386\ : Odrv4
    port map (
            O => \N__47373\,
            I => n11
        );

    \I__10385\ : InMux
    port map (
            O => \N__47370\,
            I => \N__47366\
        );

    \I__10384\ : CascadeMux
    port map (
            O => \N__47369\,
            I => \N__47362\
        );

    \I__10383\ : LocalMux
    port map (
            O => \N__47366\,
            I => \N__47359\
        );

    \I__10382\ : InMux
    port map (
            O => \N__47365\,
            I => \N__47356\
        );

    \I__10381\ : InMux
    port map (
            O => \N__47362\,
            I => \N__47353\
        );

    \I__10380\ : Span4Mux_h
    port map (
            O => \N__47359\,
            I => \N__47350\
        );

    \I__10379\ : LocalMux
    port map (
            O => \N__47356\,
            I => \N__47347\
        );

    \I__10378\ : LocalMux
    port map (
            O => \N__47353\,
            I => encoder0_position_22
        );

    \I__10377\ : Odrv4
    port map (
            O => \N__47350\,
            I => encoder0_position_22
        );

    \I__10376\ : Odrv12
    port map (
            O => \N__47347\,
            I => encoder0_position_22
        );

    \I__10375\ : CascadeMux
    port map (
            O => \N__47340\,
            I => \N__47337\
        );

    \I__10374\ : InMux
    port map (
            O => \N__47337\,
            I => \N__47332\
        );

    \I__10373\ : InMux
    port map (
            O => \N__47336\,
            I => \N__47327\
        );

    \I__10372\ : InMux
    port map (
            O => \N__47335\,
            I => \N__47327\
        );

    \I__10371\ : LocalMux
    port map (
            O => \N__47332\,
            I => n1626_adj_606
        );

    \I__10370\ : LocalMux
    port map (
            O => \N__47327\,
            I => n1626_adj_606
        );

    \I__10369\ : InMux
    port map (
            O => \N__47322\,
            I => \N__47318\
        );

    \I__10368\ : InMux
    port map (
            O => \N__47321\,
            I => \N__47315\
        );

    \I__10367\ : LocalMux
    port map (
            O => \N__47318\,
            I => \N__47312\
        );

    \I__10366\ : LocalMux
    port map (
            O => \N__47315\,
            I => \N__47309\
        );

    \I__10365\ : Span12Mux_h
    port map (
            O => \N__47312\,
            I => \N__47306\
        );

    \I__10364\ : Odrv4
    port map (
            O => \N__47309\,
            I => duty_6
        );

    \I__10363\ : Odrv12
    port map (
            O => \N__47306\,
            I => duty_6
        );

    \I__10362\ : InMux
    port map (
            O => \N__47301\,
            I => \N__47298\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__47298\,
            I => \N__47295\
        );

    \I__10360\ : Span12Mux_h
    port map (
            O => \N__47295\,
            I => \N__47292\
        );

    \I__10359\ : Odrv12
    port map (
            O => \N__47292\,
            I => n19_adj_591
        );

    \I__10358\ : InMux
    port map (
            O => \N__47289\,
            I => \bfn_14_20_0_\
        );

    \I__10357\ : InMux
    port map (
            O => \N__47286\,
            I => n12541
        );

    \I__10356\ : CascadeMux
    port map (
            O => \N__47283\,
            I => \N__47280\
        );

    \I__10355\ : InMux
    port map (
            O => \N__47280\,
            I => \N__47277\
        );

    \I__10354\ : LocalMux
    port map (
            O => \N__47277\,
            I => \N__47273\
        );

    \I__10353\ : CascadeMux
    port map (
            O => \N__47276\,
            I => \N__47270\
        );

    \I__10352\ : Span4Mux_h
    port map (
            O => \N__47273\,
            I => \N__47267\
        );

    \I__10351\ : InMux
    port map (
            O => \N__47270\,
            I => \N__47264\
        );

    \I__10350\ : Odrv4
    port map (
            O => \N__47267\,
            I => n1624_adj_604
        );

    \I__10349\ : LocalMux
    port map (
            O => \N__47264\,
            I => n1624_adj_604
        );

    \I__10348\ : InMux
    port map (
            O => \N__47259\,
            I => \N__47256\
        );

    \I__10347\ : LocalMux
    port map (
            O => \N__47256\,
            I => n14502
        );

    \I__10346\ : InMux
    port map (
            O => \N__47253\,
            I => \N__47250\
        );

    \I__10345\ : LocalMux
    port map (
            O => \N__47250\,
            I => \N__47247\
        );

    \I__10344\ : Span4Mux_h
    port map (
            O => \N__47247\,
            I => \N__47242\
        );

    \I__10343\ : InMux
    port map (
            O => \N__47246\,
            I => \N__47239\
        );

    \I__10342\ : InMux
    port map (
            O => \N__47245\,
            I => \N__47236\
        );

    \I__10341\ : Odrv4
    port map (
            O => \N__47242\,
            I => n1623_adj_603
        );

    \I__10340\ : LocalMux
    port map (
            O => \N__47239\,
            I => n1623_adj_603
        );

    \I__10339\ : LocalMux
    port map (
            O => \N__47236\,
            I => n1623_adj_603
        );

    \I__10338\ : CascadeMux
    port map (
            O => \N__47229\,
            I => \n1624_adj_604_cascade_\
        );

    \I__10337\ : InMux
    port map (
            O => \N__47226\,
            I => \N__47223\
        );

    \I__10336\ : LocalMux
    port map (
            O => \N__47223\,
            I => n13748
        );

    \I__10335\ : CascadeMux
    port map (
            O => \N__47220\,
            I => \N__47217\
        );

    \I__10334\ : InMux
    port map (
            O => \N__47217\,
            I => \N__47214\
        );

    \I__10333\ : LocalMux
    port map (
            O => \N__47214\,
            I => n14508
        );

    \I__10332\ : CascadeMux
    port map (
            O => \N__47211\,
            I => \N__47208\
        );

    \I__10331\ : InMux
    port map (
            O => \N__47208\,
            I => \N__47204\
        );

    \I__10330\ : CascadeMux
    port map (
            O => \N__47207\,
            I => \N__47201\
        );

    \I__10329\ : LocalMux
    port map (
            O => \N__47204\,
            I => \N__47197\
        );

    \I__10328\ : InMux
    port map (
            O => \N__47201\,
            I => \N__47194\
        );

    \I__10327\ : InMux
    port map (
            O => \N__47200\,
            I => \N__47191\
        );

    \I__10326\ : Odrv4
    port map (
            O => \N__47197\,
            I => n1627_adj_607
        );

    \I__10325\ : LocalMux
    port map (
            O => \N__47194\,
            I => n1627_adj_607
        );

    \I__10324\ : LocalMux
    port map (
            O => \N__47191\,
            I => n1627_adj_607
        );

    \I__10323\ : CascadeMux
    port map (
            O => \N__47184\,
            I => \n1523_cascade_\
        );

    \I__10322\ : InMux
    port map (
            O => \N__47181\,
            I => \N__47177\
        );

    \I__10321\ : CascadeMux
    port map (
            O => \N__47180\,
            I => \N__47174\
        );

    \I__10320\ : LocalMux
    port map (
            O => \N__47177\,
            I => \N__47170\
        );

    \I__10319\ : InMux
    port map (
            O => \N__47174\,
            I => \N__47167\
        );

    \I__10318\ : InMux
    port map (
            O => \N__47173\,
            I => \N__47164\
        );

    \I__10317\ : Odrv4
    port map (
            O => \N__47170\,
            I => n1622_adj_602
        );

    \I__10316\ : LocalMux
    port map (
            O => \N__47167\,
            I => n1622_adj_602
        );

    \I__10315\ : LocalMux
    port map (
            O => \N__47164\,
            I => n1622_adj_602
        );

    \I__10314\ : InMux
    port map (
            O => \N__47157\,
            I => \N__47154\
        );

    \I__10313\ : LocalMux
    port map (
            O => \N__47154\,
            I => n14426
        );

    \I__10312\ : CascadeMux
    port map (
            O => \N__47151\,
            I => \n14428_cascade_\
        );

    \I__10311\ : CascadeMux
    port map (
            O => \N__47148\,
            I => \n1554_cascade_\
        );

    \I__10310\ : CascadeMux
    port map (
            O => \N__47145\,
            I => \N__47141\
        );

    \I__10309\ : InMux
    port map (
            O => \N__47144\,
            I => \N__47138\
        );

    \I__10308\ : InMux
    port map (
            O => \N__47141\,
            I => \N__47135\
        );

    \I__10307\ : LocalMux
    port map (
            O => \N__47138\,
            I => \N__47132\
        );

    \I__10306\ : LocalMux
    port map (
            O => \N__47135\,
            I => \N__47129\
        );

    \I__10305\ : Span4Mux_h
    port map (
            O => \N__47132\,
            I => \N__47126\
        );

    \I__10304\ : Span4Mux_h
    port map (
            O => \N__47129\,
            I => \N__47123\
        );

    \I__10303\ : Odrv4
    port map (
            O => \N__47126\,
            I => n21_adj_667
        );

    \I__10302\ : Odrv4
    port map (
            O => \N__47123\,
            I => n21_adj_667
        );

    \I__10301\ : InMux
    port map (
            O => \N__47118\,
            I => \N__47112\
        );

    \I__10300\ : InMux
    port map (
            O => \N__47117\,
            I => \N__47112\
        );

    \I__10299\ : LocalMux
    port map (
            O => \N__47112\,
            I => \N__47109\
        );

    \I__10298\ : Odrv4
    port map (
            O => \N__47109\,
            I => pwm_setpoint_10
        );

    \I__10297\ : CascadeMux
    port map (
            O => \N__47106\,
            I => \n21_adj_667_cascade_\
        );

    \I__10296\ : InMux
    port map (
            O => \N__47103\,
            I => \N__47100\
        );

    \I__10295\ : LocalMux
    port map (
            O => \N__47100\,
            I => \N__47097\
        );

    \I__10294\ : Odrv12
    port map (
            O => \N__47097\,
            I => n6_adj_656
        );

    \I__10293\ : InMux
    port map (
            O => \N__47094\,
            I => \N__47091\
        );

    \I__10292\ : LocalMux
    port map (
            O => \N__47091\,
            I => \N__47088\
        );

    \I__10291\ : Odrv4
    port map (
            O => \N__47088\,
            I => n15203
        );

    \I__10290\ : CascadeMux
    port map (
            O => \N__47085\,
            I => \n14420_cascade_\
        );

    \I__10289\ : InMux
    port map (
            O => \N__47082\,
            I => \N__47078\
        );

    \I__10288\ : CascadeMux
    port map (
            O => \N__47081\,
            I => \N__47075\
        );

    \I__10287\ : LocalMux
    port map (
            O => \N__47078\,
            I => \N__47072\
        );

    \I__10286\ : InMux
    port map (
            O => \N__47075\,
            I => \N__47069\
        );

    \I__10285\ : Odrv4
    port map (
            O => \N__47072\,
            I => n1630_adj_610
        );

    \I__10284\ : LocalMux
    port map (
            O => \N__47069\,
            I => n1630_adj_610
        );

    \I__10283\ : InMux
    port map (
            O => \N__47064\,
            I => \N__47060\
        );

    \I__10282\ : CascadeMux
    port map (
            O => \N__47063\,
            I => \N__47057\
        );

    \I__10281\ : LocalMux
    port map (
            O => \N__47060\,
            I => \N__47053\
        );

    \I__10280\ : InMux
    port map (
            O => \N__47057\,
            I => \N__47050\
        );

    \I__10279\ : InMux
    port map (
            O => \N__47056\,
            I => \N__47047\
        );

    \I__10278\ : Odrv4
    port map (
            O => \N__47053\,
            I => n1629_adj_609
        );

    \I__10277\ : LocalMux
    port map (
            O => \N__47050\,
            I => n1629_adj_609
        );

    \I__10276\ : LocalMux
    port map (
            O => \N__47047\,
            I => n1629_adj_609
        );

    \I__10275\ : CascadeMux
    port map (
            O => \N__47040\,
            I => \n1630_adj_610_cascade_\
        );

    \I__10274\ : InMux
    port map (
            O => \N__47037\,
            I => \N__47034\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__47034\,
            I => \PWM.n17\
        );

    \I__10272\ : CascadeMux
    port map (
            O => \N__47031\,
            I => \PWM.n26_cascade_\
        );

    \I__10271\ : InMux
    port map (
            O => \N__47028\,
            I => \N__47025\
        );

    \I__10270\ : LocalMux
    port map (
            O => \N__47025\,
            I => \PWM.n27\
        );

    \I__10269\ : CascadeMux
    port map (
            O => \N__47022\,
            I => \PWM.n29_cascade_\
        );

    \I__10268\ : InMux
    port map (
            O => \N__47019\,
            I => \N__47016\
        );

    \I__10267\ : LocalMux
    port map (
            O => \N__47016\,
            I => \PWM.n28\
        );

    \I__10266\ : InMux
    port map (
            O => \N__47013\,
            I => \N__47010\
        );

    \I__10265\ : LocalMux
    port map (
            O => \N__47010\,
            I => commutation_state_prev_2
        );

    \I__10264\ : InMux
    port map (
            O => \N__47007\,
            I => \N__47001\
        );

    \I__10263\ : InMux
    port map (
            O => \N__47006\,
            I => \N__46997\
        );

    \I__10262\ : InMux
    port map (
            O => \N__47005\,
            I => \N__46992\
        );

    \I__10261\ : InMux
    port map (
            O => \N__47004\,
            I => \N__46992\
        );

    \I__10260\ : LocalMux
    port map (
            O => \N__47001\,
            I => \N__46989\
        );

    \I__10259\ : InMux
    port map (
            O => \N__47000\,
            I => \N__46985\
        );

    \I__10258\ : LocalMux
    port map (
            O => \N__46997\,
            I => \N__46980\
        );

    \I__10257\ : LocalMux
    port map (
            O => \N__46992\,
            I => \N__46980\
        );

    \I__10256\ : Span4Mux_h
    port map (
            O => \N__46989\,
            I => \N__46977\
        );

    \I__10255\ : InMux
    port map (
            O => \N__46988\,
            I => \N__46974\
        );

    \I__10254\ : LocalMux
    port map (
            O => \N__46985\,
            I => \N__46971\
        );

    \I__10253\ : Span4Mux_h
    port map (
            O => \N__46980\,
            I => \N__46968\
        );

    \I__10252\ : Odrv4
    port map (
            O => \N__46977\,
            I => h2
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__46974\,
            I => h2
        );

    \I__10250\ : Odrv4
    port map (
            O => \N__46971\,
            I => h2
        );

    \I__10249\ : Odrv4
    port map (
            O => \N__46968\,
            I => h2
        );

    \I__10248\ : InMux
    port map (
            O => \N__46959\,
            I => \N__46952\
        );

    \I__10247\ : InMux
    port map (
            O => \N__46958\,
            I => \N__46949\
        );

    \I__10246\ : InMux
    port map (
            O => \N__46957\,
            I => \N__46944\
        );

    \I__10245\ : InMux
    port map (
            O => \N__46956\,
            I => \N__46944\
        );

    \I__10244\ : InMux
    port map (
            O => \N__46955\,
            I => \N__46941\
        );

    \I__10243\ : LocalMux
    port map (
            O => \N__46952\,
            I => \N__46934\
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__46949\,
            I => \N__46934\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__46944\,
            I => \N__46934\
        );

    \I__10240\ : LocalMux
    port map (
            O => \N__46941\,
            I => \N__46931\
        );

    \I__10239\ : Sp12to4
    port map (
            O => \N__46934\,
            I => \N__46928\
        );

    \I__10238\ : Sp12to4
    port map (
            O => \N__46931\,
            I => \N__46924\
        );

    \I__10237\ : Span12Mux_s10_v
    port map (
            O => \N__46928\,
            I => \N__46921\
        );

    \I__10236\ : InMux
    port map (
            O => \N__46927\,
            I => \N__46918\
        );

    \I__10235\ : Span12Mux_s6_v
    port map (
            O => \N__46924\,
            I => \N__46915\
        );

    \I__10234\ : Span12Mux_h
    port map (
            O => \N__46921\,
            I => \N__46912\
        );

    \I__10233\ : LocalMux
    port map (
            O => \N__46918\,
            I => h3
        );

    \I__10232\ : Odrv12
    port map (
            O => \N__46915\,
            I => h3
        );

    \I__10231\ : Odrv12
    port map (
            O => \N__46912\,
            I => h3
        );

    \I__10230\ : CascadeMux
    port map (
            O => \N__46905\,
            I => \N__46900\
        );

    \I__10229\ : CascadeMux
    port map (
            O => \N__46904\,
            I => \N__46896\
        );

    \I__10228\ : InMux
    port map (
            O => \N__46903\,
            I => \N__46893\
        );

    \I__10227\ : InMux
    port map (
            O => \N__46900\,
            I => \N__46887\
        );

    \I__10226\ : InMux
    port map (
            O => \N__46899\,
            I => \N__46887\
        );

    \I__10225\ : InMux
    port map (
            O => \N__46896\,
            I => \N__46884\
        );

    \I__10224\ : LocalMux
    port map (
            O => \N__46893\,
            I => \N__46881\
        );

    \I__10223\ : InMux
    port map (
            O => \N__46892\,
            I => \N__46878\
        );

    \I__10222\ : LocalMux
    port map (
            O => \N__46887\,
            I => \N__46875\
        );

    \I__10221\ : LocalMux
    port map (
            O => \N__46884\,
            I => \N__46870\
        );

    \I__10220\ : Span4Mux_s2_v
    port map (
            O => \N__46881\,
            I => \N__46870\
        );

    \I__10219\ : LocalMux
    port map (
            O => \N__46878\,
            I => \N__46867\
        );

    \I__10218\ : Span4Mux_s2_v
    port map (
            O => \N__46875\,
            I => \N__46863\
        );

    \I__10217\ : Span4Mux_h
    port map (
            O => \N__46870\,
            I => \N__46858\
        );

    \I__10216\ : Span4Mux_s2_v
    port map (
            O => \N__46867\,
            I => \N__46858\
        );

    \I__10215\ : InMux
    port map (
            O => \N__46866\,
            I => \N__46855\
        );

    \I__10214\ : Sp12to4
    port map (
            O => \N__46863\,
            I => \N__46850\
        );

    \I__10213\ : Sp12to4
    port map (
            O => \N__46858\,
            I => \N__46850\
        );

    \I__10212\ : LocalMux
    port map (
            O => \N__46855\,
            I => h1
        );

    \I__10211\ : Odrv12
    port map (
            O => \N__46850\,
            I => h1
        );

    \I__10210\ : CEMux
    port map (
            O => \N__46845\,
            I => \N__46842\
        );

    \I__10209\ : LocalMux
    port map (
            O => \N__46842\,
            I => \N__46839\
        );

    \I__10208\ : Odrv12
    port map (
            O => \N__46839\,
            I => n6_adj_721
        );

    \I__10207\ : SRMux
    port map (
            O => \N__46836\,
            I => \N__46833\
        );

    \I__10206\ : LocalMux
    port map (
            O => \N__46833\,
            I => \commutation_state_7__N_261\
        );

    \I__10205\ : InMux
    port map (
            O => \N__46830\,
            I => \N__46826\
        );

    \I__10204\ : InMux
    port map (
            O => \N__46829\,
            I => \N__46823\
        );

    \I__10203\ : LocalMux
    port map (
            O => \N__46826\,
            I => \N__46818\
        );

    \I__10202\ : LocalMux
    port map (
            O => \N__46823\,
            I => \N__46818\
        );

    \I__10201\ : Span4Mux_s2_v
    port map (
            O => \N__46818\,
            I => \N__46815\
        );

    \I__10200\ : Span4Mux_v
    port map (
            O => \N__46815\,
            I => \N__46812\
        );

    \I__10199\ : Odrv4
    port map (
            O => \N__46812\,
            I => pwm_setpoint_5
        );

    \I__10198\ : InMux
    port map (
            O => \N__46809\,
            I => \N__46806\
        );

    \I__10197\ : LocalMux
    port map (
            O => \N__46806\,
            I => \N__46802\
        );

    \I__10196\ : CascadeMux
    port map (
            O => \N__46805\,
            I => \N__46799\
        );

    \I__10195\ : Span4Mux_v
    port map (
            O => \N__46802\,
            I => \N__46796\
        );

    \I__10194\ : InMux
    port map (
            O => \N__46799\,
            I => \N__46793\
        );

    \I__10193\ : Odrv4
    port map (
            O => \N__46796\,
            I => n11_adj_660
        );

    \I__10192\ : LocalMux
    port map (
            O => \N__46793\,
            I => n11_adj_660
        );

    \I__10191\ : InMux
    port map (
            O => \N__46788\,
            I => \N__46785\
        );

    \I__10190\ : LocalMux
    port map (
            O => \N__46785\,
            I => \N__46781\
        );

    \I__10189\ : InMux
    port map (
            O => \N__46784\,
            I => \N__46778\
        );

    \I__10188\ : Span4Mux_s2_v
    port map (
            O => \N__46781\,
            I => \N__46775\
        );

    \I__10187\ : LocalMux
    port map (
            O => \N__46778\,
            I => pwm_setpoint_14
        );

    \I__10186\ : Odrv4
    port map (
            O => \N__46775\,
            I => pwm_setpoint_14
        );

    \I__10185\ : CascadeMux
    port map (
            O => \N__46770\,
            I => \N__46767\
        );

    \I__10184\ : InMux
    port map (
            O => \N__46767\,
            I => \N__46760\
        );

    \I__10183\ : InMux
    port map (
            O => \N__46766\,
            I => \N__46760\
        );

    \I__10182\ : InMux
    port map (
            O => \N__46765\,
            I => \N__46757\
        );

    \I__10181\ : LocalMux
    port map (
            O => \N__46760\,
            I => n29_adj_672
        );

    \I__10180\ : LocalMux
    port map (
            O => \N__46757\,
            I => n29_adj_672
        );

    \I__10179\ : CascadeMux
    port map (
            O => \N__46752\,
            I => \N__46749\
        );

    \I__10178\ : InMux
    port map (
            O => \N__46749\,
            I => \N__46745\
        );

    \I__10177\ : InMux
    port map (
            O => \N__46748\,
            I => \N__46742\
        );

    \I__10176\ : LocalMux
    port map (
            O => \N__46745\,
            I => duty_19
        );

    \I__10175\ : LocalMux
    port map (
            O => \N__46742\,
            I => duty_19
        );

    \I__10174\ : InMux
    port map (
            O => \N__46737\,
            I => \N__46734\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__46734\,
            I => \N__46731\
        );

    \I__10172\ : Odrv4
    port map (
            O => \N__46731\,
            I => n6_adj_578
        );

    \I__10171\ : InMux
    port map (
            O => \N__46728\,
            I => \N__46725\
        );

    \I__10170\ : LocalMux
    port map (
            O => \N__46725\,
            I => \PWM.n13991\
        );

    \I__10169\ : CascadeMux
    port map (
            O => \N__46722\,
            I => \N__46715\
        );

    \I__10168\ : CascadeMux
    port map (
            O => \N__46721\,
            I => \N__46712\
        );

    \I__10167\ : InMux
    port map (
            O => \N__46720\,
            I => \N__46699\
        );

    \I__10166\ : InMux
    port map (
            O => \N__46719\,
            I => \N__46699\
        );

    \I__10165\ : InMux
    port map (
            O => \N__46718\,
            I => \N__46699\
        );

    \I__10164\ : InMux
    port map (
            O => \N__46715\,
            I => \N__46699\
        );

    \I__10163\ : InMux
    port map (
            O => \N__46712\,
            I => \N__46699\
        );

    \I__10162\ : InMux
    port map (
            O => \N__46711\,
            I => \N__46694\
        );

    \I__10161\ : InMux
    port map (
            O => \N__46710\,
            I => \N__46694\
        );

    \I__10160\ : LocalMux
    port map (
            O => \N__46699\,
            I => \N__46687\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__46694\,
            I => \N__46687\
        );

    \I__10158\ : InMux
    port map (
            O => \N__46693\,
            I => \N__46682\
        );

    \I__10157\ : InMux
    port map (
            O => \N__46692\,
            I => \N__46682\
        );

    \I__10156\ : Span4Mux_v
    port map (
            O => \N__46687\,
            I => \N__46677\
        );

    \I__10155\ : LocalMux
    port map (
            O => \N__46682\,
            I => \N__46677\
        );

    \I__10154\ : Span4Mux_h
    port map (
            O => \N__46677\,
            I => \N__46674\
        );

    \I__10153\ : Odrv4
    port map (
            O => \N__46674\,
            I => n4_adj_599
        );

    \I__10152\ : InMux
    port map (
            O => \N__46671\,
            I => \N__46668\
        );

    \I__10151\ : LocalMux
    port map (
            O => \N__46668\,
            I => commutation_state_prev_1
        );

    \I__10150\ : InMux
    port map (
            O => \N__46665\,
            I => \N__46661\
        );

    \I__10149\ : InMux
    port map (
            O => \N__46664\,
            I => \N__46655\
        );

    \I__10148\ : LocalMux
    port map (
            O => \N__46661\,
            I => \N__46652\
        );

    \I__10147\ : InMux
    port map (
            O => \N__46660\,
            I => \N__46649\
        );

    \I__10146\ : InMux
    port map (
            O => \N__46659\,
            I => \N__46644\
        );

    \I__10145\ : InMux
    port map (
            O => \N__46658\,
            I => \N__46644\
        );

    \I__10144\ : LocalMux
    port map (
            O => \N__46655\,
            I => \N__46641\
        );

    \I__10143\ : Span4Mux_v
    port map (
            O => \N__46652\,
            I => \N__46638\
        );

    \I__10142\ : LocalMux
    port map (
            O => \N__46649\,
            I => \N__46633\
        );

    \I__10141\ : LocalMux
    port map (
            O => \N__46644\,
            I => \N__46633\
        );

    \I__10140\ : Span4Mux_v
    port map (
            O => \N__46641\,
            I => \N__46630\
        );

    \I__10139\ : Odrv4
    port map (
            O => \N__46638\,
            I => n5137
        );

    \I__10138\ : Odrv4
    port map (
            O => \N__46633\,
            I => n5137
        );

    \I__10137\ : Odrv4
    port map (
            O => \N__46630\,
            I => n5137
        );

    \I__10136\ : InMux
    port map (
            O => \N__46623\,
            I => \N__46617\
        );

    \I__10135\ : InMux
    port map (
            O => \N__46622\,
            I => \N__46617\
        );

    \I__10134\ : LocalMux
    port map (
            O => \N__46617\,
            I => \N__46611\
        );

    \I__10133\ : InMux
    port map (
            O => \N__46616\,
            I => \N__46608\
        );

    \I__10132\ : InMux
    port map (
            O => \N__46615\,
            I => \N__46605\
        );

    \I__10131\ : InMux
    port map (
            O => \N__46614\,
            I => \N__46602\
        );

    \I__10130\ : Span4Mux_v
    port map (
            O => \N__46611\,
            I => \N__46598\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__46608\,
            I => \N__46591\
        );

    \I__10128\ : LocalMux
    port map (
            O => \N__46605\,
            I => \N__46591\
        );

    \I__10127\ : LocalMux
    port map (
            O => \N__46602\,
            I => \N__46591\
        );

    \I__10126\ : InMux
    port map (
            O => \N__46601\,
            I => \N__46588\
        );

    \I__10125\ : Span4Mux_v
    port map (
            O => \N__46598\,
            I => \N__46583\
        );

    \I__10124\ : Span4Mux_v
    port map (
            O => \N__46591\,
            I => \N__46583\
        );

    \I__10123\ : LocalMux
    port map (
            O => \N__46588\,
            I => dti
        );

    \I__10122\ : Odrv4
    port map (
            O => \N__46583\,
            I => dti
        );

    \I__10121\ : CascadeMux
    port map (
            O => \N__46578\,
            I => \n5201_cascade_\
        );

    \I__10120\ : InMux
    port map (
            O => \N__46575\,
            I => \N__46572\
        );

    \I__10119\ : LocalMux
    port map (
            O => \N__46572\,
            I => \N__46568\
        );

    \I__10118\ : InMux
    port map (
            O => \N__46571\,
            I => \N__46565\
        );

    \I__10117\ : Span4Mux_v
    port map (
            O => \N__46568\,
            I => \N__46562\
        );

    \I__10116\ : LocalMux
    port map (
            O => \N__46565\,
            I => \N__46559\
        );

    \I__10115\ : Sp12to4
    port map (
            O => \N__46562\,
            I => \N__46556\
        );

    \I__10114\ : Span4Mux_h
    port map (
            O => \N__46559\,
            I => \N__46553\
        );

    \I__10113\ : Odrv12
    port map (
            O => \N__46556\,
            I => pwm_setpoint_13
        );

    \I__10112\ : Odrv4
    port map (
            O => \N__46553\,
            I => pwm_setpoint_13
        );

    \I__10111\ : InMux
    port map (
            O => \N__46548\,
            I => \N__46544\
        );

    \I__10110\ : InMux
    port map (
            O => \N__46547\,
            I => \N__46541\
        );

    \I__10109\ : LocalMux
    port map (
            O => \N__46544\,
            I => \N__46535\
        );

    \I__10108\ : LocalMux
    port map (
            O => \N__46541\,
            I => \N__46535\
        );

    \I__10107\ : InMux
    port map (
            O => \N__46540\,
            I => \N__46532\
        );

    \I__10106\ : Odrv4
    port map (
            O => \N__46535\,
            I => n27_adj_671
        );

    \I__10105\ : LocalMux
    port map (
            O => \N__46532\,
            I => n27_adj_671
        );

    \I__10104\ : InMux
    port map (
            O => \N__46527\,
            I => \N__46523\
        );

    \I__10103\ : InMux
    port map (
            O => \N__46526\,
            I => \N__46520\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__46523\,
            I => \N__46517\
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__46520\,
            I => duty_2
        );

    \I__10100\ : Odrv4
    port map (
            O => \N__46517\,
            I => duty_2
        );

    \I__10099\ : InMux
    port map (
            O => \N__46512\,
            I => \N__46509\
        );

    \I__10098\ : LocalMux
    port map (
            O => \N__46509\,
            I => \N__46506\
        );

    \I__10097\ : Span4Mux_v
    port map (
            O => \N__46506\,
            I => \N__46503\
        );

    \I__10096\ : Odrv4
    port map (
            O => \N__46503\,
            I => n23_adj_595
        );

    \I__10095\ : InMux
    port map (
            O => \N__46500\,
            I => \N__46496\
        );

    \I__10094\ : InMux
    port map (
            O => \N__46499\,
            I => \N__46493\
        );

    \I__10093\ : LocalMux
    port map (
            O => \N__46496\,
            I => \N__46490\
        );

    \I__10092\ : LocalMux
    port map (
            O => \N__46493\,
            I => duty_15
        );

    \I__10091\ : Odrv12
    port map (
            O => \N__46490\,
            I => duty_15
        );

    \I__10090\ : InMux
    port map (
            O => \N__46485\,
            I => \N__46482\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__46482\,
            I => \N__46479\
        );

    \I__10088\ : Odrv12
    port map (
            O => \N__46479\,
            I => \pwm_setpoint_23_N_171_15\
        );

    \I__10087\ : InMux
    port map (
            O => \N__46476\,
            I => \N__46470\
        );

    \I__10086\ : InMux
    port map (
            O => \N__46475\,
            I => \N__46470\
        );

    \I__10085\ : LocalMux
    port map (
            O => \N__46470\,
            I => \N__46467\
        );

    \I__10084\ : Span4Mux_s2_v
    port map (
            O => \N__46467\,
            I => \N__46464\
        );

    \I__10083\ : Odrv4
    port map (
            O => \N__46464\,
            I => pwm_setpoint_15
        );

    \I__10082\ : InMux
    port map (
            O => \N__46461\,
            I => \N__46458\
        );

    \I__10081\ : LocalMux
    port map (
            O => \N__46458\,
            I => \N__46453\
        );

    \I__10080\ : InMux
    port map (
            O => \N__46457\,
            I => \N__46450\
        );

    \I__10079\ : InMux
    port map (
            O => \N__46456\,
            I => \N__46447\
        );

    \I__10078\ : Span4Mux_v
    port map (
            O => \N__46453\,
            I => \N__46442\
        );

    \I__10077\ : LocalMux
    port map (
            O => \N__46450\,
            I => \N__46442\
        );

    \I__10076\ : LocalMux
    port map (
            O => \N__46447\,
            I => \N__46439\
        );

    \I__10075\ : Span4Mux_h
    port map (
            O => \N__46442\,
            I => \N__46434\
        );

    \I__10074\ : Span4Mux_h
    port map (
            O => \N__46439\,
            I => \N__46434\
        );

    \I__10073\ : Span4Mux_h
    port map (
            O => \N__46434\,
            I => \N__46431\
        );

    \I__10072\ : Odrv4
    port map (
            O => \N__46431\,
            I => \quad_counter0.a_new_0\
        );

    \I__10071\ : InMux
    port map (
            O => \N__46428\,
            I => \N__46425\
        );

    \I__10070\ : LocalMux
    port map (
            O => \N__46425\,
            I => \N__46421\
        );

    \I__10069\ : InMux
    port map (
            O => \N__46424\,
            I => \N__46418\
        );

    \I__10068\ : Span4Mux_h
    port map (
            O => \N__46421\,
            I => \N__46412\
        );

    \I__10067\ : LocalMux
    port map (
            O => \N__46418\,
            I => \N__46412\
        );

    \I__10066\ : InMux
    port map (
            O => \N__46417\,
            I => \N__46409\
        );

    \I__10065\ : Span4Mux_v
    port map (
            O => \N__46412\,
            I => \N__46406\
        );

    \I__10064\ : LocalMux
    port map (
            O => \N__46409\,
            I => \quad_counter0.b_new_0\
        );

    \I__10063\ : Odrv4
    port map (
            O => \N__46406\,
            I => \quad_counter0.b_new_0\
        );

    \I__10062\ : CascadeMux
    port map (
            O => \N__46401\,
            I => \N__46397\
        );

    \I__10061\ : InMux
    port map (
            O => \N__46400\,
            I => \N__46390\
        );

    \I__10060\ : InMux
    port map (
            O => \N__46397\,
            I => \N__46387\
        );

    \I__10059\ : InMux
    port map (
            O => \N__46396\,
            I => \N__46380\
        );

    \I__10058\ : InMux
    port map (
            O => \N__46395\,
            I => \N__46380\
        );

    \I__10057\ : InMux
    port map (
            O => \N__46394\,
            I => \N__46380\
        );

    \I__10056\ : CascadeMux
    port map (
            O => \N__46393\,
            I => \N__46377\
        );

    \I__10055\ : LocalMux
    port map (
            O => \N__46390\,
            I => \N__46372\
        );

    \I__10054\ : LocalMux
    port map (
            O => \N__46387\,
            I => \N__46372\
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__46380\,
            I => \N__46369\
        );

    \I__10052\ : InMux
    port map (
            O => \N__46377\,
            I => \N__46366\
        );

    \I__10051\ : Span4Mux_v
    port map (
            O => \N__46372\,
            I => \N__46361\
        );

    \I__10050\ : Span4Mux_v
    port map (
            O => \N__46369\,
            I => \N__46361\
        );

    \I__10049\ : LocalMux
    port map (
            O => \N__46366\,
            I => a_new_1
        );

    \I__10048\ : Odrv4
    port map (
            O => \N__46361\,
            I => a_new_1
        );

    \I__10047\ : InMux
    port map (
            O => \N__46356\,
            I => \N__46353\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__46353\,
            I => \N__46350\
        );

    \I__10045\ : Odrv12
    port map (
            O => \N__46350\,
            I => \quad_counter0.a_prev_N_543\
        );

    \I__10044\ : CascadeMux
    port map (
            O => \N__46347\,
            I => \N__46344\
        );

    \I__10043\ : InMux
    port map (
            O => \N__46344\,
            I => \N__46341\
        );

    \I__10042\ : LocalMux
    port map (
            O => \N__46341\,
            I => \N__46337\
        );

    \I__10041\ : InMux
    port map (
            O => \N__46340\,
            I => \N__46334\
        );

    \I__10040\ : Span4Mux_v
    port map (
            O => \N__46337\,
            I => \N__46327\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__46334\,
            I => \N__46327\
        );

    \I__10038\ : InMux
    port map (
            O => \N__46333\,
            I => \N__46322\
        );

    \I__10037\ : InMux
    port map (
            O => \N__46332\,
            I => \N__46322\
        );

    \I__10036\ : Span4Mux_v
    port map (
            O => \N__46327\,
            I => \N__46319\
        );

    \I__10035\ : LocalMux
    port map (
            O => \N__46322\,
            I => \N__46316\
        );

    \I__10034\ : Span4Mux_h
    port map (
            O => \N__46319\,
            I => \N__46313\
        );

    \I__10033\ : Odrv12
    port map (
            O => \N__46316\,
            I => \quad_counter0.b_new_1\
        );

    \I__10032\ : Odrv4
    port map (
            O => \N__46313\,
            I => \quad_counter0.b_new_1\
        );

    \I__10031\ : CascadeMux
    port map (
            O => \N__46308\,
            I => \N__46303\
        );

    \I__10030\ : InMux
    port map (
            O => \N__46307\,
            I => \N__46300\
        );

    \I__10029\ : InMux
    port map (
            O => \N__46306\,
            I => \N__46297\
        );

    \I__10028\ : InMux
    port map (
            O => \N__46303\,
            I => \N__46294\
        );

    \I__10027\ : LocalMux
    port map (
            O => \N__46300\,
            I => \N__46291\
        );

    \I__10026\ : LocalMux
    port map (
            O => \N__46297\,
            I => \N__46288\
        );

    \I__10025\ : LocalMux
    port map (
            O => \N__46294\,
            I => \quad_counter0.debounce_cnt\
        );

    \I__10024\ : Odrv12
    port map (
            O => \N__46291\,
            I => \quad_counter0.debounce_cnt\
        );

    \I__10023\ : Odrv12
    port map (
            O => \N__46288\,
            I => \quad_counter0.debounce_cnt\
        );

    \I__10022\ : CascadeMux
    port map (
            O => \N__46281\,
            I => \quad_counter0.a_prev_N_543_cascade_\
        );

    \I__10021\ : InMux
    port map (
            O => \N__46278\,
            I => \N__46274\
        );

    \I__10020\ : InMux
    port map (
            O => \N__46277\,
            I => \N__46271\
        );

    \I__10019\ : LocalMux
    port map (
            O => \N__46274\,
            I => \N__46266\
        );

    \I__10018\ : LocalMux
    port map (
            O => \N__46271\,
            I => \N__46263\
        );

    \I__10017\ : InMux
    port map (
            O => \N__46270\,
            I => \N__46260\
        );

    \I__10016\ : InMux
    port map (
            O => \N__46269\,
            I => \N__46257\
        );

    \I__10015\ : Span4Mux_h
    port map (
            O => \N__46266\,
            I => \N__46254\
        );

    \I__10014\ : Span4Mux_h
    port map (
            O => \N__46263\,
            I => \N__46251\
        );

    \I__10013\ : LocalMux
    port map (
            O => \N__46260\,
            I => \N__46248\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__46257\,
            I => b_prev
        );

    \I__10011\ : Odrv4
    port map (
            O => \N__46254\,
            I => b_prev
        );

    \I__10010\ : Odrv4
    port map (
            O => \N__46251\,
            I => b_prev
        );

    \I__10009\ : Odrv12
    port map (
            O => \N__46248\,
            I => b_prev
        );

    \I__10008\ : CascadeMux
    port map (
            O => \N__46239\,
            I => \N__46236\
        );

    \I__10007\ : InMux
    port map (
            O => \N__46236\,
            I => \N__46233\
        );

    \I__10006\ : LocalMux
    port map (
            O => \N__46233\,
            I => \N__46230\
        );

    \I__10005\ : Span4Mux_v
    port map (
            O => \N__46230\,
            I => \N__46227\
        );

    \I__10004\ : Odrv4
    port map (
            O => \N__46227\,
            I => n15121
        );

    \I__10003\ : InMux
    port map (
            O => \N__46224\,
            I => \N__46221\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__46221\,
            I => \N__46218\
        );

    \I__10001\ : Span4Mux_h
    port map (
            O => \N__46218\,
            I => \N__46215\
        );

    \I__10000\ : Odrv4
    port map (
            O => \N__46215\,
            I => \pwm_setpoint_23_N_171_6\
        );

    \I__9999\ : InMux
    port map (
            O => \N__46212\,
            I => \N__46209\
        );

    \I__9998\ : LocalMux
    port map (
            O => \N__46209\,
            I => \N__46205\
        );

    \I__9997\ : InMux
    port map (
            O => \N__46208\,
            I => \N__46202\
        );

    \I__9996\ : Odrv4
    port map (
            O => \N__46205\,
            I => pwm_setpoint_6
        );

    \I__9995\ : LocalMux
    port map (
            O => \N__46202\,
            I => pwm_setpoint_6
        );

    \I__9994\ : InMux
    port map (
            O => \N__46197\,
            I => \N__46191\
        );

    \I__9993\ : InMux
    port map (
            O => \N__46196\,
            I => \N__46191\
        );

    \I__9992\ : LocalMux
    port map (
            O => \N__46191\,
            I => \N__46188\
        );

    \I__9991\ : Odrv4
    port map (
            O => \N__46188\,
            I => pwm_setpoint_2
        );

    \I__9990\ : InMux
    port map (
            O => \N__46185\,
            I => \N__46179\
        );

    \I__9989\ : InMux
    port map (
            O => \N__46184\,
            I => \N__46179\
        );

    \I__9988\ : LocalMux
    port map (
            O => \N__46179\,
            I => \N__46176\
        );

    \I__9987\ : Odrv4
    port map (
            O => \N__46176\,
            I => pwm_setpoint_3
        );

    \I__9986\ : CascadeMux
    port map (
            O => \N__46173\,
            I => \n14034_cascade_\
        );

    \I__9985\ : CascadeMux
    port map (
            O => \N__46170\,
            I => \n14116_cascade_\
        );

    \I__9984\ : InMux
    port map (
            O => \N__46167\,
            I => \N__46164\
        );

    \I__9983\ : LocalMux
    port map (
            O => \N__46164\,
            I => n10_adj_598
        );

    \I__9982\ : InMux
    port map (
            O => \N__46161\,
            I => \N__46158\
        );

    \I__9981\ : LocalMux
    port map (
            O => \N__46158\,
            I => \N__46155\
        );

    \I__9980\ : Odrv4
    port map (
            O => \N__46155\,
            I => \pwm_setpoint_23_N_171_2\
        );

    \I__9979\ : InMux
    port map (
            O => \N__46152\,
            I => \N__46149\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__46149\,
            I => \N__46146\
        );

    \I__9977\ : Odrv4
    port map (
            O => \N__46146\,
            I => \pwm_setpoint_23_N_171_3\
        );

    \I__9976\ : InMux
    port map (
            O => \N__46143\,
            I => \N__46139\
        );

    \I__9975\ : InMux
    port map (
            O => \N__46142\,
            I => \N__46136\
        );

    \I__9974\ : LocalMux
    port map (
            O => \N__46139\,
            I => duty_3
        );

    \I__9973\ : LocalMux
    port map (
            O => \N__46136\,
            I => duty_3
        );

    \I__9972\ : CascadeMux
    port map (
            O => \N__46131\,
            I => \N__46128\
        );

    \I__9971\ : InMux
    port map (
            O => \N__46128\,
            I => \N__46125\
        );

    \I__9970\ : LocalMux
    port map (
            O => \N__46125\,
            I => n10_adj_681
        );

    \I__9969\ : CascadeMux
    port map (
            O => \N__46122\,
            I => \n16_adj_710_cascade_\
        );

    \I__9968\ : InMux
    port map (
            O => \N__46119\,
            I => \N__46116\
        );

    \I__9967\ : LocalMux
    port map (
            O => \N__46116\,
            I => \N__46113\
        );

    \I__9966\ : Odrv4
    port map (
            O => \N__46113\,
            I => n15_adj_711
        );

    \I__9965\ : InMux
    port map (
            O => \N__46110\,
            I => n12509
        );

    \I__9964\ : CascadeMux
    port map (
            O => \N__46107\,
            I => \N__46104\
        );

    \I__9963\ : InMux
    port map (
            O => \N__46104\,
            I => \N__46101\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__46101\,
            I => \N__46097\
        );

    \I__9961\ : InMux
    port map (
            O => \N__46100\,
            I => \N__46093\
        );

    \I__9960\ : Span4Mux_v
    port map (
            O => \N__46097\,
            I => \N__46090\
        );

    \I__9959\ : InMux
    port map (
            O => \N__46096\,
            I => \N__46087\
        );

    \I__9958\ : LocalMux
    port map (
            O => \N__46093\,
            I => n930
        );

    \I__9957\ : Odrv4
    port map (
            O => \N__46090\,
            I => n930
        );

    \I__9956\ : LocalMux
    port map (
            O => \N__46087\,
            I => n930
        );

    \I__9955\ : InMux
    port map (
            O => \N__46080\,
            I => \N__46077\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__46077\,
            I => n997
        );

    \I__9953\ : InMux
    port map (
            O => \N__46074\,
            I => n12510
        );

    \I__9952\ : CascadeMux
    port map (
            O => \N__46071\,
            I => \N__46068\
        );

    \I__9951\ : InMux
    port map (
            O => \N__46068\,
            I => \N__46065\
        );

    \I__9950\ : LocalMux
    port map (
            O => \N__46065\,
            I => \N__46061\
        );

    \I__9949\ : InMux
    port map (
            O => \N__46064\,
            I => \N__46058\
        );

    \I__9948\ : Span4Mux_h
    port map (
            O => \N__46061\,
            I => \N__46055\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__46058\,
            I => n929
        );

    \I__9946\ : Odrv4
    port map (
            O => \N__46055\,
            I => n929
        );

    \I__9945\ : InMux
    port map (
            O => \N__46050\,
            I => \N__46047\
        );

    \I__9944\ : LocalMux
    port map (
            O => \N__46047\,
            I => n996
        );

    \I__9943\ : InMux
    port map (
            O => \N__46044\,
            I => n12511
        );

    \I__9942\ : CascadeMux
    port map (
            O => \N__46041\,
            I => \N__46038\
        );

    \I__9941\ : InMux
    port map (
            O => \N__46038\,
            I => \N__46033\
        );

    \I__9940\ : InMux
    port map (
            O => \N__46037\,
            I => \N__46028\
        );

    \I__9939\ : InMux
    port map (
            O => \N__46036\,
            I => \N__46028\
        );

    \I__9938\ : LocalMux
    port map (
            O => \N__46033\,
            I => n928
        );

    \I__9937\ : LocalMux
    port map (
            O => \N__46028\,
            I => n928
        );

    \I__9936\ : InMux
    port map (
            O => \N__46023\,
            I => \N__46020\
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__46020\,
            I => n995
        );

    \I__9934\ : InMux
    port map (
            O => \N__46017\,
            I => n12512
        );

    \I__9933\ : CascadeMux
    port map (
            O => \N__46014\,
            I => \N__46009\
        );

    \I__9932\ : CascadeMux
    port map (
            O => \N__46013\,
            I => \N__46005\
        );

    \I__9931\ : InMux
    port map (
            O => \N__46012\,
            I => \N__45999\
        );

    \I__9930\ : InMux
    port map (
            O => \N__46009\,
            I => \N__45996\
        );

    \I__9929\ : InMux
    port map (
            O => \N__46008\,
            I => \N__45993\
        );

    \I__9928\ : InMux
    port map (
            O => \N__46005\,
            I => \N__45984\
        );

    \I__9927\ : InMux
    port map (
            O => \N__46004\,
            I => \N__45984\
        );

    \I__9926\ : InMux
    port map (
            O => \N__46003\,
            I => \N__45984\
        );

    \I__9925\ : InMux
    port map (
            O => \N__46002\,
            I => \N__45984\
        );

    \I__9924\ : LocalMux
    port map (
            O => \N__45999\,
            I => n960
        );

    \I__9923\ : LocalMux
    port map (
            O => \N__45996\,
            I => n960
        );

    \I__9922\ : LocalMux
    port map (
            O => \N__45993\,
            I => n960
        );

    \I__9921\ : LocalMux
    port map (
            O => \N__45984\,
            I => n960
        );

    \I__9920\ : CascadeMux
    port map (
            O => \N__45975\,
            I => \N__45972\
        );

    \I__9919\ : InMux
    port map (
            O => \N__45972\,
            I => \N__45969\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__45969\,
            I => \N__45965\
        );

    \I__9917\ : InMux
    port map (
            O => \N__45968\,
            I => \N__45962\
        );

    \I__9916\ : Odrv4
    port map (
            O => \N__45965\,
            I => n927
        );

    \I__9915\ : LocalMux
    port map (
            O => \N__45962\,
            I => n927
        );

    \I__9914\ : InMux
    port map (
            O => \N__45957\,
            I => n12513
        );

    \I__9913\ : InMux
    port map (
            O => \N__45954\,
            I => \N__45951\
        );

    \I__9912\ : LocalMux
    port map (
            O => \N__45951\,
            I => \N__45948\
        );

    \I__9911\ : Odrv12
    port map (
            O => \N__45948\,
            I => encoder0_position_scaled_0
        );

    \I__9910\ : InMux
    port map (
            O => \N__45945\,
            I => \N__45942\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__45942\,
            I => n25_adj_551
        );

    \I__9908\ : CascadeMux
    port map (
            O => \N__45939\,
            I => \n11872_cascade_\
        );

    \I__9907\ : CascadeMux
    port map (
            O => \N__45936\,
            I => \n11933_cascade_\
        );

    \I__9906\ : CascadeMux
    port map (
            O => \N__45933\,
            I => \n13728_cascade_\
        );

    \I__9905\ : CascadeMux
    port map (
            O => \N__45930\,
            I => \n1059_cascade_\
        );

    \I__9904\ : CascadeMux
    port map (
            O => \N__45927\,
            I => \n1132_cascade_\
        );

    \I__9903\ : InMux
    port map (
            O => \N__45924\,
            I => \N__45920\
        );

    \I__9902\ : InMux
    port map (
            O => \N__45923\,
            I => \N__45917\
        );

    \I__9901\ : LocalMux
    port map (
            O => \N__45920\,
            I => n295
        );

    \I__9900\ : LocalMux
    port map (
            O => \N__45917\,
            I => n295
        );

    \I__9899\ : InMux
    port map (
            O => \N__45912\,
            I => \N__45909\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__45909\,
            I => n1001
        );

    \I__9897\ : InMux
    port map (
            O => \N__45906\,
            I => \bfn_13_24_0_\
        );

    \I__9896\ : CascadeMux
    port map (
            O => \N__45903\,
            I => \N__45900\
        );

    \I__9895\ : InMux
    port map (
            O => \N__45900\,
            I => \N__45896\
        );

    \I__9894\ : InMux
    port map (
            O => \N__45899\,
            I => \N__45893\
        );

    \I__9893\ : LocalMux
    port map (
            O => \N__45896\,
            I => n933
        );

    \I__9892\ : LocalMux
    port map (
            O => \N__45893\,
            I => n933
        );

    \I__9891\ : InMux
    port map (
            O => \N__45888\,
            I => \N__45885\
        );

    \I__9890\ : LocalMux
    port map (
            O => \N__45885\,
            I => n1000
        );

    \I__9889\ : InMux
    port map (
            O => \N__45882\,
            I => n12507
        );

    \I__9888\ : CascadeMux
    port map (
            O => \N__45879\,
            I => \N__45876\
        );

    \I__9887\ : InMux
    port map (
            O => \N__45876\,
            I => \N__45872\
        );

    \I__9886\ : InMux
    port map (
            O => \N__45875\,
            I => \N__45869\
        );

    \I__9885\ : LocalMux
    port map (
            O => \N__45872\,
            I => n932
        );

    \I__9884\ : LocalMux
    port map (
            O => \N__45869\,
            I => n932
        );

    \I__9883\ : InMux
    port map (
            O => \N__45864\,
            I => \N__45861\
        );

    \I__9882\ : LocalMux
    port map (
            O => \N__45861\,
            I => n999
        );

    \I__9881\ : InMux
    port map (
            O => \N__45858\,
            I => n12508
        );

    \I__9880\ : CascadeMux
    port map (
            O => \N__45855\,
            I => \N__45851\
        );

    \I__9879\ : InMux
    port map (
            O => \N__45854\,
            I => \N__45847\
        );

    \I__9878\ : InMux
    port map (
            O => \N__45851\,
            I => \N__45844\
        );

    \I__9877\ : InMux
    port map (
            O => \N__45850\,
            I => \N__45841\
        );

    \I__9876\ : LocalMux
    port map (
            O => \N__45847\,
            I => n931
        );

    \I__9875\ : LocalMux
    port map (
            O => \N__45844\,
            I => n931
        );

    \I__9874\ : LocalMux
    port map (
            O => \N__45841\,
            I => n931
        );

    \I__9873\ : CascadeMux
    port map (
            O => \N__45834\,
            I => \N__45831\
        );

    \I__9872\ : InMux
    port map (
            O => \N__45831\,
            I => \N__45828\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__45828\,
            I => \N__45825\
        );

    \I__9870\ : Odrv4
    port map (
            O => \N__45825\,
            I => n998
        );

    \I__9869\ : InMux
    port map (
            O => \N__45822\,
            I => \N__45819\
        );

    \I__9868\ : LocalMux
    port map (
            O => \N__45819\,
            I => \N__45816\
        );

    \I__9867\ : Span4Mux_v
    port map (
            O => \N__45816\,
            I => \N__45813\
        );

    \I__9866\ : Span4Mux_h
    port map (
            O => \N__45813\,
            I => \N__45810\
        );

    \I__9865\ : Sp12to4
    port map (
            O => \N__45810\,
            I => \N__45807\
        );

    \I__9864\ : Odrv12
    port map (
            O => \N__45807\,
            I => \ENCODER0_B_N\
        );

    \I__9863\ : InMux
    port map (
            O => \N__45804\,
            I => \N__45801\
        );

    \I__9862\ : LocalMux
    port map (
            O => \N__45801\,
            I => \N__45796\
        );

    \I__9861\ : InMux
    port map (
            O => \N__45800\,
            I => \N__45793\
        );

    \I__9860\ : CascadeMux
    port map (
            O => \N__45799\,
            I => \N__45790\
        );

    \I__9859\ : Span4Mux_h
    port map (
            O => \N__45796\,
            I => \N__45787\
        );

    \I__9858\ : LocalMux
    port map (
            O => \N__45793\,
            I => \N__45784\
        );

    \I__9857\ : InMux
    port map (
            O => \N__45790\,
            I => \N__45781\
        );

    \I__9856\ : Span4Mux_v
    port map (
            O => \N__45787\,
            I => \N__45776\
        );

    \I__9855\ : Span4Mux_v
    port map (
            O => \N__45784\,
            I => \N__45776\
        );

    \I__9854\ : LocalMux
    port map (
            O => \N__45781\,
            I => encoder0_position_1
        );

    \I__9853\ : Odrv4
    port map (
            O => \N__45776\,
            I => encoder0_position_1
        );

    \I__9852\ : CascadeMux
    port map (
            O => \N__45771\,
            I => \N__45768\
        );

    \I__9851\ : InMux
    port map (
            O => \N__45768\,
            I => \N__45765\
        );

    \I__9850\ : LocalMux
    port map (
            O => \N__45765\,
            I => \N__45762\
        );

    \I__9849\ : Odrv12
    port map (
            O => \N__45762\,
            I => n32_adj_650
        );

    \I__9848\ : InMux
    port map (
            O => \N__45759\,
            I => \N__45754\
        );

    \I__9847\ : InMux
    port map (
            O => \N__45758\,
            I => \N__45751\
        );

    \I__9846\ : CascadeMux
    port map (
            O => \N__45757\,
            I => \N__45748\
        );

    \I__9845\ : LocalMux
    port map (
            O => \N__45754\,
            I => \N__45743\
        );

    \I__9844\ : LocalMux
    port map (
            O => \N__45751\,
            I => \N__45743\
        );

    \I__9843\ : InMux
    port map (
            O => \N__45748\,
            I => \N__45740\
        );

    \I__9842\ : Span4Mux_h
    port map (
            O => \N__45743\,
            I => \N__45737\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__45740\,
            I => encoder0_position_16
        );

    \I__9840\ : Odrv4
    port map (
            O => \N__45737\,
            I => encoder0_position_16
        );

    \I__9839\ : CascadeMux
    port map (
            O => \N__45732\,
            I => \N__45729\
        );

    \I__9838\ : InMux
    port map (
            O => \N__45729\,
            I => \N__45726\
        );

    \I__9837\ : LocalMux
    port map (
            O => \N__45726\,
            I => \N__45723\
        );

    \I__9836\ : Span4Mux_v
    port map (
            O => \N__45723\,
            I => \N__45720\
        );

    \I__9835\ : Odrv4
    port map (
            O => \N__45720\,
            I => n17_adj_635
        );

    \I__9834\ : CascadeMux
    port map (
            O => \N__45717\,
            I => \n1129_cascade_\
        );

    \I__9833\ : CascadeMux
    port map (
            O => \N__45714\,
            I => \n1625_adj_605_cascade_\
        );

    \I__9832\ : InMux
    port map (
            O => \N__45711\,
            I => \N__45708\
        );

    \I__9831\ : LocalMux
    port map (
            O => \N__45708\,
            I => \N__45705\
        );

    \I__9830\ : Odrv4
    port map (
            O => \N__45705\,
            I => n1698
        );

    \I__9829\ : InMux
    port map (
            O => \N__45702\,
            I => \N__45698\
        );

    \I__9828\ : CascadeMux
    port map (
            O => \N__45701\,
            I => \N__45695\
        );

    \I__9827\ : LocalMux
    port map (
            O => \N__45698\,
            I => \N__45692\
        );

    \I__9826\ : InMux
    port map (
            O => \N__45695\,
            I => \N__45689\
        );

    \I__9825\ : Odrv4
    port map (
            O => \N__45692\,
            I => n1730
        );

    \I__9824\ : LocalMux
    port map (
            O => \N__45689\,
            I => n1730
        );

    \I__9823\ : CascadeMux
    port map (
            O => \N__45684\,
            I => \n1730_cascade_\
        );

    \I__9822\ : CascadeMux
    port map (
            O => \N__45681\,
            I => \N__45678\
        );

    \I__9821\ : InMux
    port map (
            O => \N__45678\,
            I => \N__45674\
        );

    \I__9820\ : CascadeMux
    port map (
            O => \N__45677\,
            I => \N__45671\
        );

    \I__9819\ : LocalMux
    port map (
            O => \N__45674\,
            I => \N__45667\
        );

    \I__9818\ : InMux
    port map (
            O => \N__45671\,
            I => \N__45664\
        );

    \I__9817\ : InMux
    port map (
            O => \N__45670\,
            I => \N__45661\
        );

    \I__9816\ : Odrv4
    port map (
            O => \N__45667\,
            I => n1729
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__45664\,
            I => n1729
        );

    \I__9814\ : LocalMux
    port map (
            O => \N__45661\,
            I => n1729
        );

    \I__9813\ : InMux
    port map (
            O => \N__45654\,
            I => \N__45651\
        );

    \I__9812\ : LocalMux
    port map (
            O => \N__45651\,
            I => \N__45648\
        );

    \I__9811\ : Odrv4
    port map (
            O => \N__45648\,
            I => n14514
        );

    \I__9810\ : CascadeMux
    port map (
            O => \N__45645\,
            I => \N__45642\
        );

    \I__9809\ : InMux
    port map (
            O => \N__45642\,
            I => \N__45639\
        );

    \I__9808\ : LocalMux
    port map (
            O => \N__45639\,
            I => \N__45636\
        );

    \I__9807\ : Span4Mux_v
    port map (
            O => \N__45636\,
            I => \N__45633\
        );

    \I__9806\ : Odrv4
    port map (
            O => \N__45633\,
            I => n11_adj_629
        );

    \I__9805\ : InMux
    port map (
            O => \N__45630\,
            I => \N__45627\
        );

    \I__9804\ : LocalMux
    port map (
            O => \N__45627\,
            I => \N__45624\
        );

    \I__9803\ : Odrv12
    port map (
            O => \N__45624\,
            I => n1701
        );

    \I__9802\ : InMux
    port map (
            O => \N__45621\,
            I => \N__45618\
        );

    \I__9801\ : LocalMux
    port map (
            O => \N__45618\,
            I => \N__45610\
        );

    \I__9800\ : CascadeMux
    port map (
            O => \N__45617\,
            I => \N__45605\
        );

    \I__9799\ : CascadeMux
    port map (
            O => \N__45616\,
            I => \N__45599\
        );

    \I__9798\ : CascadeMux
    port map (
            O => \N__45615\,
            I => \N__45594\
        );

    \I__9797\ : CascadeMux
    port map (
            O => \N__45614\,
            I => \N__45591\
        );

    \I__9796\ : CascadeMux
    port map (
            O => \N__45613\,
            I => \N__45588\
        );

    \I__9795\ : Span12Mux_h
    port map (
            O => \N__45610\,
            I => \N__45583\
        );

    \I__9794\ : InMux
    port map (
            O => \N__45609\,
            I => \N__45578\
        );

    \I__9793\ : InMux
    port map (
            O => \N__45608\,
            I => \N__45578\
        );

    \I__9792\ : InMux
    port map (
            O => \N__45605\,
            I => \N__45575\
        );

    \I__9791\ : InMux
    port map (
            O => \N__45604\,
            I => \N__45564\
        );

    \I__9790\ : InMux
    port map (
            O => \N__45603\,
            I => \N__45564\
        );

    \I__9789\ : InMux
    port map (
            O => \N__45602\,
            I => \N__45564\
        );

    \I__9788\ : InMux
    port map (
            O => \N__45599\,
            I => \N__45564\
        );

    \I__9787\ : InMux
    port map (
            O => \N__45598\,
            I => \N__45564\
        );

    \I__9786\ : InMux
    port map (
            O => \N__45597\,
            I => \N__45559\
        );

    \I__9785\ : InMux
    port map (
            O => \N__45594\,
            I => \N__45559\
        );

    \I__9784\ : InMux
    port map (
            O => \N__45591\,
            I => \N__45550\
        );

    \I__9783\ : InMux
    port map (
            O => \N__45588\,
            I => \N__45550\
        );

    \I__9782\ : InMux
    port map (
            O => \N__45587\,
            I => \N__45550\
        );

    \I__9781\ : InMux
    port map (
            O => \N__45586\,
            I => \N__45550\
        );

    \I__9780\ : Odrv12
    port map (
            O => \N__45583\,
            I => n1653
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__45578\,
            I => n1653
        );

    \I__9778\ : LocalMux
    port map (
            O => \N__45575\,
            I => n1653
        );

    \I__9777\ : LocalMux
    port map (
            O => \N__45564\,
            I => n1653
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__45559\,
            I => n1653
        );

    \I__9775\ : LocalMux
    port map (
            O => \N__45550\,
            I => n1653
        );

    \I__9774\ : InMux
    port map (
            O => \N__45537\,
            I => \N__45534\
        );

    \I__9773\ : LocalMux
    port map (
            O => \N__45534\,
            I => \N__45530\
        );

    \I__9772\ : CascadeMux
    port map (
            O => \N__45533\,
            I => \N__45527\
        );

    \I__9771\ : Span4Mux_h
    port map (
            O => \N__45530\,
            I => \N__45523\
        );

    \I__9770\ : InMux
    port map (
            O => \N__45527\,
            I => \N__45520\
        );

    \I__9769\ : InMux
    port map (
            O => \N__45526\,
            I => \N__45517\
        );

    \I__9768\ : Odrv4
    port map (
            O => \N__45523\,
            I => n1733
        );

    \I__9767\ : LocalMux
    port map (
            O => \N__45520\,
            I => n1733
        );

    \I__9766\ : LocalMux
    port map (
            O => \N__45517\,
            I => n1733
        );

    \I__9765\ : InMux
    port map (
            O => \N__45510\,
            I => \N__45507\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__45507\,
            I => \N__45503\
        );

    \I__9763\ : CascadeMux
    port map (
            O => \N__45506\,
            I => \N__45496\
        );

    \I__9762\ : Span4Mux_v
    port map (
            O => \N__45503\,
            I => \N__45493\
        );

    \I__9761\ : InMux
    port map (
            O => \N__45502\,
            I => \N__45490\
        );

    \I__9760\ : CascadeMux
    port map (
            O => \N__45501\,
            I => \N__45487\
        );

    \I__9759\ : InMux
    port map (
            O => \N__45500\,
            I => \N__45481\
        );

    \I__9758\ : CascadeMux
    port map (
            O => \N__45499\,
            I => \N__45477\
        );

    \I__9757\ : InMux
    port map (
            O => \N__45496\,
            I => \N__45473\
        );

    \I__9756\ : Span4Mux_h
    port map (
            O => \N__45493\,
            I => \N__45468\
        );

    \I__9755\ : LocalMux
    port map (
            O => \N__45490\,
            I => \N__45468\
        );

    \I__9754\ : InMux
    port map (
            O => \N__45487\,
            I => \N__45465\
        );

    \I__9753\ : CascadeMux
    port map (
            O => \N__45486\,
            I => \N__45462\
        );

    \I__9752\ : CascadeMux
    port map (
            O => \N__45485\,
            I => \N__45458\
        );

    \I__9751\ : InMux
    port map (
            O => \N__45484\,
            I => \N__45451\
        );

    \I__9750\ : LocalMux
    port map (
            O => \N__45481\,
            I => \N__45448\
        );

    \I__9749\ : InMux
    port map (
            O => \N__45480\,
            I => \N__45445\
        );

    \I__9748\ : InMux
    port map (
            O => \N__45477\,
            I => \N__45440\
        );

    \I__9747\ : InMux
    port map (
            O => \N__45476\,
            I => \N__45440\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__45473\,
            I => \N__45433\
        );

    \I__9745\ : Span4Mux_v
    port map (
            O => \N__45468\,
            I => \N__45433\
        );

    \I__9744\ : LocalMux
    port map (
            O => \N__45465\,
            I => \N__45433\
        );

    \I__9743\ : InMux
    port map (
            O => \N__45462\,
            I => \N__45422\
        );

    \I__9742\ : InMux
    port map (
            O => \N__45461\,
            I => \N__45422\
        );

    \I__9741\ : InMux
    port map (
            O => \N__45458\,
            I => \N__45422\
        );

    \I__9740\ : InMux
    port map (
            O => \N__45457\,
            I => \N__45422\
        );

    \I__9739\ : InMux
    port map (
            O => \N__45456\,
            I => \N__45422\
        );

    \I__9738\ : InMux
    port map (
            O => \N__45455\,
            I => \N__45417\
        );

    \I__9737\ : InMux
    port map (
            O => \N__45454\,
            I => \N__45417\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__45451\,
            I => \N__45410\
        );

    \I__9735\ : Span4Mux_h
    port map (
            O => \N__45448\,
            I => \N__45410\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__45445\,
            I => \N__45410\
        );

    \I__9733\ : LocalMux
    port map (
            O => \N__45440\,
            I => n1752
        );

    \I__9732\ : Odrv4
    port map (
            O => \N__45433\,
            I => n1752
        );

    \I__9731\ : LocalMux
    port map (
            O => \N__45422\,
            I => n1752
        );

    \I__9730\ : LocalMux
    port map (
            O => \N__45417\,
            I => n1752
        );

    \I__9729\ : Odrv4
    port map (
            O => \N__45410\,
            I => n1752
        );

    \I__9728\ : InMux
    port map (
            O => \N__45399\,
            I => \N__45396\
        );

    \I__9727\ : LocalMux
    port map (
            O => \N__45396\,
            I => \N__45393\
        );

    \I__9726\ : Span4Mux_h
    port map (
            O => \N__45393\,
            I => \N__45390\
        );

    \I__9725\ : Span4Mux_h
    port map (
            O => \N__45390\,
            I => \N__45386\
        );

    \I__9724\ : CascadeMux
    port map (
            O => \N__45389\,
            I => \N__45383\
        );

    \I__9723\ : Span4Mux_v
    port map (
            O => \N__45386\,
            I => \N__45380\
        );

    \I__9722\ : InMux
    port map (
            O => \N__45383\,
            I => \N__45377\
        );

    \I__9721\ : Odrv4
    port map (
            O => \N__45380\,
            I => n15630
        );

    \I__9720\ : LocalMux
    port map (
            O => \N__45377\,
            I => n15630
        );

    \I__9719\ : CascadeMux
    port map (
            O => \N__45372\,
            I => \N__45368\
        );

    \I__9718\ : InMux
    port map (
            O => \N__45371\,
            I => \N__45365\
        );

    \I__9717\ : InMux
    port map (
            O => \N__45368\,
            I => \N__45361\
        );

    \I__9716\ : LocalMux
    port map (
            O => \N__45365\,
            I => \N__45358\
        );

    \I__9715\ : InMux
    port map (
            O => \N__45364\,
            I => \N__45355\
        );

    \I__9714\ : LocalMux
    port map (
            O => \N__45361\,
            I => n1621_adj_601
        );

    \I__9713\ : Odrv4
    port map (
            O => \N__45358\,
            I => n1621_adj_601
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__45355\,
            I => n1621_adj_601
        );

    \I__9711\ : InMux
    port map (
            O => \N__45348\,
            I => n12590
        );

    \I__9710\ : InMux
    port map (
            O => \N__45345\,
            I => \N__45342\
        );

    \I__9709\ : LocalMux
    port map (
            O => \N__45342\,
            I => \N__45338\
        );

    \I__9708\ : CascadeMux
    port map (
            O => \N__45341\,
            I => \N__45335\
        );

    \I__9707\ : Span4Mux_v
    port map (
            O => \N__45338\,
            I => \N__45332\
        );

    \I__9706\ : InMux
    port map (
            O => \N__45335\,
            I => \N__45329\
        );

    \I__9705\ : Odrv4
    port map (
            O => \N__45332\,
            I => n1719
        );

    \I__9704\ : LocalMux
    port map (
            O => \N__45329\,
            I => n1719
        );

    \I__9703\ : InMux
    port map (
            O => \N__45324\,
            I => \N__45321\
        );

    \I__9702\ : LocalMux
    port map (
            O => \N__45321\,
            I => n1695
        );

    \I__9701\ : CascadeMux
    port map (
            O => \N__45318\,
            I => \N__45315\
        );

    \I__9700\ : InMux
    port map (
            O => \N__45315\,
            I => \N__45311\
        );

    \I__9699\ : InMux
    port map (
            O => \N__45314\,
            I => \N__45307\
        );

    \I__9698\ : LocalMux
    port map (
            O => \N__45311\,
            I => \N__45304\
        );

    \I__9697\ : InMux
    port map (
            O => \N__45310\,
            I => \N__45301\
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__45307\,
            I => n1727
        );

    \I__9695\ : Odrv4
    port map (
            O => \N__45304\,
            I => n1727
        );

    \I__9694\ : LocalMux
    port map (
            O => \N__45301\,
            I => n1727
        );

    \I__9693\ : InMux
    port map (
            O => \N__45294\,
            I => \N__45291\
        );

    \I__9692\ : LocalMux
    port map (
            O => \N__45291\,
            I => \N__45288\
        );

    \I__9691\ : Odrv4
    port map (
            O => \N__45288\,
            I => n1696
        );

    \I__9690\ : CascadeMux
    port map (
            O => \N__45285\,
            I => \n1653_cascade_\
        );

    \I__9689\ : CascadeMux
    port map (
            O => \N__45282\,
            I => \N__45279\
        );

    \I__9688\ : InMux
    port map (
            O => \N__45279\,
            I => \N__45274\
        );

    \I__9687\ : InMux
    port map (
            O => \N__45278\,
            I => \N__45269\
        );

    \I__9686\ : InMux
    port map (
            O => \N__45277\,
            I => \N__45269\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__45274\,
            I => n1728
        );

    \I__9684\ : LocalMux
    port map (
            O => \N__45269\,
            I => n1728
        );

    \I__9683\ : CascadeMux
    port map (
            O => \N__45264\,
            I => \N__45261\
        );

    \I__9682\ : InMux
    port map (
            O => \N__45261\,
            I => \N__45258\
        );

    \I__9681\ : LocalMux
    port map (
            O => \N__45258\,
            I => \N__45255\
        );

    \I__9680\ : Odrv4
    port map (
            O => \N__45255\,
            I => n1697
        );

    \I__9679\ : InMux
    port map (
            O => \N__45252\,
            I => \N__45249\
        );

    \I__9678\ : LocalMux
    port map (
            O => \N__45249\,
            I => n1692
        );

    \I__9677\ : CascadeMux
    port map (
            O => \N__45246\,
            I => \N__45242\
        );

    \I__9676\ : InMux
    port map (
            O => \N__45245\,
            I => \N__45239\
        );

    \I__9675\ : InMux
    port map (
            O => \N__45242\,
            I => \N__45236\
        );

    \I__9674\ : LocalMux
    port map (
            O => \N__45239\,
            I => \N__45232\
        );

    \I__9673\ : LocalMux
    port map (
            O => \N__45236\,
            I => \N__45229\
        );

    \I__9672\ : InMux
    port map (
            O => \N__45235\,
            I => \N__45226\
        );

    \I__9671\ : Odrv4
    port map (
            O => \N__45232\,
            I => n1724
        );

    \I__9670\ : Odrv4
    port map (
            O => \N__45229\,
            I => n1724
        );

    \I__9669\ : LocalMux
    port map (
            O => \N__45226\,
            I => n1724
        );

    \I__9668\ : CascadeMux
    port map (
            O => \N__45219\,
            I => \N__45216\
        );

    \I__9667\ : InMux
    port map (
            O => \N__45216\,
            I => \N__45213\
        );

    \I__9666\ : LocalMux
    port map (
            O => \N__45213\,
            I => n1693_adj_614
        );

    \I__9665\ : CascadeMux
    port map (
            O => \N__45210\,
            I => \N__45206\
        );

    \I__9664\ : CascadeMux
    port map (
            O => \N__45209\,
            I => \N__45203\
        );

    \I__9663\ : InMux
    port map (
            O => \N__45206\,
            I => \N__45200\
        );

    \I__9662\ : InMux
    port map (
            O => \N__45203\,
            I => \N__45197\
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__45200\,
            I => \N__45193\
        );

    \I__9660\ : LocalMux
    port map (
            O => \N__45197\,
            I => \N__45190\
        );

    \I__9659\ : InMux
    port map (
            O => \N__45196\,
            I => \N__45187\
        );

    \I__9658\ : Odrv4
    port map (
            O => \N__45193\,
            I => n1725
        );

    \I__9657\ : Odrv4
    port map (
            O => \N__45190\,
            I => n1725
        );

    \I__9656\ : LocalMux
    port map (
            O => \N__45187\,
            I => n1725
        );

    \I__9655\ : InMux
    port map (
            O => \N__45180\,
            I => \N__45177\
        );

    \I__9654\ : LocalMux
    port map (
            O => \N__45177\,
            I => \N__45174\
        );

    \I__9653\ : Span4Mux_h
    port map (
            O => \N__45174\,
            I => \N__45171\
        );

    \I__9652\ : Span4Mux_v
    port map (
            O => \N__45171\,
            I => \N__45168\
        );

    \I__9651\ : Span4Mux_v
    port map (
            O => \N__45168\,
            I => \N__45164\
        );

    \I__9650\ : InMux
    port map (
            O => \N__45167\,
            I => \N__45161\
        );

    \I__9649\ : Odrv4
    port map (
            O => \N__45164\,
            I => n15611
        );

    \I__9648\ : LocalMux
    port map (
            O => \N__45161\,
            I => n15611
        );

    \I__9647\ : CascadeMux
    port map (
            O => \N__45156\,
            I => \N__45152\
        );

    \I__9646\ : InMux
    port map (
            O => \N__45155\,
            I => \N__45149\
        );

    \I__9645\ : InMux
    port map (
            O => \N__45152\,
            I => \N__45146\
        );

    \I__9644\ : LocalMux
    port map (
            O => \N__45149\,
            I => n1625_adj_605
        );

    \I__9643\ : LocalMux
    port map (
            O => \N__45146\,
            I => n1625_adj_605
        );

    \I__9642\ : InMux
    port map (
            O => \N__45141\,
            I => n12581
        );

    \I__9641\ : InMux
    port map (
            O => \N__45138\,
            I => n12582
        );

    \I__9640\ : InMux
    port map (
            O => \N__45135\,
            I => \N__45132\
        );

    \I__9639\ : LocalMux
    port map (
            O => \N__45132\,
            I => n1694
        );

    \I__9638\ : InMux
    port map (
            O => \N__45129\,
            I => n12583
        );

    \I__9637\ : InMux
    port map (
            O => \N__45126\,
            I => \bfn_13_18_0_\
        );

    \I__9636\ : InMux
    port map (
            O => \N__45123\,
            I => n12585
        );

    \I__9635\ : InMux
    port map (
            O => \N__45120\,
            I => \N__45117\
        );

    \I__9634\ : LocalMux
    port map (
            O => \N__45117\,
            I => n1691
        );

    \I__9633\ : InMux
    port map (
            O => \N__45114\,
            I => n12586
        );

    \I__9632\ : CascadeMux
    port map (
            O => \N__45111\,
            I => \N__45108\
        );

    \I__9631\ : InMux
    port map (
            O => \N__45108\,
            I => \N__45105\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__45105\,
            I => n1690
        );

    \I__9629\ : InMux
    port map (
            O => \N__45102\,
            I => n12587
        );

    \I__9628\ : CascadeMux
    port map (
            O => \N__45099\,
            I => \N__45096\
        );

    \I__9627\ : InMux
    port map (
            O => \N__45096\,
            I => \N__45093\
        );

    \I__9626\ : LocalMux
    port map (
            O => \N__45093\,
            I => n1689
        );

    \I__9625\ : InMux
    port map (
            O => \N__45090\,
            I => n12588
        );

    \I__9624\ : InMux
    port map (
            O => \N__45087\,
            I => \N__45084\
        );

    \I__9623\ : LocalMux
    port map (
            O => \N__45084\,
            I => n1688
        );

    \I__9622\ : InMux
    port map (
            O => \N__45081\,
            I => n12589
        );

    \I__9621\ : InMux
    port map (
            O => \N__45078\,
            I => \N__45072\
        );

    \I__9620\ : InMux
    port map (
            O => \N__45077\,
            I => \N__45072\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__45072\,
            I => n33_adj_675
        );

    \I__9618\ : CascadeMux
    port map (
            O => \N__45069\,
            I => \N__45066\
        );

    \I__9617\ : InMux
    port map (
            O => \N__45066\,
            I => \N__45063\
        );

    \I__9616\ : LocalMux
    port map (
            O => \N__45063\,
            I => n15104
        );

    \I__9615\ : InMux
    port map (
            O => \N__45060\,
            I => \N__45054\
        );

    \I__9614\ : InMux
    port map (
            O => \N__45059\,
            I => \N__45054\
        );

    \I__9613\ : LocalMux
    port map (
            O => \N__45054\,
            I => n31_adj_674
        );

    \I__9612\ : CascadeMux
    port map (
            O => \N__45051\,
            I => \N__45046\
        );

    \I__9611\ : InMux
    port map (
            O => \N__45050\,
            I => \N__45039\
        );

    \I__9610\ : InMux
    port map (
            O => \N__45049\,
            I => \N__45039\
        );

    \I__9609\ : InMux
    port map (
            O => \N__45046\,
            I => \N__45039\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__45039\,
            I => n35
        );

    \I__9607\ : InMux
    port map (
            O => \N__45036\,
            I => \N__45033\
        );

    \I__9606\ : LocalMux
    port map (
            O => \N__45033\,
            I => n15247
        );

    \I__9605\ : CascadeMux
    port map (
            O => \N__45030\,
            I => \n15099_cascade_\
        );

    \I__9604\ : InMux
    port map (
            O => \N__45027\,
            I => \N__45024\
        );

    \I__9603\ : LocalMux
    port map (
            O => \N__45024\,
            I => n15220
        );

    \I__9602\ : InMux
    port map (
            O => \N__45021\,
            I => \N__45015\
        );

    \I__9601\ : InMux
    port map (
            O => \N__45020\,
            I => \N__45015\
        );

    \I__9600\ : LocalMux
    port map (
            O => \N__45015\,
            I => \N__45012\
        );

    \I__9599\ : Odrv4
    port map (
            O => \N__45012\,
            I => pwm_setpoint_18
        );

    \I__9598\ : CascadeMux
    port map (
            O => \N__45009\,
            I => \n15257_cascade_\
        );

    \I__9597\ : InMux
    port map (
            O => \N__45006\,
            I => \N__45000\
        );

    \I__9596\ : InMux
    port map (
            O => \N__45005\,
            I => \N__45000\
        );

    \I__9595\ : LocalMux
    port map (
            O => \N__45000\,
            I => n37
        );

    \I__9594\ : InMux
    port map (
            O => \N__44997\,
            I => \N__44994\
        );

    \I__9593\ : LocalMux
    port map (
            O => \N__44994\,
            I => \N__44991\
        );

    \I__9592\ : Odrv4
    port map (
            O => \N__44991\,
            I => n15258
        );

    \I__9591\ : InMux
    port map (
            O => \N__44988\,
            I => \bfn_13_17_0_\
        );

    \I__9590\ : InMux
    port map (
            O => \N__44985\,
            I => \N__44982\
        );

    \I__9589\ : LocalMux
    port map (
            O => \N__44982\,
            I => \N__44979\
        );

    \I__9588\ : Odrv4
    port map (
            O => \N__44979\,
            I => n1700
        );

    \I__9587\ : InMux
    port map (
            O => \N__44976\,
            I => n12577
        );

    \I__9586\ : InMux
    port map (
            O => \N__44973\,
            I => \N__44970\
        );

    \I__9585\ : LocalMux
    port map (
            O => \N__44970\,
            I => \N__44967\
        );

    \I__9584\ : Odrv4
    port map (
            O => \N__44967\,
            I => n1699
        );

    \I__9583\ : InMux
    port map (
            O => \N__44964\,
            I => n12578
        );

    \I__9582\ : InMux
    port map (
            O => \N__44961\,
            I => n12579
        );

    \I__9581\ : InMux
    port map (
            O => \N__44958\,
            I => n12580
        );

    \I__9580\ : InMux
    port map (
            O => \N__44955\,
            I => \N__44951\
        );

    \I__9579\ : InMux
    port map (
            O => \N__44954\,
            I => \N__44948\
        );

    \I__9578\ : LocalMux
    port map (
            O => \N__44951\,
            I => \N__44943\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__44948\,
            I => \N__44943\
        );

    \I__9576\ : Span4Mux_s3_v
    port map (
            O => \N__44943\,
            I => \N__44940\
        );

    \I__9575\ : Odrv4
    port map (
            O => \N__44940\,
            I => duty_12
        );

    \I__9574\ : InMux
    port map (
            O => \N__44937\,
            I => \N__44934\
        );

    \I__9573\ : LocalMux
    port map (
            O => \N__44934\,
            I => \N__44931\
        );

    \I__9572\ : Span4Mux_h
    port map (
            O => \N__44931\,
            I => \N__44928\
        );

    \I__9571\ : Odrv4
    port map (
            O => \N__44928\,
            I => n13_adj_585
        );

    \I__9570\ : CascadeMux
    port map (
            O => \N__44925\,
            I => \n31_adj_674_cascade_\
        );

    \I__9569\ : InMux
    port map (
            O => \N__44922\,
            I => \N__44919\
        );

    \I__9568\ : LocalMux
    port map (
            O => \N__44919\,
            I => n15230
        );

    \I__9567\ : InMux
    port map (
            O => \N__44916\,
            I => \N__44913\
        );

    \I__9566\ : LocalMux
    port map (
            O => \N__44913\,
            I => n15237
        );

    \I__9565\ : CascadeMux
    port map (
            O => \N__44910\,
            I => \n15195_cascade_\
        );

    \I__9564\ : InMux
    port map (
            O => \N__44907\,
            I => \N__44904\
        );

    \I__9563\ : LocalMux
    port map (
            O => \N__44904\,
            I => \N__44901\
        );

    \I__9562\ : Odrv4
    port map (
            O => \N__44901\,
            I => n15241
        );

    \I__9561\ : InMux
    port map (
            O => \N__44898\,
            I => \N__44895\
        );

    \I__9560\ : LocalMux
    port map (
            O => \N__44895\,
            I => n15097
        );

    \I__9559\ : InMux
    port map (
            O => \N__44892\,
            I => \N__44889\
        );

    \I__9558\ : LocalMux
    port map (
            O => \N__44889\,
            I => n10_adj_659
        );

    \I__9557\ : InMux
    port map (
            O => \N__44886\,
            I => \N__44883\
        );

    \I__9556\ : LocalMux
    port map (
            O => \N__44883\,
            I => n30_adj_673
        );

    \I__9555\ : InMux
    port map (
            O => \N__44880\,
            I => \N__44875\
        );

    \I__9554\ : InMux
    port map (
            O => \N__44879\,
            I => \N__44870\
        );

    \I__9553\ : InMux
    port map (
            O => \N__44878\,
            I => \N__44870\
        );

    \I__9552\ : LocalMux
    port map (
            O => \N__44875\,
            I => pwm_setpoint_21
        );

    \I__9551\ : LocalMux
    port map (
            O => \N__44870\,
            I => pwm_setpoint_21
        );

    \I__9550\ : InMux
    port map (
            O => \N__44865\,
            I => \N__44862\
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__44862\,
            I => \N__44859\
        );

    \I__9548\ : Odrv4
    port map (
            O => \N__44859\,
            I => \pwm_setpoint_23_N_171_12\
        );

    \I__9547\ : InMux
    port map (
            O => \N__44856\,
            I => \N__44853\
        );

    \I__9546\ : LocalMux
    port map (
            O => \N__44853\,
            I => n39_adj_676
        );

    \I__9545\ : CascadeMux
    port map (
            O => \N__44850\,
            I => \N__44847\
        );

    \I__9544\ : InMux
    port map (
            O => \N__44847\,
            I => \N__44844\
        );

    \I__9543\ : LocalMux
    port map (
            O => \N__44844\,
            I => \N__44841\
        );

    \I__9542\ : Odrv4
    port map (
            O => \N__44841\,
            I => n41_adj_678
        );

    \I__9541\ : InMux
    port map (
            O => \N__44838\,
            I => \N__44835\
        );

    \I__9540\ : LocalMux
    port map (
            O => \N__44835\,
            I => \N__44832\
        );

    \I__9539\ : Odrv12
    port map (
            O => \N__44832\,
            I => n15091
        );

    \I__9538\ : InMux
    port map (
            O => \N__44829\,
            I => \N__44826\
        );

    \I__9537\ : LocalMux
    port map (
            O => \N__44826\,
            I => \N__44823\
        );

    \I__9536\ : Odrv4
    port map (
            O => \N__44823\,
            I => n4_adj_655
        );

    \I__9535\ : InMux
    port map (
            O => \N__44820\,
            I => \N__44816\
        );

    \I__9534\ : InMux
    port map (
            O => \N__44819\,
            I => \N__44813\
        );

    \I__9533\ : LocalMux
    port map (
            O => \N__44816\,
            I => pwm_setpoint_12
        );

    \I__9532\ : LocalMux
    port map (
            O => \N__44813\,
            I => pwm_setpoint_12
        );

    \I__9531\ : InMux
    port map (
            O => \N__44808\,
            I => \N__44802\
        );

    \I__9530\ : InMux
    port map (
            O => \N__44807\,
            I => \N__44802\
        );

    \I__9529\ : LocalMux
    port map (
            O => \N__44802\,
            I => n25_adj_670
        );

    \I__9528\ : InMux
    port map (
            O => \N__44799\,
            I => \N__44796\
        );

    \I__9527\ : LocalMux
    port map (
            O => \N__44796\,
            I => \N__44793\
        );

    \I__9526\ : Odrv4
    port map (
            O => \N__44793\,
            I => n15110
        );

    \I__9525\ : InMux
    port map (
            O => \N__44790\,
            I => \N__44785\
        );

    \I__9524\ : InMux
    port map (
            O => \N__44789\,
            I => \N__44782\
        );

    \I__9523\ : InMux
    port map (
            O => \N__44788\,
            I => \N__44779\
        );

    \I__9522\ : LocalMux
    port map (
            O => \N__44785\,
            I => \N__44774\
        );

    \I__9521\ : LocalMux
    port map (
            O => \N__44782\,
            I => \N__44774\
        );

    \I__9520\ : LocalMux
    port map (
            O => \N__44779\,
            I => n23_adj_668
        );

    \I__9519\ : Odrv4
    port map (
            O => \N__44774\,
            I => n23_adj_668
        );

    \I__9518\ : CascadeMux
    port map (
            O => \N__44769\,
            I => \n25_adj_670_cascade_\
        );

    \I__9517\ : InMux
    port map (
            O => \N__44766\,
            I => \N__44760\
        );

    \I__9516\ : InMux
    port map (
            O => \N__44765\,
            I => \N__44760\
        );

    \I__9515\ : LocalMux
    port map (
            O => \N__44760\,
            I => n43
        );

    \I__9514\ : CascadeMux
    port map (
            O => \N__44757\,
            I => \N__44754\
        );

    \I__9513\ : InMux
    port map (
            O => \N__44754\,
            I => \N__44751\
        );

    \I__9512\ : LocalMux
    port map (
            O => \N__44751\,
            I => n15146
        );

    \I__9511\ : InMux
    port map (
            O => \N__44748\,
            I => \N__44744\
        );

    \I__9510\ : InMux
    port map (
            O => \N__44747\,
            I => \N__44741\
        );

    \I__9509\ : LocalMux
    port map (
            O => \N__44744\,
            I => \N__44738\
        );

    \I__9508\ : LocalMux
    port map (
            O => \N__44741\,
            I => n13_adj_662
        );

    \I__9507\ : Odrv4
    port map (
            O => \N__44738\,
            I => n13_adj_662
        );

    \I__9506\ : InMux
    port map (
            O => \N__44733\,
            I => \N__44729\
        );

    \I__9505\ : InMux
    port map (
            O => \N__44732\,
            I => \N__44726\
        );

    \I__9504\ : LocalMux
    port map (
            O => \N__44729\,
            I => n15_adj_663
        );

    \I__9503\ : LocalMux
    port map (
            O => \N__44726\,
            I => n15_adj_663
        );

    \I__9502\ : InMux
    port map (
            O => \N__44721\,
            I => \N__44718\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__44718\,
            I => n15229
        );

    \I__9500\ : InMux
    port map (
            O => \N__44715\,
            I => \N__44712\
        );

    \I__9499\ : LocalMux
    port map (
            O => \N__44712\,
            I => \N__44708\
        );

    \I__9498\ : InMux
    port map (
            O => \N__44711\,
            I => \N__44705\
        );

    \I__9497\ : Odrv4
    port map (
            O => \N__44708\,
            I => pwm_setpoint_22
        );

    \I__9496\ : LocalMux
    port map (
            O => \N__44705\,
            I => pwm_setpoint_22
        );

    \I__9495\ : CascadeMux
    port map (
            O => \N__44700\,
            I => \n45_cascade_\
        );

    \I__9494\ : InMux
    port map (
            O => \N__44697\,
            I => \N__44691\
        );

    \I__9493\ : InMux
    port map (
            O => \N__44696\,
            I => \N__44691\
        );

    \I__9492\ : LocalMux
    port map (
            O => \N__44691\,
            I => pwm_setpoint_20
        );

    \I__9491\ : CascadeMux
    port map (
            O => \N__44688\,
            I => \n41_adj_678_cascade_\
        );

    \I__9490\ : InMux
    port map (
            O => \N__44685\,
            I => \N__44682\
        );

    \I__9489\ : LocalMux
    port map (
            O => \N__44682\,
            I => n40_adj_677
        );

    \I__9488\ : InMux
    port map (
            O => \N__44679\,
            I => \N__44674\
        );

    \I__9487\ : InMux
    port map (
            O => \N__44678\,
            I => \N__44669\
        );

    \I__9486\ : InMux
    port map (
            O => \N__44677\,
            I => \N__44669\
        );

    \I__9485\ : LocalMux
    port map (
            O => \N__44674\,
            I => n45
        );

    \I__9484\ : LocalMux
    port map (
            O => \N__44669\,
            I => n45
        );

    \I__9483\ : InMux
    port map (
            O => \N__44664\,
            I => \N__44661\
        );

    \I__9482\ : LocalMux
    port map (
            O => \N__44661\,
            I => n15223
        );

    \I__9481\ : InMux
    port map (
            O => \N__44658\,
            I => \N__44655\
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__44655\,
            I => \N__44652\
        );

    \I__9479\ : Odrv4
    port map (
            O => \N__44652\,
            I => n15165
        );

    \I__9478\ : InMux
    port map (
            O => \N__44649\,
            I => \N__44646\
        );

    \I__9477\ : LocalMux
    port map (
            O => \N__44646\,
            I => n15243
        );

    \I__9476\ : InMux
    port map (
            O => \N__44643\,
            I => \N__44640\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__44640\,
            I => \N__44636\
        );

    \I__9474\ : InMux
    port map (
            O => \N__44639\,
            I => \N__44633\
        );

    \I__9473\ : Span4Mux_h
    port map (
            O => \N__44636\,
            I => \N__44628\
        );

    \I__9472\ : LocalMux
    port map (
            O => \N__44633\,
            I => \N__44628\
        );

    \I__9471\ : Odrv4
    port map (
            O => \N__44628\,
            I => duty_22
        );

    \I__9470\ : InMux
    port map (
            O => \N__44625\,
            I => \N__44622\
        );

    \I__9469\ : LocalMux
    port map (
            O => \N__44622\,
            I => n3_adj_575
        );

    \I__9468\ : InMux
    port map (
            O => \N__44619\,
            I => \N__44613\
        );

    \I__9467\ : InMux
    port map (
            O => \N__44618\,
            I => \N__44613\
        );

    \I__9466\ : LocalMux
    port map (
            O => \N__44613\,
            I => \N__44610\
        );

    \I__9465\ : Odrv4
    port map (
            O => \N__44610\,
            I => pwm_setpoint_19
        );

    \I__9464\ : CascadeMux
    port map (
            O => \N__44607\,
            I => \n39_adj_676_cascade_\
        );

    \I__9463\ : InMux
    port map (
            O => \N__44604\,
            I => \N__44601\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__44601\,
            I => n15254
        );

    \I__9461\ : InMux
    port map (
            O => \N__44598\,
            I => \N__44595\
        );

    \I__9460\ : LocalMux
    port map (
            O => \N__44595\,
            I => \N__44592\
        );

    \I__9459\ : Span4Mux_s3_v
    port map (
            O => \N__44592\,
            I => \N__44588\
        );

    \I__9458\ : InMux
    port map (
            O => \N__44591\,
            I => \N__44585\
        );

    \I__9457\ : Odrv4
    port map (
            O => \N__44588\,
            I => duty_17
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__44585\,
            I => duty_17
        );

    \I__9455\ : InMux
    port map (
            O => \N__44580\,
            I => \N__44577\
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__44577\,
            I => n8_adj_580
        );

    \I__9453\ : InMux
    port map (
            O => \N__44574\,
            I => \N__44571\
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__44571\,
            I => \N__44567\
        );

    \I__9451\ : InMux
    port map (
            O => \N__44570\,
            I => \N__44564\
        );

    \I__9450\ : Odrv4
    port map (
            O => \N__44567\,
            I => duty_21
        );

    \I__9449\ : LocalMux
    port map (
            O => \N__44564\,
            I => duty_21
        );

    \I__9448\ : InMux
    port map (
            O => \N__44559\,
            I => \N__44556\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__44556\,
            I => n4_adj_576
        );

    \I__9446\ : InMux
    port map (
            O => \N__44553\,
            I => \N__44550\
        );

    \I__9445\ : LocalMux
    port map (
            O => \N__44550\,
            I => \N__44547\
        );

    \I__9444\ : Span4Mux_s2_v
    port map (
            O => \N__44547\,
            I => \N__44544\
        );

    \I__9443\ : Span4Mux_h
    port map (
            O => \N__44544\,
            I => \N__44540\
        );

    \I__9442\ : InMux
    port map (
            O => \N__44543\,
            I => \N__44537\
        );

    \I__9441\ : Odrv4
    port map (
            O => \N__44540\,
            I => duty_18
        );

    \I__9440\ : LocalMux
    port map (
            O => \N__44537\,
            I => duty_18
        );

    \I__9439\ : InMux
    port map (
            O => \N__44532\,
            I => \N__44529\
        );

    \I__9438\ : LocalMux
    port map (
            O => \N__44529\,
            I => n7_adj_579
        );

    \I__9437\ : InMux
    port map (
            O => \N__44526\,
            I => \N__44523\
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__44523\,
            I => \pwm_setpoint_23_N_171_19\
        );

    \I__9435\ : InMux
    port map (
            O => \N__44520\,
            I => \N__44517\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__44517\,
            I => \pwm_setpoint_23_N_171_20\
        );

    \I__9433\ : InMux
    port map (
            O => \N__44514\,
            I => \N__44511\
        );

    \I__9432\ : LocalMux
    port map (
            O => \N__44511\,
            I => \N__44508\
        );

    \I__9431\ : Odrv4
    port map (
            O => \N__44508\,
            I => \pwm_setpoint_23_N_171_0\
        );

    \I__9430\ : InMux
    port map (
            O => \N__44505\,
            I => \N__44502\
        );

    \I__9429\ : LocalMux
    port map (
            O => \N__44502\,
            I => \N__44498\
        );

    \I__9428\ : InMux
    port map (
            O => \N__44501\,
            I => \N__44495\
        );

    \I__9427\ : Odrv12
    port map (
            O => \N__44498\,
            I => duty_0
        );

    \I__9426\ : LocalMux
    port map (
            O => \N__44495\,
            I => duty_0
        );

    \I__9425\ : InMux
    port map (
            O => \N__44490\,
            I => \N__44487\
        );

    \I__9424\ : LocalMux
    port map (
            O => \N__44487\,
            I => pwm_setpoint_0
        );

    \I__9423\ : InMux
    port map (
            O => \N__44484\,
            I => \N__44478\
        );

    \I__9422\ : InMux
    port map (
            O => \N__44483\,
            I => \N__44478\
        );

    \I__9421\ : LocalMux
    port map (
            O => \N__44478\,
            I => duty_20
        );

    \I__9420\ : InMux
    port map (
            O => \N__44475\,
            I => \N__44472\
        );

    \I__9419\ : LocalMux
    port map (
            O => \N__44472\,
            I => n5_adj_577
        );

    \I__9418\ : InMux
    port map (
            O => \N__44469\,
            I => \N__44466\
        );

    \I__9417\ : LocalMux
    port map (
            O => \N__44466\,
            I => \N__44463\
        );

    \I__9416\ : Span4Mux_h
    port map (
            O => \N__44463\,
            I => \N__44460\
        );

    \I__9415\ : Odrv4
    port map (
            O => \N__44460\,
            I => n10_adj_566
        );

    \I__9414\ : InMux
    port map (
            O => \N__44457\,
            I => n12487
        );

    \I__9413\ : InMux
    port map (
            O => \N__44454\,
            I => \N__44451\
        );

    \I__9412\ : LocalMux
    port map (
            O => \N__44451\,
            I => \N__44447\
        );

    \I__9411\ : InMux
    port map (
            O => \N__44450\,
            I => \N__44444\
        );

    \I__9410\ : Span4Mux_v
    port map (
            O => \N__44447\,
            I => \N__44439\
        );

    \I__9409\ : LocalMux
    port map (
            O => \N__44444\,
            I => \N__44439\
        );

    \I__9408\ : Span4Mux_h
    port map (
            O => \N__44439\,
            I => \N__44436\
        );

    \I__9407\ : Odrv4
    port map (
            O => \N__44436\,
            I => duty_16
        );

    \I__9406\ : InMux
    port map (
            O => \N__44433\,
            I => \bfn_12_27_0_\
        );

    \I__9405\ : InMux
    port map (
            O => \N__44430\,
            I => \N__44427\
        );

    \I__9404\ : LocalMux
    port map (
            O => \N__44427\,
            I => \N__44424\
        );

    \I__9403\ : Span4Mux_v
    port map (
            O => \N__44424\,
            I => \N__44421\
        );

    \I__9402\ : Odrv4
    port map (
            O => \N__44421\,
            I => n8_adj_568
        );

    \I__9401\ : InMux
    port map (
            O => \N__44418\,
            I => n12489
        );

    \I__9400\ : InMux
    port map (
            O => \N__44415\,
            I => \N__44412\
        );

    \I__9399\ : LocalMux
    port map (
            O => \N__44412\,
            I => \N__44409\
        );

    \I__9398\ : Odrv4
    port map (
            O => \N__44409\,
            I => n7_adj_569
        );

    \I__9397\ : InMux
    port map (
            O => \N__44406\,
            I => n12490
        );

    \I__9396\ : InMux
    port map (
            O => \N__44403\,
            I => \N__44400\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__44400\,
            I => \N__44397\
        );

    \I__9394\ : Odrv4
    port map (
            O => \N__44397\,
            I => n6_adj_570
        );

    \I__9393\ : InMux
    port map (
            O => \N__44394\,
            I => n12491
        );

    \I__9392\ : InMux
    port map (
            O => \N__44391\,
            I => \N__44388\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__44388\,
            I => \N__44385\
        );

    \I__9390\ : Span4Mux_v
    port map (
            O => \N__44385\,
            I => \N__44382\
        );

    \I__9389\ : Odrv4
    port map (
            O => \N__44382\,
            I => n5_adj_571
        );

    \I__9388\ : InMux
    port map (
            O => \N__44379\,
            I => n12492
        );

    \I__9387\ : InMux
    port map (
            O => \N__44376\,
            I => \N__44373\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__44373\,
            I => \N__44370\
        );

    \I__9385\ : Odrv4
    port map (
            O => \N__44370\,
            I => n4_adj_572
        );

    \I__9384\ : InMux
    port map (
            O => \N__44367\,
            I => n12493
        );

    \I__9383\ : InMux
    port map (
            O => \N__44364\,
            I => \N__44361\
        );

    \I__9382\ : LocalMux
    port map (
            O => \N__44361\,
            I => \N__44358\
        );

    \I__9381\ : Odrv4
    port map (
            O => \N__44358\,
            I => n3_adj_573
        );

    \I__9380\ : InMux
    port map (
            O => \N__44355\,
            I => n12494
        );

    \I__9379\ : InMux
    port map (
            O => \N__44352\,
            I => \N__44349\
        );

    \I__9378\ : LocalMux
    port map (
            O => \N__44349\,
            I => \N__44346\
        );

    \I__9377\ : Odrv4
    port map (
            O => \N__44346\,
            I => n2_adj_574
        );

    \I__9376\ : InMux
    port map (
            O => \N__44343\,
            I => n12495
        );

    \I__9375\ : InMux
    port map (
            O => \N__44340\,
            I => \N__44337\
        );

    \I__9374\ : LocalMux
    port map (
            O => \N__44337\,
            I => \N__44334\
        );

    \I__9373\ : Span4Mux_h
    port map (
            O => \N__44334\,
            I => \N__44330\
        );

    \I__9372\ : InMux
    port map (
            O => \N__44333\,
            I => \N__44327\
        );

    \I__9371\ : Odrv4
    port map (
            O => \N__44330\,
            I => duty_7
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__44327\,
            I => duty_7
        );

    \I__9369\ : InMux
    port map (
            O => \N__44322\,
            I => n12479
        );

    \I__9368\ : InMux
    port map (
            O => \N__44319\,
            I => \N__44316\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__44316\,
            I => \N__44313\
        );

    \I__9366\ : Odrv4
    port map (
            O => \N__44313\,
            I => n17_adj_559
        );

    \I__9365\ : InMux
    port map (
            O => \N__44310\,
            I => \N__44306\
        );

    \I__9364\ : InMux
    port map (
            O => \N__44309\,
            I => \N__44303\
        );

    \I__9363\ : LocalMux
    port map (
            O => \N__44306\,
            I => \N__44300\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__44303\,
            I => \N__44297\
        );

    \I__9361\ : Span4Mux_h
    port map (
            O => \N__44300\,
            I => \N__44294\
        );

    \I__9360\ : Span4Mux_h
    port map (
            O => \N__44297\,
            I => \N__44291\
        );

    \I__9359\ : Span4Mux_h
    port map (
            O => \N__44294\,
            I => \N__44288\
        );

    \I__9358\ : Odrv4
    port map (
            O => \N__44291\,
            I => duty_8
        );

    \I__9357\ : Odrv4
    port map (
            O => \N__44288\,
            I => duty_8
        );

    \I__9356\ : InMux
    port map (
            O => \N__44283\,
            I => \bfn_12_26_0_\
        );

    \I__9355\ : InMux
    port map (
            O => \N__44280\,
            I => \N__44277\
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__44277\,
            I => \N__44274\
        );

    \I__9353\ : Odrv4
    port map (
            O => \N__44274\,
            I => n16_adj_560
        );

    \I__9352\ : InMux
    port map (
            O => \N__44271\,
            I => \N__44267\
        );

    \I__9351\ : InMux
    port map (
            O => \N__44270\,
            I => \N__44264\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__44267\,
            I => \N__44261\
        );

    \I__9349\ : LocalMux
    port map (
            O => \N__44264\,
            I => \N__44258\
        );

    \I__9348\ : Span4Mux_v
    port map (
            O => \N__44261\,
            I => \N__44255\
        );

    \I__9347\ : Span12Mux_s6_v
    port map (
            O => \N__44258\,
            I => \N__44252\
        );

    \I__9346\ : Odrv4
    port map (
            O => \N__44255\,
            I => duty_9
        );

    \I__9345\ : Odrv12
    port map (
            O => \N__44252\,
            I => duty_9
        );

    \I__9344\ : InMux
    port map (
            O => \N__44247\,
            I => n12481
        );

    \I__9343\ : InMux
    port map (
            O => \N__44244\,
            I => \N__44241\
        );

    \I__9342\ : LocalMux
    port map (
            O => \N__44241\,
            I => \N__44238\
        );

    \I__9341\ : Odrv4
    port map (
            O => \N__44238\,
            I => n15_adj_561
        );

    \I__9340\ : InMux
    port map (
            O => \N__44235\,
            I => \N__44232\
        );

    \I__9339\ : LocalMux
    port map (
            O => \N__44232\,
            I => \N__44228\
        );

    \I__9338\ : InMux
    port map (
            O => \N__44231\,
            I => \N__44225\
        );

    \I__9337\ : Span4Mux_s3_v
    port map (
            O => \N__44228\,
            I => \N__44222\
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__44225\,
            I => \N__44219\
        );

    \I__9335\ : Odrv4
    port map (
            O => \N__44222\,
            I => duty_10
        );

    \I__9334\ : Odrv4
    port map (
            O => \N__44219\,
            I => duty_10
        );

    \I__9333\ : InMux
    port map (
            O => \N__44214\,
            I => n12482
        );

    \I__9332\ : InMux
    port map (
            O => \N__44211\,
            I => \N__44208\
        );

    \I__9331\ : LocalMux
    port map (
            O => \N__44208\,
            I => \N__44205\
        );

    \I__9330\ : Odrv4
    port map (
            O => \N__44205\,
            I => n14_adj_562
        );

    \I__9329\ : InMux
    port map (
            O => \N__44202\,
            I => \N__44198\
        );

    \I__9328\ : InMux
    port map (
            O => \N__44201\,
            I => \N__44195\
        );

    \I__9327\ : LocalMux
    port map (
            O => \N__44198\,
            I => \N__44192\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__44195\,
            I => \N__44189\
        );

    \I__9325\ : Span4Mux_v
    port map (
            O => \N__44192\,
            I => \N__44186\
        );

    \I__9324\ : Span4Mux_v
    port map (
            O => \N__44189\,
            I => \N__44181\
        );

    \I__9323\ : Span4Mux_h
    port map (
            O => \N__44186\,
            I => \N__44181\
        );

    \I__9322\ : Odrv4
    port map (
            O => \N__44181\,
            I => duty_11
        );

    \I__9321\ : InMux
    port map (
            O => \N__44178\,
            I => n12483
        );

    \I__9320\ : CascadeMux
    port map (
            O => \N__44175\,
            I => \N__44172\
        );

    \I__9319\ : InMux
    port map (
            O => \N__44172\,
            I => \N__44169\
        );

    \I__9318\ : LocalMux
    port map (
            O => \N__44169\,
            I => \N__44166\
        );

    \I__9317\ : Odrv4
    port map (
            O => \N__44166\,
            I => n13_adj_563
        );

    \I__9316\ : InMux
    port map (
            O => \N__44163\,
            I => n12484
        );

    \I__9315\ : InMux
    port map (
            O => \N__44160\,
            I => \N__44157\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__44157\,
            I => \N__44154\
        );

    \I__9313\ : Odrv12
    port map (
            O => \N__44154\,
            I => n12_adj_564
        );

    \I__9312\ : InMux
    port map (
            O => \N__44151\,
            I => \N__44147\
        );

    \I__9311\ : InMux
    port map (
            O => \N__44150\,
            I => \N__44144\
        );

    \I__9310\ : LocalMux
    port map (
            O => \N__44147\,
            I => \N__44139\
        );

    \I__9309\ : LocalMux
    port map (
            O => \N__44144\,
            I => \N__44139\
        );

    \I__9308\ : Span4Mux_v
    port map (
            O => \N__44139\,
            I => \N__44136\
        );

    \I__9307\ : Odrv4
    port map (
            O => \N__44136\,
            I => duty_13
        );

    \I__9306\ : InMux
    port map (
            O => \N__44133\,
            I => n12485
        );

    \I__9305\ : InMux
    port map (
            O => \N__44130\,
            I => \N__44127\
        );

    \I__9304\ : LocalMux
    port map (
            O => \N__44127\,
            I => \N__44124\
        );

    \I__9303\ : Odrv12
    port map (
            O => \N__44124\,
            I => n11_adj_565
        );

    \I__9302\ : InMux
    port map (
            O => \N__44121\,
            I => \N__44117\
        );

    \I__9301\ : InMux
    port map (
            O => \N__44120\,
            I => \N__44114\
        );

    \I__9300\ : LocalMux
    port map (
            O => \N__44117\,
            I => \N__44111\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__44114\,
            I => \N__44108\
        );

    \I__9298\ : Span4Mux_h
    port map (
            O => \N__44111\,
            I => \N__44105\
        );

    \I__9297\ : Span4Mux_v
    port map (
            O => \N__44108\,
            I => \N__44100\
        );

    \I__9296\ : Span4Mux_h
    port map (
            O => \N__44105\,
            I => \N__44100\
        );

    \I__9295\ : Odrv4
    port map (
            O => \N__44100\,
            I => duty_14
        );

    \I__9294\ : InMux
    port map (
            O => \N__44097\,
            I => n12486
        );

    \I__9293\ : InMux
    port map (
            O => \N__44094\,
            I => \N__44086\
        );

    \I__9292\ : InMux
    port map (
            O => \N__44093\,
            I => \N__44083\
        );

    \I__9291\ : InMux
    port map (
            O => \N__44092\,
            I => \N__44076\
        );

    \I__9290\ : InMux
    port map (
            O => \N__44091\,
            I => \N__44076\
        );

    \I__9289\ : InMux
    port map (
            O => \N__44090\,
            I => \N__44076\
        );

    \I__9288\ : InMux
    port map (
            O => \N__44089\,
            I => \N__44073\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__44086\,
            I => n861
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__44083\,
            I => n861
        );

    \I__9285\ : LocalMux
    port map (
            O => \N__44076\,
            I => n861
        );

    \I__9284\ : LocalMux
    port map (
            O => \N__44073\,
            I => n861
        );

    \I__9283\ : CascadeMux
    port map (
            O => \N__44064\,
            I => \N__44060\
        );

    \I__9282\ : CascadeMux
    port map (
            O => \N__44063\,
            I => \N__44057\
        );

    \I__9281\ : InMux
    port map (
            O => \N__44060\,
            I => \N__44054\
        );

    \I__9280\ : InMux
    port map (
            O => \N__44057\,
            I => \N__44051\
        );

    \I__9279\ : LocalMux
    port map (
            O => \N__44054\,
            I => n829
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__44051\,
            I => n829
        );

    \I__9277\ : InMux
    port map (
            O => \N__44046\,
            I => \N__44043\
        );

    \I__9276\ : LocalMux
    port map (
            O => \N__44043\,
            I => n896
        );

    \I__9275\ : InMux
    port map (
            O => \N__44040\,
            I => \bfn_12_25_0_\
        );

    \I__9274\ : InMux
    port map (
            O => \N__44037\,
            I => \N__44034\
        );

    \I__9273\ : LocalMux
    port map (
            O => \N__44034\,
            I => \N__44031\
        );

    \I__9272\ : Odrv4
    port map (
            O => \N__44031\,
            I => n24_adj_552
        );

    \I__9271\ : InMux
    port map (
            O => \N__44028\,
            I => n12473
        );

    \I__9270\ : InMux
    port map (
            O => \N__44025\,
            I => \N__44022\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__44022\,
            I => n23_adj_553
        );

    \I__9268\ : InMux
    port map (
            O => \N__44019\,
            I => n12474
        );

    \I__9267\ : InMux
    port map (
            O => \N__44016\,
            I => \N__44013\
        );

    \I__9266\ : LocalMux
    port map (
            O => \N__44013\,
            I => n22_adj_554
        );

    \I__9265\ : InMux
    port map (
            O => \N__44010\,
            I => n12475
        );

    \I__9264\ : InMux
    port map (
            O => \N__44007\,
            I => \N__44004\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__44004\,
            I => \N__44001\
        );

    \I__9262\ : Odrv4
    port map (
            O => \N__44001\,
            I => n21_adj_555
        );

    \I__9261\ : InMux
    port map (
            O => \N__43998\,
            I => \N__43995\
        );

    \I__9260\ : LocalMux
    port map (
            O => \N__43995\,
            I => \N__43992\
        );

    \I__9259\ : Span4Mux_v
    port map (
            O => \N__43992\,
            I => \N__43988\
        );

    \I__9258\ : InMux
    port map (
            O => \N__43991\,
            I => \N__43985\
        );

    \I__9257\ : Odrv4
    port map (
            O => \N__43988\,
            I => duty_4
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__43985\,
            I => duty_4
        );

    \I__9255\ : InMux
    port map (
            O => \N__43980\,
            I => n12476
        );

    \I__9254\ : InMux
    port map (
            O => \N__43977\,
            I => \N__43974\
        );

    \I__9253\ : LocalMux
    port map (
            O => \N__43974\,
            I => \N__43971\
        );

    \I__9252\ : Odrv4
    port map (
            O => \N__43971\,
            I => n20_adj_556
        );

    \I__9251\ : InMux
    port map (
            O => \N__43968\,
            I => \N__43965\
        );

    \I__9250\ : LocalMux
    port map (
            O => \N__43965\,
            I => \N__43962\
        );

    \I__9249\ : Span4Mux_v
    port map (
            O => \N__43962\,
            I => \N__43959\
        );

    \I__9248\ : Sp12to4
    port map (
            O => \N__43959\,
            I => \N__43955\
        );

    \I__9247\ : InMux
    port map (
            O => \N__43958\,
            I => \N__43952\
        );

    \I__9246\ : Odrv12
    port map (
            O => \N__43955\,
            I => duty_5
        );

    \I__9245\ : LocalMux
    port map (
            O => \N__43952\,
            I => duty_5
        );

    \I__9244\ : InMux
    port map (
            O => \N__43947\,
            I => n12477
        );

    \I__9243\ : InMux
    port map (
            O => \N__43944\,
            I => \N__43941\
        );

    \I__9242\ : LocalMux
    port map (
            O => \N__43941\,
            I => n19_adj_557
        );

    \I__9241\ : InMux
    port map (
            O => \N__43938\,
            I => n12478
        );

    \I__9240\ : InMux
    port map (
            O => \N__43935\,
            I => \N__43932\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__43932\,
            I => \N__43929\
        );

    \I__9238\ : Span4Mux_h
    port map (
            O => \N__43929\,
            I => \N__43926\
        );

    \I__9237\ : Span4Mux_h
    port map (
            O => \N__43926\,
            I => \N__43923\
        );

    \I__9236\ : Odrv4
    port map (
            O => \N__43923\,
            I => n18_adj_558
        );

    \I__9235\ : CascadeMux
    port map (
            O => \N__43920\,
            I => \N__43917\
        );

    \I__9234\ : InMux
    port map (
            O => \N__43917\,
            I => \N__43913\
        );

    \I__9233\ : InMux
    port map (
            O => \N__43916\,
            I => \N__43910\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__43913\,
            I => \N__43906\
        );

    \I__9231\ : LocalMux
    port map (
            O => \N__43910\,
            I => \N__43903\
        );

    \I__9230\ : InMux
    port map (
            O => \N__43909\,
            I => \N__43900\
        );

    \I__9229\ : Span4Mux_h
    port map (
            O => \N__43906\,
            I => \N__43897\
        );

    \I__9228\ : Span4Mux_v
    port map (
            O => \N__43903\,
            I => \N__43894\
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__43900\,
            I => encoder0_position_25
        );

    \I__9226\ : Odrv4
    port map (
            O => \N__43897\,
            I => encoder0_position_25
        );

    \I__9225\ : Odrv4
    port map (
            O => \N__43894\,
            I => encoder0_position_25
        );

    \I__9224\ : InMux
    port map (
            O => \N__43887\,
            I => \N__43884\
        );

    \I__9223\ : LocalMux
    port map (
            O => \N__43884\,
            I => \N__43881\
        );

    \I__9222\ : Span4Mux_h
    port map (
            O => \N__43881\,
            I => \N__43878\
        );

    \I__9221\ : Odrv4
    port map (
            O => \N__43878\,
            I => n8
        );

    \I__9220\ : InMux
    port map (
            O => \N__43875\,
            I => \N__43871\
        );

    \I__9219\ : InMux
    port map (
            O => \N__43874\,
            I => \N__43868\
        );

    \I__9218\ : LocalMux
    port map (
            O => \N__43871\,
            I => n41
        );

    \I__9217\ : LocalMux
    port map (
            O => \N__43868\,
            I => n41
        );

    \I__9216\ : InMux
    port map (
            O => \N__43863\,
            I => \N__43860\
        );

    \I__9215\ : LocalMux
    port map (
            O => \N__43860\,
            I => n901
        );

    \I__9214\ : CascadeMux
    port map (
            O => \N__43857\,
            I => \n41_cascade_\
        );

    \I__9213\ : CascadeMux
    port map (
            O => \N__43854\,
            I => \n933_cascade_\
        );

    \I__9212\ : CascadeMux
    port map (
            O => \N__43851\,
            I => \N__43848\
        );

    \I__9211\ : InMux
    port map (
            O => \N__43848\,
            I => \N__43845\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__43845\,
            I => \N__43842\
        );

    \I__9209\ : Odrv12
    port map (
            O => \N__43842\,
            I => n10
        );

    \I__9208\ : InMux
    port map (
            O => \N__43839\,
            I => \N__43834\
        );

    \I__9207\ : InMux
    port map (
            O => \N__43838\,
            I => \N__43831\
        );

    \I__9206\ : InMux
    port map (
            O => \N__43837\,
            I => \N__43828\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__43834\,
            I => \N__43825\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__43831\,
            I => \N__43822\
        );

    \I__9203\ : LocalMux
    port map (
            O => \N__43828\,
            I => \N__43817\
        );

    \I__9202\ : Span4Mux_v
    port map (
            O => \N__43825\,
            I => \N__43817\
        );

    \I__9201\ : Span4Mux_h
    port map (
            O => \N__43822\,
            I => \N__43814\
        );

    \I__9200\ : Odrv4
    port map (
            O => \N__43817\,
            I => encoder0_position_23
        );

    \I__9199\ : Odrv4
    port map (
            O => \N__43814\,
            I => encoder0_position_23
        );

    \I__9198\ : CascadeMux
    port map (
            O => \N__43809\,
            I => \N__43805\
        );

    \I__9197\ : InMux
    port map (
            O => \N__43808\,
            I => \N__43802\
        );

    \I__9196\ : InMux
    port map (
            O => \N__43805\,
            I => \N__43798\
        );

    \I__9195\ : LocalMux
    port map (
            O => \N__43802\,
            I => \N__43795\
        );

    \I__9194\ : InMux
    port map (
            O => \N__43801\,
            I => \N__43792\
        );

    \I__9193\ : LocalMux
    port map (
            O => \N__43798\,
            I => \N__43787\
        );

    \I__9192\ : Span4Mux_v
    port map (
            O => \N__43795\,
            I => \N__43787\
        );

    \I__9191\ : LocalMux
    port map (
            O => \N__43792\,
            I => \N__43784\
        );

    \I__9190\ : Odrv4
    port map (
            O => \N__43787\,
            I => encoder0_position_24
        );

    \I__9189\ : Odrv12
    port map (
            O => \N__43784\,
            I => encoder0_position_24
        );

    \I__9188\ : InMux
    port map (
            O => \N__43779\,
            I => \N__43776\
        );

    \I__9187\ : LocalMux
    port map (
            O => \N__43776\,
            I => \N__43773\
        );

    \I__9186\ : Span4Mux_v
    port map (
            O => \N__43773\,
            I => \N__43770\
        );

    \I__9185\ : Span4Mux_h
    port map (
            O => \N__43770\,
            I => \N__43767\
        );

    \I__9184\ : Odrv4
    port map (
            O => \N__43767\,
            I => n9
        );

    \I__9183\ : CascadeMux
    port map (
            O => \N__43764\,
            I => \n295_cascade_\
        );

    \I__9182\ : CascadeMux
    port map (
            O => \N__43761\,
            I => \n11955_cascade_\
        );

    \I__9181\ : InMux
    port map (
            O => \N__43758\,
            I => \N__43755\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__43755\,
            I => n14460
        );

    \I__9179\ : CascadeMux
    port map (
            O => \N__43752\,
            I => \n960_cascade_\
        );

    \I__9178\ : CascadeMux
    port map (
            O => \N__43749\,
            I => \N__43745\
        );

    \I__9177\ : InMux
    port map (
            O => \N__43748\,
            I => \N__43742\
        );

    \I__9176\ : InMux
    port map (
            O => \N__43745\,
            I => \N__43739\
        );

    \I__9175\ : LocalMux
    port map (
            O => \N__43742\,
            I => \N__43736\
        );

    \I__9174\ : LocalMux
    port map (
            O => \N__43739\,
            I => \N__43730\
        );

    \I__9173\ : Span4Mux_h
    port map (
            O => \N__43736\,
            I => \N__43730\
        );

    \I__9172\ : InMux
    port map (
            O => \N__43735\,
            I => \N__43727\
        );

    \I__9171\ : Span4Mux_v
    port map (
            O => \N__43730\,
            I => \N__43724\
        );

    \I__9170\ : LocalMux
    port map (
            O => \N__43727\,
            I => n1818
        );

    \I__9169\ : Odrv4
    port map (
            O => \N__43724\,
            I => n1818
        );

    \I__9168\ : CascadeMux
    port map (
            O => \N__43719\,
            I => \N__43716\
        );

    \I__9167\ : InMux
    port map (
            O => \N__43716\,
            I => \N__43713\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__43713\,
            I => \N__43710\
        );

    \I__9165\ : Span4Mux_v
    port map (
            O => \N__43710\,
            I => \N__43707\
        );

    \I__9164\ : Odrv4
    port map (
            O => \N__43707\,
            I => n10_adj_628
        );

    \I__9163\ : InMux
    port map (
            O => \N__43704\,
            I => \N__43701\
        );

    \I__9162\ : LocalMux
    port map (
            O => \N__43701\,
            I => \N__43698\
        );

    \I__9161\ : Span4Mux_h
    port map (
            O => \N__43698\,
            I => \N__43695\
        );

    \I__9160\ : Odrv4
    port map (
            O => \N__43695\,
            I => n17
        );

    \I__9159\ : InMux
    port map (
            O => \N__43692\,
            I => \N__43689\
        );

    \I__9158\ : LocalMux
    port map (
            O => \N__43689\,
            I => \N__43684\
        );

    \I__9157\ : InMux
    port map (
            O => \N__43688\,
            I => \N__43681\
        );

    \I__9156\ : InMux
    port map (
            O => \N__43687\,
            I => \N__43678\
        );

    \I__9155\ : Span4Mux_v
    port map (
            O => \N__43684\,
            I => \N__43671\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__43681\,
            I => \N__43671\
        );

    \I__9153\ : LocalMux
    port map (
            O => \N__43678\,
            I => \N__43671\
        );

    \I__9152\ : Odrv4
    port map (
            O => \N__43671\,
            I => n303
        );

    \I__9151\ : InMux
    port map (
            O => \N__43668\,
            I => \N__43665\
        );

    \I__9150\ : LocalMux
    port map (
            O => \N__43665\,
            I => \N__43662\
        );

    \I__9149\ : Span4Mux_v
    port map (
            O => \N__43662\,
            I => \N__43659\
        );

    \I__9148\ : Odrv4
    port map (
            O => \N__43659\,
            I => n15
        );

    \I__9147\ : CascadeMux
    port map (
            O => \N__43656\,
            I => \N__43652\
        );

    \I__9146\ : InMux
    port map (
            O => \N__43655\,
            I => \N__43649\
        );

    \I__9145\ : InMux
    port map (
            O => \N__43652\,
            I => \N__43645\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__43649\,
            I => \N__43642\
        );

    \I__9143\ : InMux
    port map (
            O => \N__43648\,
            I => \N__43639\
        );

    \I__9142\ : LocalMux
    port map (
            O => \N__43645\,
            I => \N__43634\
        );

    \I__9141\ : Span4Mux_v
    port map (
            O => \N__43642\,
            I => \N__43634\
        );

    \I__9140\ : LocalMux
    port map (
            O => \N__43639\,
            I => \N__43631\
        );

    \I__9139\ : Odrv4
    port map (
            O => \N__43634\,
            I => encoder0_position_18
        );

    \I__9138\ : Odrv12
    port map (
            O => \N__43631\,
            I => encoder0_position_18
        );

    \I__9137\ : InMux
    port map (
            O => \N__43626\,
            I => \N__43623\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__43623\,
            I => n899
        );

    \I__9135\ : CascadeMux
    port map (
            O => \N__43620\,
            I => \N__43616\
        );

    \I__9134\ : CascadeMux
    port map (
            O => \N__43619\,
            I => \N__43613\
        );

    \I__9133\ : InMux
    port map (
            O => \N__43616\,
            I => \N__43610\
        );

    \I__9132\ : InMux
    port map (
            O => \N__43613\,
            I => \N__43607\
        );

    \I__9131\ : LocalMux
    port map (
            O => \N__43610\,
            I => \N__43604\
        );

    \I__9130\ : LocalMux
    port map (
            O => \N__43607\,
            I => n832
        );

    \I__9129\ : Odrv4
    port map (
            O => \N__43604\,
            I => n832
        );

    \I__9128\ : InMux
    port map (
            O => \N__43599\,
            I => \N__43596\
        );

    \I__9127\ : LocalMux
    port map (
            O => \N__43596\,
            I => n900
        );

    \I__9126\ : CascadeMux
    port map (
            O => \N__43593\,
            I => \N__43589\
        );

    \I__9125\ : CascadeMux
    port map (
            O => \N__43592\,
            I => \N__43586\
        );

    \I__9124\ : InMux
    port map (
            O => \N__43589\,
            I => \N__43582\
        );

    \I__9123\ : InMux
    port map (
            O => \N__43586\,
            I => \N__43579\
        );

    \I__9122\ : InMux
    port map (
            O => \N__43585\,
            I => \N__43576\
        );

    \I__9121\ : LocalMux
    port map (
            O => \N__43582\,
            I => \N__43571\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__43579\,
            I => \N__43571\
        );

    \I__9119\ : LocalMux
    port map (
            O => \N__43576\,
            I => n833
        );

    \I__9118\ : Odrv4
    port map (
            O => \N__43571\,
            I => n833
        );

    \I__9117\ : CascadeMux
    port map (
            O => \N__43566\,
            I => \n932_cascade_\
        );

    \I__9116\ : InMux
    port map (
            O => \N__43563\,
            I => n12597
        );

    \I__9115\ : CascadeMux
    port map (
            O => \N__43560\,
            I => \N__43557\
        );

    \I__9114\ : InMux
    port map (
            O => \N__43557\,
            I => \N__43554\
        );

    \I__9113\ : LocalMux
    port map (
            O => \N__43554\,
            I => \N__43550\
        );

    \I__9112\ : InMux
    port map (
            O => \N__43553\,
            I => \N__43547\
        );

    \I__9111\ : Span4Mux_v
    port map (
            O => \N__43550\,
            I => \N__43544\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__43547\,
            I => n1726
        );

    \I__9109\ : Odrv4
    port map (
            O => \N__43544\,
            I => n1726
        );

    \I__9108\ : CascadeMux
    port map (
            O => \N__43539\,
            I => \N__43536\
        );

    \I__9107\ : InMux
    port map (
            O => \N__43536\,
            I => \N__43533\
        );

    \I__9106\ : LocalMux
    port map (
            O => \N__43533\,
            I => \N__43530\
        );

    \I__9105\ : Span4Mux_h
    port map (
            O => \N__43530\,
            I => \N__43527\
        );

    \I__9104\ : Odrv4
    port map (
            O => \N__43527\,
            I => n1793
        );

    \I__9103\ : InMux
    port map (
            O => \N__43524\,
            I => \bfn_12_21_0_\
        );

    \I__9102\ : InMux
    port map (
            O => \N__43521\,
            I => \N__43518\
        );

    \I__9101\ : LocalMux
    port map (
            O => \N__43518\,
            I => \N__43515\
        );

    \I__9100\ : Span4Mux_h
    port map (
            O => \N__43515\,
            I => \N__43512\
        );

    \I__9099\ : Odrv4
    port map (
            O => \N__43512\,
            I => n1792
        );

    \I__9098\ : InMux
    port map (
            O => \N__43509\,
            I => n12599
        );

    \I__9097\ : InMux
    port map (
            O => \N__43506\,
            I => \N__43503\
        );

    \I__9096\ : LocalMux
    port map (
            O => \N__43503\,
            I => \N__43500\
        );

    \I__9095\ : Span4Mux_h
    port map (
            O => \N__43500\,
            I => \N__43497\
        );

    \I__9094\ : Odrv4
    port map (
            O => \N__43497\,
            I => n1791
        );

    \I__9093\ : InMux
    port map (
            O => \N__43494\,
            I => n12600
        );

    \I__9092\ : CascadeMux
    port map (
            O => \N__43491\,
            I => \N__43488\
        );

    \I__9091\ : InMux
    port map (
            O => \N__43488\,
            I => \N__43484\
        );

    \I__9090\ : InMux
    port map (
            O => \N__43487\,
            I => \N__43480\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__43484\,
            I => \N__43477\
        );

    \I__9088\ : InMux
    port map (
            O => \N__43483\,
            I => \N__43474\
        );

    \I__9087\ : LocalMux
    port map (
            O => \N__43480\,
            I => n1723
        );

    \I__9086\ : Odrv4
    port map (
            O => \N__43477\,
            I => n1723
        );

    \I__9085\ : LocalMux
    port map (
            O => \N__43474\,
            I => n1723
        );

    \I__9084\ : InMux
    port map (
            O => \N__43467\,
            I => \N__43464\
        );

    \I__9083\ : LocalMux
    port map (
            O => \N__43464\,
            I => \N__43461\
        );

    \I__9082\ : Odrv4
    port map (
            O => \N__43461\,
            I => n1790
        );

    \I__9081\ : InMux
    port map (
            O => \N__43458\,
            I => n12601
        );

    \I__9080\ : CascadeMux
    port map (
            O => \N__43455\,
            I => \N__43452\
        );

    \I__9079\ : InMux
    port map (
            O => \N__43452\,
            I => \N__43449\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__43449\,
            I => \N__43445\
        );

    \I__9077\ : InMux
    port map (
            O => \N__43448\,
            I => \N__43442\
        );

    \I__9076\ : Odrv4
    port map (
            O => \N__43445\,
            I => n1722
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__43442\,
            I => n1722
        );

    \I__9074\ : InMux
    port map (
            O => \N__43437\,
            I => \N__43434\
        );

    \I__9073\ : LocalMux
    port map (
            O => \N__43434\,
            I => \N__43431\
        );

    \I__9072\ : Odrv4
    port map (
            O => \N__43431\,
            I => n1789
        );

    \I__9071\ : InMux
    port map (
            O => \N__43428\,
            I => n12602
        );

    \I__9070\ : CascadeMux
    port map (
            O => \N__43425\,
            I => \N__43422\
        );

    \I__9069\ : InMux
    port map (
            O => \N__43422\,
            I => \N__43419\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__43419\,
            I => \N__43415\
        );

    \I__9067\ : InMux
    port map (
            O => \N__43418\,
            I => \N__43412\
        );

    \I__9066\ : Odrv4
    port map (
            O => \N__43415\,
            I => n1721
        );

    \I__9065\ : LocalMux
    port map (
            O => \N__43412\,
            I => n1721
        );

    \I__9064\ : InMux
    port map (
            O => \N__43407\,
            I => \N__43404\
        );

    \I__9063\ : LocalMux
    port map (
            O => \N__43404\,
            I => \N__43401\
        );

    \I__9062\ : Odrv12
    port map (
            O => \N__43401\,
            I => n1788
        );

    \I__9061\ : InMux
    port map (
            O => \N__43398\,
            I => n12603
        );

    \I__9060\ : CascadeMux
    port map (
            O => \N__43395\,
            I => \N__43392\
        );

    \I__9059\ : InMux
    port map (
            O => \N__43392\,
            I => \N__43387\
        );

    \I__9058\ : InMux
    port map (
            O => \N__43391\,
            I => \N__43384\
        );

    \I__9057\ : InMux
    port map (
            O => \N__43390\,
            I => \N__43381\
        );

    \I__9056\ : LocalMux
    port map (
            O => \N__43387\,
            I => \N__43376\
        );

    \I__9055\ : LocalMux
    port map (
            O => \N__43384\,
            I => \N__43376\
        );

    \I__9054\ : LocalMux
    port map (
            O => \N__43381\,
            I => \N__43373\
        );

    \I__9053\ : Odrv4
    port map (
            O => \N__43376\,
            I => n1720
        );

    \I__9052\ : Odrv4
    port map (
            O => \N__43373\,
            I => n1720
        );

    \I__9051\ : InMux
    port map (
            O => \N__43368\,
            I => \N__43365\
        );

    \I__9050\ : LocalMux
    port map (
            O => \N__43365\,
            I => n1787
        );

    \I__9049\ : InMux
    port map (
            O => \N__43362\,
            I => n12604
        );

    \I__9048\ : InMux
    port map (
            O => \N__43359\,
            I => n12605
        );

    \I__9047\ : CascadeMux
    port map (
            O => \N__43356\,
            I => \n1731_cascade_\
        );

    \I__9046\ : InMux
    port map (
            O => \N__43353\,
            I => \N__43350\
        );

    \I__9045\ : LocalMux
    port map (
            O => \N__43350\,
            I => n11991
        );

    \I__9044\ : InMux
    port map (
            O => \N__43347\,
            I => \N__43344\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__43344\,
            I => \N__43341\
        );

    \I__9042\ : Span4Mux_h
    port map (
            O => \N__43341\,
            I => \N__43338\
        );

    \I__9041\ : Odrv4
    port map (
            O => \N__43338\,
            I => n1801
        );

    \I__9040\ : InMux
    port map (
            O => \N__43335\,
            I => \bfn_12_20_0_\
        );

    \I__9039\ : InMux
    port map (
            O => \N__43332\,
            I => \N__43329\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__43329\,
            I => \N__43326\
        );

    \I__9037\ : Span4Mux_h
    port map (
            O => \N__43326\,
            I => \N__43323\
        );

    \I__9036\ : Odrv4
    port map (
            O => \N__43323\,
            I => n1800
        );

    \I__9035\ : InMux
    port map (
            O => \N__43320\,
            I => n12591
        );

    \I__9034\ : CascadeMux
    port map (
            O => \N__43317\,
            I => \N__43314\
        );

    \I__9033\ : InMux
    port map (
            O => \N__43314\,
            I => \N__43311\
        );

    \I__9032\ : LocalMux
    port map (
            O => \N__43311\,
            I => \N__43307\
        );

    \I__9031\ : CascadeMux
    port map (
            O => \N__43310\,
            I => \N__43304\
        );

    \I__9030\ : Span4Mux_v
    port map (
            O => \N__43307\,
            I => \N__43300\
        );

    \I__9029\ : InMux
    port map (
            O => \N__43304\,
            I => \N__43297\
        );

    \I__9028\ : InMux
    port map (
            O => \N__43303\,
            I => \N__43294\
        );

    \I__9027\ : Odrv4
    port map (
            O => \N__43300\,
            I => n1732
        );

    \I__9026\ : LocalMux
    port map (
            O => \N__43297\,
            I => n1732
        );

    \I__9025\ : LocalMux
    port map (
            O => \N__43294\,
            I => n1732
        );

    \I__9024\ : InMux
    port map (
            O => \N__43287\,
            I => \N__43284\
        );

    \I__9023\ : LocalMux
    port map (
            O => \N__43284\,
            I => \N__43281\
        );

    \I__9022\ : Span4Mux_h
    port map (
            O => \N__43281\,
            I => \N__43278\
        );

    \I__9021\ : Odrv4
    port map (
            O => \N__43278\,
            I => n1799
        );

    \I__9020\ : InMux
    port map (
            O => \N__43275\,
            I => n12592
        );

    \I__9019\ : InMux
    port map (
            O => \N__43272\,
            I => \N__43268\
        );

    \I__9018\ : CascadeMux
    port map (
            O => \N__43271\,
            I => \N__43265\
        );

    \I__9017\ : LocalMux
    port map (
            O => \N__43268\,
            I => \N__43262\
        );

    \I__9016\ : InMux
    port map (
            O => \N__43265\,
            I => \N__43259\
        );

    \I__9015\ : Odrv4
    port map (
            O => \N__43262\,
            I => n1731
        );

    \I__9014\ : LocalMux
    port map (
            O => \N__43259\,
            I => n1731
        );

    \I__9013\ : InMux
    port map (
            O => \N__43254\,
            I => \N__43251\
        );

    \I__9012\ : LocalMux
    port map (
            O => \N__43251\,
            I => \N__43248\
        );

    \I__9011\ : Odrv4
    port map (
            O => \N__43248\,
            I => n1798
        );

    \I__9010\ : InMux
    port map (
            O => \N__43245\,
            I => n12593
        );

    \I__9009\ : InMux
    port map (
            O => \N__43242\,
            I => \N__43239\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__43239\,
            I => n1797
        );

    \I__9007\ : InMux
    port map (
            O => \N__43236\,
            I => n12594
        );

    \I__9006\ : InMux
    port map (
            O => \N__43233\,
            I => \N__43230\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__43230\,
            I => \N__43227\
        );

    \I__9004\ : Odrv4
    port map (
            O => \N__43227\,
            I => n1796
        );

    \I__9003\ : InMux
    port map (
            O => \N__43224\,
            I => n12595
        );

    \I__9002\ : CascadeMux
    port map (
            O => \N__43221\,
            I => \N__43218\
        );

    \I__9001\ : InMux
    port map (
            O => \N__43218\,
            I => \N__43215\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__43215\,
            I => \N__43212\
        );

    \I__8999\ : Odrv4
    port map (
            O => \N__43212\,
            I => n1795
        );

    \I__8998\ : InMux
    port map (
            O => \N__43209\,
            I => n12596
        );

    \I__8997\ : InMux
    port map (
            O => \N__43206\,
            I => \N__43203\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__43203\,
            I => \N__43200\
        );

    \I__8995\ : Odrv12
    port map (
            O => \N__43200\,
            I => n1794
        );

    \I__8994\ : CascadeMux
    port map (
            O => \N__43197\,
            I => \n1721_cascade_\
        );

    \I__8993\ : InMux
    port map (
            O => \N__43194\,
            I => \N__43190\
        );

    \I__8992\ : CascadeMux
    port map (
            O => \N__43193\,
            I => \N__43187\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__43190\,
            I => \N__43183\
        );

    \I__8990\ : InMux
    port map (
            O => \N__43187\,
            I => \N__43180\
        );

    \I__8989\ : InMux
    port map (
            O => \N__43186\,
            I => \N__43177\
        );

    \I__8988\ : Odrv4
    port map (
            O => \N__43183\,
            I => n1820
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__43180\,
            I => n1820
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__43177\,
            I => n1820
        );

    \I__8985\ : CascadeMux
    port map (
            O => \N__43170\,
            I => \N__43166\
        );

    \I__8984\ : CascadeMux
    port map (
            O => \N__43169\,
            I => \N__43163\
        );

    \I__8983\ : InMux
    port map (
            O => \N__43166\,
            I => \N__43159\
        );

    \I__8982\ : InMux
    port map (
            O => \N__43163\,
            I => \N__43156\
        );

    \I__8981\ : InMux
    port map (
            O => \N__43162\,
            I => \N__43153\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__43159\,
            I => n1827
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__43156\,
            I => n1827
        );

    \I__8978\ : LocalMux
    port map (
            O => \N__43153\,
            I => n1827
        );

    \I__8977\ : CascadeMux
    port map (
            O => \N__43146\,
            I => \n1722_cascade_\
        );

    \I__8976\ : CascadeMux
    port map (
            O => \N__43143\,
            I => \N__43139\
        );

    \I__8975\ : CascadeMux
    port map (
            O => \N__43142\,
            I => \N__43136\
        );

    \I__8974\ : InMux
    port map (
            O => \N__43139\,
            I => \N__43132\
        );

    \I__8973\ : InMux
    port map (
            O => \N__43136\,
            I => \N__43129\
        );

    \I__8972\ : InMux
    port map (
            O => \N__43135\,
            I => \N__43126\
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__43132\,
            I => n1821
        );

    \I__8970\ : LocalMux
    port map (
            O => \N__43129\,
            I => n1821
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__43126\,
            I => n1821
        );

    \I__8968\ : CascadeMux
    port map (
            O => \N__43119\,
            I => \N__43116\
        );

    \I__8967\ : InMux
    port map (
            O => \N__43116\,
            I => \N__43113\
        );

    \I__8966\ : LocalMux
    port map (
            O => \N__43113\,
            I => \N__43108\
        );

    \I__8965\ : InMux
    port map (
            O => \N__43112\,
            I => \N__43105\
        );

    \I__8964\ : CascadeMux
    port map (
            O => \N__43111\,
            I => \N__43102\
        );

    \I__8963\ : Span4Mux_h
    port map (
            O => \N__43108\,
            I => \N__43099\
        );

    \I__8962\ : LocalMux
    port map (
            O => \N__43105\,
            I => \N__43096\
        );

    \I__8961\ : InMux
    port map (
            O => \N__43102\,
            I => \N__43093\
        );

    \I__8960\ : Odrv4
    port map (
            O => \N__43099\,
            I => n1830
        );

    \I__8959\ : Odrv4
    port map (
            O => \N__43096\,
            I => n1830
        );

    \I__8958\ : LocalMux
    port map (
            O => \N__43093\,
            I => n1830
        );

    \I__8957\ : CascadeMux
    port map (
            O => \N__43086\,
            I => \n1752_cascade_\
        );

    \I__8956\ : InMux
    port map (
            O => \N__43083\,
            I => \N__43079\
        );

    \I__8955\ : CascadeMux
    port map (
            O => \N__43082\,
            I => \N__43076\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__43079\,
            I => \N__43072\
        );

    \I__8953\ : InMux
    port map (
            O => \N__43076\,
            I => \N__43069\
        );

    \I__8952\ : InMux
    port map (
            O => \N__43075\,
            I => \N__43066\
        );

    \I__8951\ : Odrv4
    port map (
            O => \N__43072\,
            I => n1826
        );

    \I__8950\ : LocalMux
    port map (
            O => \N__43069\,
            I => n1826
        );

    \I__8949\ : LocalMux
    port map (
            O => \N__43066\,
            I => n1826
        );

    \I__8948\ : CascadeMux
    port map (
            O => \N__43059\,
            I => \N__43054\
        );

    \I__8947\ : CascadeMux
    port map (
            O => \N__43058\,
            I => \N__43051\
        );

    \I__8946\ : InMux
    port map (
            O => \N__43057\,
            I => \N__43046\
        );

    \I__8945\ : InMux
    port map (
            O => \N__43054\,
            I => \N__43046\
        );

    \I__8944\ : InMux
    port map (
            O => \N__43051\,
            I => \N__43043\
        );

    \I__8943\ : LocalMux
    port map (
            O => \N__43046\,
            I => \N__43040\
        );

    \I__8942\ : LocalMux
    port map (
            O => \N__43043\,
            I => n1824
        );

    \I__8941\ : Odrv4
    port map (
            O => \N__43040\,
            I => n1824
        );

    \I__8940\ : CascadeMux
    port map (
            O => \N__43035\,
            I => \N__43032\
        );

    \I__8939\ : InMux
    port map (
            O => \N__43032\,
            I => \N__43028\
        );

    \I__8938\ : CascadeMux
    port map (
            O => \N__43031\,
            I => \N__43024\
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__43028\,
            I => \N__43021\
        );

    \I__8936\ : InMux
    port map (
            O => \N__43027\,
            I => \N__43018\
        );

    \I__8935\ : InMux
    port map (
            O => \N__43024\,
            I => \N__43015\
        );

    \I__8934\ : Span4Mux_h
    port map (
            O => \N__43021\,
            I => \N__43010\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__43018\,
            I => \N__43010\
        );

    \I__8932\ : LocalMux
    port map (
            O => \N__43015\,
            I => n1823
        );

    \I__8931\ : Odrv4
    port map (
            O => \N__43010\,
            I => n1823
        );

    \I__8930\ : CascadeMux
    port map (
            O => \N__43005\,
            I => \n1726_cascade_\
        );

    \I__8929\ : CascadeMux
    port map (
            O => \N__43002\,
            I => \n14244_cascade_\
        );

    \I__8928\ : CascadeMux
    port map (
            O => \N__42999\,
            I => \n14250_cascade_\
        );

    \I__8927\ : InMux
    port map (
            O => \N__42996\,
            I => \N__42993\
        );

    \I__8926\ : LocalMux
    port map (
            O => \N__42993\,
            I => n14254
        );

    \I__8925\ : InMux
    port map (
            O => \N__42990\,
            I => \N__42987\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__42987\,
            I => \N__42984\
        );

    \I__8923\ : Odrv12
    port map (
            O => \N__42984\,
            I => \pwm_setpoint_23_N_171_17\
        );

    \I__8922\ : InMux
    port map (
            O => \N__42981\,
            I => \N__42972\
        );

    \I__8921\ : InMux
    port map (
            O => \N__42980\,
            I => \N__42972\
        );

    \I__8920\ : InMux
    port map (
            O => \N__42979\,
            I => \N__42972\
        );

    \I__8919\ : LocalMux
    port map (
            O => \N__42972\,
            I => pwm_setpoint_16
        );

    \I__8918\ : CascadeMux
    port map (
            O => \N__42969\,
            I => \N__42966\
        );

    \I__8917\ : InMux
    port map (
            O => \N__42966\,
            I => \N__42961\
        );

    \I__8916\ : InMux
    port map (
            O => \N__42965\,
            I => \N__42958\
        );

    \I__8915\ : InMux
    port map (
            O => \N__42964\,
            I => \N__42955\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__42961\,
            I => \N__42952\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__42958\,
            I => \N__42947\
        );

    \I__8912\ : LocalMux
    port map (
            O => \N__42955\,
            I => \N__42947\
        );

    \I__8911\ : Span4Mux_s3_v
    port map (
            O => \N__42952\,
            I => \N__42942\
        );

    \I__8910\ : Span4Mux_s3_v
    port map (
            O => \N__42947\,
            I => \N__42942\
        );

    \I__8909\ : Odrv4
    port map (
            O => \N__42942\,
            I => pwm_setpoint_7
        );

    \I__8908\ : InMux
    port map (
            O => \N__42939\,
            I => \N__42936\
        );

    \I__8907\ : LocalMux
    port map (
            O => \N__42936\,
            I => \N__42933\
        );

    \I__8906\ : Odrv12
    port map (
            O => \N__42933\,
            I => \pwm_setpoint_23_N_171_10\
        );

    \I__8905\ : InMux
    port map (
            O => \N__42930\,
            I => \N__42926\
        );

    \I__8904\ : InMux
    port map (
            O => \N__42929\,
            I => \N__42923\
        );

    \I__8903\ : LocalMux
    port map (
            O => \N__42926\,
            I => \N__42920\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__42923\,
            I => \N__42917\
        );

    \I__8901\ : Span4Mux_s2_v
    port map (
            O => \N__42920\,
            I => \N__42914\
        );

    \I__8900\ : Span4Mux_h
    port map (
            O => \N__42917\,
            I => \N__42911\
        );

    \I__8899\ : Odrv4
    port map (
            O => \N__42914\,
            I => pwm_setpoint_11
        );

    \I__8898\ : Odrv4
    port map (
            O => \N__42911\,
            I => pwm_setpoint_11
        );

    \I__8897\ : InMux
    port map (
            O => \N__42906\,
            I => \N__42903\
        );

    \I__8896\ : LocalMux
    port map (
            O => \N__42903\,
            I => \N__42900\
        );

    \I__8895\ : Odrv4
    port map (
            O => \N__42900\,
            I => n15204
        );

    \I__8894\ : InMux
    port map (
            O => \N__42897\,
            I => \N__42891\
        );

    \I__8893\ : InMux
    port map (
            O => \N__42896\,
            I => \N__42891\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__42891\,
            I => pwm_setpoint_17
        );

    \I__8891\ : CascadeMux
    port map (
            O => \N__42888\,
            I => \n35_cascade_\
        );

    \I__8890\ : InMux
    port map (
            O => \N__42885\,
            I => \N__42882\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__42882\,
            I => n12_adj_661
        );

    \I__8888\ : InMux
    port map (
            O => \N__42879\,
            I => \N__42875\
        );

    \I__8887\ : CascadeMux
    port map (
            O => \N__42878\,
            I => \N__42872\
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__42875\,
            I => \N__42869\
        );

    \I__8885\ : InMux
    port map (
            O => \N__42872\,
            I => \N__42866\
        );

    \I__8884\ : Odrv4
    port map (
            O => \N__42869\,
            I => n1825
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__42866\,
            I => n1825
        );

    \I__8882\ : CascadeMux
    port map (
            O => \N__42861\,
            I => \n1825_cascade_\
        );

    \I__8881\ : InMux
    port map (
            O => \N__42858\,
            I => \N__42855\
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__42855\,
            I => \N__42852\
        );

    \I__8879\ : Odrv4
    port map (
            O => \N__42852\,
            I => n14520
        );

    \I__8878\ : InMux
    port map (
            O => \N__42849\,
            I => \N__42845\
        );

    \I__8877\ : CascadeMux
    port map (
            O => \N__42848\,
            I => \N__42842\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__42845\,
            I => \N__42838\
        );

    \I__8875\ : InMux
    port map (
            O => \N__42842\,
            I => \N__42835\
        );

    \I__8874\ : InMux
    port map (
            O => \N__42841\,
            I => \N__42832\
        );

    \I__8873\ : Odrv4
    port map (
            O => \N__42838\,
            I => n1828
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__42835\,
            I => n1828
        );

    \I__8871\ : LocalMux
    port map (
            O => \N__42832\,
            I => n1828
        );

    \I__8870\ : InMux
    port map (
            O => \N__42825\,
            I => \N__42822\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__42822\,
            I => \N__42819\
        );

    \I__8868\ : Odrv12
    port map (
            O => \N__42819\,
            I => \pwm_setpoint_23_N_171_22\
        );

    \I__8867\ : InMux
    port map (
            O => \N__42816\,
            I => \N__42810\
        );

    \I__8866\ : InMux
    port map (
            O => \N__42815\,
            I => \N__42810\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__42810\,
            I => \N__42807\
        );

    \I__8864\ : Odrv4
    port map (
            O => \N__42807\,
            I => n9_adj_658
        );

    \I__8863\ : InMux
    port map (
            O => \N__42804\,
            I => \N__42800\
        );

    \I__8862\ : InMux
    port map (
            O => \N__42803\,
            I => \N__42797\
        );

    \I__8861\ : LocalMux
    port map (
            O => \N__42800\,
            I => \N__42794\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__42797\,
            I => pwm_setpoint_8
        );

    \I__8859\ : Odrv4
    port map (
            O => \N__42794\,
            I => pwm_setpoint_8
        );

    \I__8858\ : CascadeMux
    port map (
            O => \N__42789\,
            I => \N__42786\
        );

    \I__8857\ : InMux
    port map (
            O => \N__42786\,
            I => \N__42783\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__42783\,
            I => n17_adj_665
        );

    \I__8855\ : InMux
    port map (
            O => \N__42780\,
            I => \N__42774\
        );

    \I__8854\ : InMux
    port map (
            O => \N__42779\,
            I => \N__42774\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__42774\,
            I => n19_adj_666
        );

    \I__8852\ : InMux
    port map (
            O => \N__42771\,
            I => \N__42768\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__42768\,
            I => n15178
        );

    \I__8850\ : CascadeMux
    port map (
            O => \N__42765\,
            I => \n17_adj_665_cascade_\
        );

    \I__8849\ : InMux
    port map (
            O => \N__42762\,
            I => \N__42759\
        );

    \I__8848\ : LocalMux
    port map (
            O => \N__42759\,
            I => \N__42756\
        );

    \I__8847\ : Odrv12
    port map (
            O => \N__42756\,
            I => \pwm_setpoint_23_N_171_16\
        );

    \I__8846\ : InMux
    port map (
            O => \N__42753\,
            I => \N__42750\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__42750\,
            I => n15174
        );

    \I__8844\ : CascadeMux
    port map (
            O => \N__42747\,
            I => \n16_adj_664_cascade_\
        );

    \I__8843\ : CascadeMux
    port map (
            O => \N__42744\,
            I => \n24_adj_669_cascade_\
        );

    \I__8842\ : InMux
    port map (
            O => \N__42741\,
            I => \N__42738\
        );

    \I__8841\ : LocalMux
    port map (
            O => \N__42738\,
            I => \N__42735\
        );

    \I__8840\ : Span4Mux_v
    port map (
            O => \N__42735\,
            I => \N__42732\
        );

    \I__8839\ : Odrv4
    port map (
            O => \N__42732\,
            I => n8_adj_657
        );

    \I__8838\ : InMux
    port map (
            O => \N__42729\,
            I => \N__42726\
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__42726\,
            I => n15144
        );

    \I__8836\ : InMux
    port map (
            O => \N__42723\,
            I => \N__42720\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__42720\,
            I => \pwm_setpoint_23_N_171_21\
        );

    \I__8834\ : CascadeMux
    port map (
            O => \N__42717\,
            I => \N__42714\
        );

    \I__8833\ : InMux
    port map (
            O => \N__42714\,
            I => \N__42711\
        );

    \I__8832\ : LocalMux
    port map (
            O => \N__42711\,
            I => \N__42708\
        );

    \I__8831\ : Odrv4
    port map (
            O => \N__42708\,
            I => \pwm_setpoint_23_N_171_9\
        );

    \I__8830\ : InMux
    port map (
            O => \N__42705\,
            I => \N__42696\
        );

    \I__8829\ : InMux
    port map (
            O => \N__42704\,
            I => \N__42696\
        );

    \I__8828\ : InMux
    port map (
            O => \N__42703\,
            I => \N__42696\
        );

    \I__8827\ : LocalMux
    port map (
            O => \N__42696\,
            I => pwm_setpoint_9
        );

    \I__8826\ : InMux
    port map (
            O => \N__42693\,
            I => \N__42690\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__42690\,
            I => \N__42687\
        );

    \I__8824\ : Odrv4
    port map (
            O => \N__42687\,
            I => \pwm_setpoint_23_N_171_14\
        );

    \I__8823\ : InMux
    port map (
            O => \N__42684\,
            I => \N__42681\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__42681\,
            I => \N__42678\
        );

    \I__8821\ : Odrv4
    port map (
            O => \N__42678\,
            I => n9_adj_581
        );

    \I__8820\ : InMux
    port map (
            O => \N__42675\,
            I => \bfn_11_28_0_\
        );

    \I__8819\ : InMux
    port map (
            O => \N__42672\,
            I => n12442
        );

    \I__8818\ : InMux
    port map (
            O => \N__42669\,
            I => \N__42666\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__42666\,
            I => \N__42663\
        );

    \I__8816\ : Span4Mux_v
    port map (
            O => \N__42663\,
            I => \N__42660\
        );

    \I__8815\ : Odrv4
    port map (
            O => \N__42660\,
            I => \pwm_setpoint_23_N_171_18\
        );

    \I__8814\ : InMux
    port map (
            O => \N__42657\,
            I => n12443
        );

    \I__8813\ : InMux
    port map (
            O => \N__42654\,
            I => n12444
        );

    \I__8812\ : InMux
    port map (
            O => \N__42651\,
            I => n12445
        );

    \I__8811\ : InMux
    port map (
            O => \N__42648\,
            I => n12446
        );

    \I__8810\ : InMux
    port map (
            O => \N__42645\,
            I => n12447
        );

    \I__8809\ : InMux
    port map (
            O => \N__42642\,
            I => n12448
        );

    \I__8808\ : InMux
    port map (
            O => \N__42639\,
            I => \N__42636\
        );

    \I__8807\ : LocalMux
    port map (
            O => \N__42636\,
            I => \N__42633\
        );

    \I__8806\ : Span4Mux_h
    port map (
            O => \N__42633\,
            I => \N__42630\
        );

    \I__8805\ : Odrv4
    port map (
            O => \N__42630\,
            I => n17_adj_589
        );

    \I__8804\ : InMux
    port map (
            O => \N__42627\,
            I => \N__42624\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__42624\,
            I => \pwm_setpoint_23_N_171_8\
        );

    \I__8802\ : InMux
    port map (
            O => \N__42621\,
            I => \bfn_11_27_0_\
        );

    \I__8801\ : InMux
    port map (
            O => \N__42618\,
            I => \N__42615\
        );

    \I__8800\ : LocalMux
    port map (
            O => \N__42615\,
            I => \N__42612\
        );

    \I__8799\ : Span4Mux_h
    port map (
            O => \N__42612\,
            I => \N__42609\
        );

    \I__8798\ : Odrv4
    port map (
            O => \N__42609\,
            I => n16_adj_588
        );

    \I__8797\ : InMux
    port map (
            O => \N__42606\,
            I => n12434
        );

    \I__8796\ : InMux
    port map (
            O => \N__42603\,
            I => \N__42600\
        );

    \I__8795\ : LocalMux
    port map (
            O => \N__42600\,
            I => \N__42597\
        );

    \I__8794\ : Span4Mux_h
    port map (
            O => \N__42597\,
            I => \N__42594\
        );

    \I__8793\ : Odrv4
    port map (
            O => \N__42594\,
            I => n15_adj_587
        );

    \I__8792\ : InMux
    port map (
            O => \N__42591\,
            I => n12435
        );

    \I__8791\ : InMux
    port map (
            O => \N__42588\,
            I => \N__42585\
        );

    \I__8790\ : LocalMux
    port map (
            O => \N__42585\,
            I => \N__42582\
        );

    \I__8789\ : Span4Mux_h
    port map (
            O => \N__42582\,
            I => \N__42579\
        );

    \I__8788\ : Odrv4
    port map (
            O => \N__42579\,
            I => n14_adj_586
        );

    \I__8787\ : InMux
    port map (
            O => \N__42576\,
            I => \N__42573\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__42573\,
            I => \pwm_setpoint_23_N_171_11\
        );

    \I__8785\ : InMux
    port map (
            O => \N__42570\,
            I => n12436
        );

    \I__8784\ : InMux
    port map (
            O => \N__42567\,
            I => n12437
        );

    \I__8783\ : InMux
    port map (
            O => \N__42564\,
            I => \N__42561\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__42561\,
            I => n12_adj_584
        );

    \I__8781\ : InMux
    port map (
            O => \N__42558\,
            I => \N__42555\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__42555\,
            I => \pwm_setpoint_23_N_171_13\
        );

    \I__8779\ : InMux
    port map (
            O => \N__42552\,
            I => n12438
        );

    \I__8778\ : InMux
    port map (
            O => \N__42549\,
            I => \N__42546\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__42546\,
            I => \N__42543\
        );

    \I__8776\ : Span4Mux_v
    port map (
            O => \N__42543\,
            I => \N__42540\
        );

    \I__8775\ : Odrv4
    port map (
            O => \N__42540\,
            I => n11_adj_583
        );

    \I__8774\ : InMux
    port map (
            O => \N__42537\,
            I => n12439
        );

    \I__8773\ : InMux
    port map (
            O => \N__42534\,
            I => \N__42531\
        );

    \I__8772\ : LocalMux
    port map (
            O => \N__42531\,
            I => \N__42528\
        );

    \I__8771\ : Span4Mux_h
    port map (
            O => \N__42528\,
            I => \N__42525\
        );

    \I__8770\ : Span4Mux_h
    port map (
            O => \N__42525\,
            I => \N__42522\
        );

    \I__8769\ : Span4Mux_h
    port map (
            O => \N__42522\,
            I => \N__42519\
        );

    \I__8768\ : Odrv4
    port map (
            O => \N__42519\,
            I => n10_adj_582
        );

    \I__8767\ : InMux
    port map (
            O => \N__42516\,
            I => n12440
        );

    \I__8766\ : InMux
    port map (
            O => \N__42513\,
            I => \N__42510\
        );

    \I__8765\ : LocalMux
    port map (
            O => \N__42510\,
            I => \N__42507\
        );

    \I__8764\ : Odrv12
    port map (
            O => \N__42507\,
            I => encoder0_position_scaled_2
        );

    \I__8763\ : InMux
    port map (
            O => \N__42504\,
            I => \N__42501\
        );

    \I__8762\ : LocalMux
    port map (
            O => \N__42501\,
            I => n25_adj_597
        );

    \I__8761\ : InMux
    port map (
            O => \N__42498\,
            I => \bfn_11_26_0_\
        );

    \I__8760\ : InMux
    port map (
            O => \N__42495\,
            I => n12426
        );

    \I__8759\ : InMux
    port map (
            O => \N__42492\,
            I => n12427
        );

    \I__8758\ : InMux
    port map (
            O => \N__42489\,
            I => \N__42486\
        );

    \I__8757\ : LocalMux
    port map (
            O => \N__42486\,
            I => n22_adj_594
        );

    \I__8756\ : InMux
    port map (
            O => \N__42483\,
            I => n12428
        );

    \I__8755\ : InMux
    port map (
            O => \N__42480\,
            I => \N__42477\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__42477\,
            I => n21_adj_593
        );

    \I__8753\ : InMux
    port map (
            O => \N__42474\,
            I => \N__42471\
        );

    \I__8752\ : LocalMux
    port map (
            O => \N__42471\,
            I => \pwm_setpoint_23_N_171_4\
        );

    \I__8751\ : InMux
    port map (
            O => \N__42468\,
            I => n12429
        );

    \I__8750\ : InMux
    port map (
            O => \N__42465\,
            I => \N__42462\
        );

    \I__8749\ : LocalMux
    port map (
            O => \N__42462\,
            I => n20_adj_592
        );

    \I__8748\ : InMux
    port map (
            O => \N__42459\,
            I => \N__42456\
        );

    \I__8747\ : LocalMux
    port map (
            O => \N__42456\,
            I => \pwm_setpoint_23_N_171_5\
        );

    \I__8746\ : InMux
    port map (
            O => \N__42453\,
            I => n12430
        );

    \I__8745\ : InMux
    port map (
            O => \N__42450\,
            I => n12431
        );

    \I__8744\ : InMux
    port map (
            O => \N__42447\,
            I => \N__42444\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__42444\,
            I => n18_adj_590
        );

    \I__8742\ : InMux
    port map (
            O => \N__42441\,
            I => \N__42438\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__42438\,
            I => \pwm_setpoint_23_N_171_7\
        );

    \I__8740\ : InMux
    port map (
            O => \N__42435\,
            I => n12432
        );

    \I__8739\ : InMux
    port map (
            O => \N__42432\,
            I => n12506
        );

    \I__8738\ : InMux
    port map (
            O => \N__42429\,
            I => \N__42424\
        );

    \I__8737\ : InMux
    port map (
            O => \N__42428\,
            I => \N__42421\
        );

    \I__8736\ : InMux
    port map (
            O => \N__42427\,
            I => \N__42418\
        );

    \I__8735\ : LocalMux
    port map (
            O => \N__42424\,
            I => \N__42415\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__42421\,
            I => \N__42410\
        );

    \I__8733\ : LocalMux
    port map (
            O => \N__42418\,
            I => \N__42410\
        );

    \I__8732\ : Span4Mux_h
    port map (
            O => \N__42415\,
            I => \N__42407\
        );

    \I__8731\ : Span4Mux_h
    port map (
            O => \N__42410\,
            I => \N__42404\
        );

    \I__8730\ : Odrv4
    port map (
            O => \N__42407\,
            I => n2
        );

    \I__8729\ : Odrv4
    port map (
            O => \N__42404\,
            I => n2
        );

    \I__8728\ : CascadeMux
    port map (
            O => \N__42399\,
            I => \N__42396\
        );

    \I__8727\ : InMux
    port map (
            O => \N__42396\,
            I => \N__42393\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__42393\,
            I => n14568
        );

    \I__8725\ : InMux
    port map (
            O => \N__42390\,
            I => \N__42387\
        );

    \I__8724\ : LocalMux
    port map (
            O => \N__42387\,
            I => \N__42384\
        );

    \I__8723\ : Odrv4
    port map (
            O => \N__42384\,
            I => n2561
        );

    \I__8722\ : CascadeMux
    port map (
            O => \N__42381\,
            I => \N__42378\
        );

    \I__8721\ : InMux
    port map (
            O => \N__42378\,
            I => \N__42374\
        );

    \I__8720\ : InMux
    port map (
            O => \N__42377\,
            I => \N__42371\
        );

    \I__8719\ : LocalMux
    port map (
            O => \N__42374\,
            I => n828
        );

    \I__8718\ : LocalMux
    port map (
            O => \N__42371\,
            I => n828
        );

    \I__8717\ : InMux
    port map (
            O => \N__42366\,
            I => \N__42363\
        );

    \I__8716\ : LocalMux
    port map (
            O => \N__42363\,
            I => \N__42360\
        );

    \I__8715\ : Odrv12
    port map (
            O => \N__42360\,
            I => encoder0_position_scaled_3
        );

    \I__8714\ : InMux
    port map (
            O => \N__42357\,
            I => \N__42354\
        );

    \I__8713\ : LocalMux
    port map (
            O => \N__42354\,
            I => \N__42351\
        );

    \I__8712\ : Odrv12
    port map (
            O => \N__42351\,
            I => encoder0_position_scaled_6
        );

    \I__8711\ : InMux
    port map (
            O => \N__42348\,
            I => \N__42344\
        );

    \I__8710\ : InMux
    port map (
            O => \N__42347\,
            I => \N__42341\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__42344\,
            I => \N__42337\
        );

    \I__8708\ : LocalMux
    port map (
            O => \N__42341\,
            I => \N__42334\
        );

    \I__8707\ : InMux
    port map (
            O => \N__42340\,
            I => \N__42331\
        );

    \I__8706\ : Span4Mux_v
    port map (
            O => \N__42337\,
            I => \N__42326\
        );

    \I__8705\ : Span4Mux_v
    port map (
            O => \N__42334\,
            I => \N__42326\
        );

    \I__8704\ : LocalMux
    port map (
            O => \N__42331\,
            I => \N__42323\
        );

    \I__8703\ : Odrv4
    port map (
            O => \N__42326\,
            I => n6
        );

    \I__8702\ : Odrv4
    port map (
            O => \N__42323\,
            I => n6
        );

    \I__8701\ : CascadeMux
    port map (
            O => \N__42318\,
            I => \N__42313\
        );

    \I__8700\ : InMux
    port map (
            O => \N__42317\,
            I => \N__42310\
        );

    \I__8699\ : InMux
    port map (
            O => \N__42316\,
            I => \N__42307\
        );

    \I__8698\ : InMux
    port map (
            O => \N__42313\,
            I => \N__42304\
        );

    \I__8697\ : LocalMux
    port map (
            O => \N__42310\,
            I => \N__42301\
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__42307\,
            I => \N__42298\
        );

    \I__8695\ : LocalMux
    port map (
            O => \N__42304\,
            I => \N__42295\
        );

    \I__8694\ : Span4Mux_h
    port map (
            O => \N__42301\,
            I => \N__42292\
        );

    \I__8693\ : Span4Mux_h
    port map (
            O => \N__42298\,
            I => \N__42289\
        );

    \I__8692\ : Odrv4
    port map (
            O => \N__42295\,
            I => n4
        );

    \I__8691\ : Odrv4
    port map (
            O => \N__42292\,
            I => n4
        );

    \I__8690\ : Odrv4
    port map (
            O => \N__42289\,
            I => n4
        );

    \I__8689\ : CascadeMux
    port map (
            O => \N__42282\,
            I => \N__42278\
        );

    \I__8688\ : CascadeMux
    port map (
            O => \N__42281\,
            I => \N__42275\
        );

    \I__8687\ : InMux
    port map (
            O => \N__42278\,
            I => \N__42272\
        );

    \I__8686\ : InMux
    port map (
            O => \N__42275\,
            I => \N__42269\
        );

    \I__8685\ : LocalMux
    port map (
            O => \N__42272\,
            I => n40
        );

    \I__8684\ : LocalMux
    port map (
            O => \N__42269\,
            I => n40
        );

    \I__8683\ : InMux
    port map (
            O => \N__42264\,
            I => \N__42260\
        );

    \I__8682\ : InMux
    port map (
            O => \N__42263\,
            I => \N__42257\
        );

    \I__8681\ : LocalMux
    port map (
            O => \N__42260\,
            I => \N__42253\
        );

    \I__8680\ : LocalMux
    port map (
            O => \N__42257\,
            I => \N__42250\
        );

    \I__8679\ : InMux
    port map (
            O => \N__42256\,
            I => \N__42247\
        );

    \I__8678\ : Span4Mux_v
    port map (
            O => \N__42253\,
            I => \N__42244\
        );

    \I__8677\ : Span4Mux_h
    port map (
            O => \N__42250\,
            I => \N__42241\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__42247\,
            I => \N__42238\
        );

    \I__8675\ : Odrv4
    port map (
            O => \N__42244\,
            I => n5
        );

    \I__8674\ : Odrv4
    port map (
            O => \N__42241\,
            I => n5
        );

    \I__8673\ : Odrv4
    port map (
            O => \N__42238\,
            I => n5
        );

    \I__8672\ : InMux
    port map (
            O => \N__42231\,
            I => \N__42228\
        );

    \I__8671\ : LocalMux
    port map (
            O => \N__42228\,
            I => n5_adj_682
        );

    \I__8670\ : CascadeMux
    port map (
            O => \N__42225\,
            I => \N__42222\
        );

    \I__8669\ : InMux
    port map (
            O => \N__42222\,
            I => \N__42212\
        );

    \I__8668\ : InMux
    port map (
            O => \N__42221\,
            I => \N__42212\
        );

    \I__8667\ : InMux
    port map (
            O => \N__42220\,
            I => \N__42212\
        );

    \I__8666\ : InMux
    port map (
            O => \N__42219\,
            I => \N__42209\
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__42212\,
            I => \N__42204\
        );

    \I__8664\ : LocalMux
    port map (
            O => \N__42209\,
            I => \N__42204\
        );

    \I__8663\ : Span4Mux_h
    port map (
            O => \N__42204\,
            I => \N__42201\
        );

    \I__8662\ : Odrv4
    port map (
            O => \N__42201\,
            I => n3
        );

    \I__8661\ : CascadeMux
    port map (
            O => \N__42198\,
            I => \n5_adj_682_cascade_\
        );

    \I__8660\ : CascadeMux
    port map (
            O => \N__42195\,
            I => \N__42190\
        );

    \I__8659\ : InMux
    port map (
            O => \N__42194\,
            I => \N__42185\
        );

    \I__8658\ : InMux
    port map (
            O => \N__42193\,
            I => \N__42182\
        );

    \I__8657\ : InMux
    port map (
            O => \N__42190\,
            I => \N__42175\
        );

    \I__8656\ : InMux
    port map (
            O => \N__42189\,
            I => \N__42175\
        );

    \I__8655\ : InMux
    port map (
            O => \N__42188\,
            I => \N__42175\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__42185\,
            I => n13653
        );

    \I__8653\ : LocalMux
    port map (
            O => \N__42182\,
            I => n13653
        );

    \I__8652\ : LocalMux
    port map (
            O => \N__42175\,
            I => n13653
        );

    \I__8651\ : InMux
    port map (
            O => \N__42168\,
            I => \bfn_11_24_0_\
        );

    \I__8650\ : InMux
    port map (
            O => \N__42165\,
            I => n12501
        );

    \I__8649\ : InMux
    port map (
            O => \N__42162\,
            I => n12502
        );

    \I__8648\ : CascadeMux
    port map (
            O => \N__42159\,
            I => \N__42156\
        );

    \I__8647\ : InMux
    port map (
            O => \N__42156\,
            I => \N__42152\
        );

    \I__8646\ : InMux
    port map (
            O => \N__42155\,
            I => \N__42148\
        );

    \I__8645\ : LocalMux
    port map (
            O => \N__42152\,
            I => \N__42145\
        );

    \I__8644\ : InMux
    port map (
            O => \N__42151\,
            I => \N__42142\
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__42148\,
            I => n831
        );

    \I__8642\ : Odrv4
    port map (
            O => \N__42145\,
            I => n831
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__42142\,
            I => n831
        );

    \I__8640\ : InMux
    port map (
            O => \N__42135\,
            I => \N__42132\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__42132\,
            I => n898
        );

    \I__8638\ : InMux
    port map (
            O => \N__42129\,
            I => n12503
        );

    \I__8637\ : CascadeMux
    port map (
            O => \N__42126\,
            I => \N__42122\
        );

    \I__8636\ : CascadeMux
    port map (
            O => \N__42125\,
            I => \N__42119\
        );

    \I__8635\ : InMux
    port map (
            O => \N__42122\,
            I => \N__42115\
        );

    \I__8634\ : InMux
    port map (
            O => \N__42119\,
            I => \N__42112\
        );

    \I__8633\ : InMux
    port map (
            O => \N__42118\,
            I => \N__42109\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__42115\,
            I => \N__42106\
        );

    \I__8631\ : LocalMux
    port map (
            O => \N__42112\,
            I => n830
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__42109\,
            I => n830
        );

    \I__8629\ : Odrv4
    port map (
            O => \N__42106\,
            I => n830
        );

    \I__8628\ : InMux
    port map (
            O => \N__42099\,
            I => \N__42096\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__42096\,
            I => n897
        );

    \I__8626\ : InMux
    port map (
            O => \N__42093\,
            I => n12504
        );

    \I__8625\ : InMux
    port map (
            O => \N__42090\,
            I => n12505
        );

    \I__8624\ : CascadeMux
    port map (
            O => \N__42087\,
            I => \n832_cascade_\
        );

    \I__8623\ : InMux
    port map (
            O => \N__42084\,
            I => \N__42081\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__42081\,
            I => n2564
        );

    \I__8621\ : CascadeMux
    port map (
            O => \N__42078\,
            I => \n13658_cascade_\
        );

    \I__8620\ : CascadeMux
    port map (
            O => \N__42075\,
            I => \N__42070\
        );

    \I__8619\ : CascadeMux
    port map (
            O => \N__42074\,
            I => \N__42067\
        );

    \I__8618\ : CascadeMux
    port map (
            O => \N__42073\,
            I => \N__42064\
        );

    \I__8617\ : InMux
    port map (
            O => \N__42070\,
            I => \N__42060\
        );

    \I__8616\ : InMux
    port map (
            O => \N__42067\,
            I => \N__42057\
        );

    \I__8615\ : InMux
    port map (
            O => \N__42064\,
            I => \N__42054\
        );

    \I__8614\ : InMux
    port map (
            O => \N__42063\,
            I => \N__42051\
        );

    \I__8613\ : LocalMux
    port map (
            O => \N__42060\,
            I => \N__42048\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__42057\,
            I => \N__42045\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__42054\,
            I => encoder0_position_28
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__42051\,
            I => encoder0_position_28
        );

    \I__8609\ : Odrv4
    port map (
            O => \N__42048\,
            I => encoder0_position_28
        );

    \I__8608\ : Odrv12
    port map (
            O => \N__42045\,
            I => encoder0_position_28
        );

    \I__8607\ : InMux
    port map (
            O => \N__42036\,
            I => \N__42033\
        );

    \I__8606\ : LocalMux
    port map (
            O => \N__42033\,
            I => \N__42030\
        );

    \I__8605\ : Span4Mux_v
    port map (
            O => \N__42030\,
            I => \N__42027\
        );

    \I__8604\ : Odrv4
    port map (
            O => \N__42027\,
            I => encoder0_position_scaled_4
        );

    \I__8603\ : CascadeMux
    port map (
            O => \N__42024\,
            I => \n929_cascade_\
        );

    \I__8602\ : CascadeMux
    port map (
            O => \N__42021\,
            I => \N__42016\
        );

    \I__8601\ : CascadeMux
    port map (
            O => \N__42020\,
            I => \N__42013\
        );

    \I__8600\ : CascadeMux
    port map (
            O => \N__42019\,
            I => \N__42010\
        );

    \I__8599\ : InMux
    port map (
            O => \N__42016\,
            I => \N__42007\
        );

    \I__8598\ : InMux
    port map (
            O => \N__42013\,
            I => \N__42004\
        );

    \I__8597\ : InMux
    port map (
            O => \N__42010\,
            I => \N__42000\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__42007\,
            I => \N__41995\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__42004\,
            I => \N__41995\
        );

    \I__8594\ : InMux
    port map (
            O => \N__42003\,
            I => \N__41992\
        );

    \I__8593\ : LocalMux
    port map (
            O => \N__42000\,
            I => encoder0_position_30
        );

    \I__8592\ : Odrv4
    port map (
            O => \N__41995\,
            I => encoder0_position_30
        );

    \I__8591\ : LocalMux
    port map (
            O => \N__41992\,
            I => encoder0_position_30
        );

    \I__8590\ : InMux
    port map (
            O => \N__41985\,
            I => \N__41982\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__41982\,
            I => n13654
        );

    \I__8588\ : CascadeMux
    port map (
            O => \N__41979\,
            I => \n829_cascade_\
        );

    \I__8587\ : InMux
    port map (
            O => \N__41976\,
            I => \N__41973\
        );

    \I__8586\ : LocalMux
    port map (
            O => \N__41973\,
            I => n12027
        );

    \I__8585\ : CascadeMux
    port map (
            O => \N__41970\,
            I => \n861_cascade_\
        );

    \I__8584\ : InMux
    port map (
            O => \N__41967\,
            I => \N__41964\
        );

    \I__8583\ : LocalMux
    port map (
            O => \N__41964\,
            I => \N__41961\
        );

    \I__8582\ : Span4Mux_h
    port map (
            O => \N__41961\,
            I => \N__41958\
        );

    \I__8581\ : Odrv4
    port map (
            O => \N__41958\,
            I => n16
        );

    \I__8580\ : CascadeMux
    port map (
            O => \N__41955\,
            I => \N__41951\
        );

    \I__8579\ : InMux
    port map (
            O => \N__41954\,
            I => \N__41946\
        );

    \I__8578\ : InMux
    port map (
            O => \N__41951\,
            I => \N__41943\
        );

    \I__8577\ : InMux
    port map (
            O => \N__41950\,
            I => \N__41940\
        );

    \I__8576\ : InMux
    port map (
            O => \N__41949\,
            I => \N__41937\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__41946\,
            I => encoder0_position_29
        );

    \I__8574\ : LocalMux
    port map (
            O => \N__41943\,
            I => encoder0_position_29
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__41940\,
            I => encoder0_position_29
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__41937\,
            I => encoder0_position_29
        );

    \I__8571\ : CascadeMux
    port map (
            O => \N__41928\,
            I => \N__41925\
        );

    \I__8570\ : InMux
    port map (
            O => \N__41925\,
            I => \N__41922\
        );

    \I__8569\ : LocalMux
    port map (
            O => \N__41922\,
            I => n404
        );

    \I__8568\ : InMux
    port map (
            O => \N__41919\,
            I => \N__41914\
        );

    \I__8567\ : InMux
    port map (
            O => \N__41918\,
            I => \N__41909\
        );

    \I__8566\ : InMux
    port map (
            O => \N__41917\,
            I => \N__41909\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__41914\,
            I => encoder0_position_17
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__41909\,
            I => encoder0_position_17
        );

    \I__8563\ : CascadeMux
    port map (
            O => \N__41904\,
            I => \N__41901\
        );

    \I__8562\ : InMux
    port map (
            O => \N__41901\,
            I => \N__41898\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__41898\,
            I => \N__41895\
        );

    \I__8560\ : Span4Mux_h
    port map (
            O => \N__41895\,
            I => \N__41892\
        );

    \I__8559\ : Odrv4
    port map (
            O => \N__41892\,
            I => n16_adj_634
        );

    \I__8558\ : CascadeMux
    port map (
            O => \N__41889\,
            I => \N__41886\
        );

    \I__8557\ : InMux
    port map (
            O => \N__41886\,
            I => \N__41883\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__41883\,
            I => \N__41880\
        );

    \I__8555\ : Span4Mux_v
    port map (
            O => \N__41880\,
            I => \N__41877\
        );

    \I__8554\ : Odrv4
    port map (
            O => \N__41877\,
            I => n7_adj_625
        );

    \I__8553\ : CascadeMux
    port map (
            O => \N__41874\,
            I => \N__41871\
        );

    \I__8552\ : InMux
    port map (
            O => \N__41871\,
            I => \N__41868\
        );

    \I__8551\ : LocalMux
    port map (
            O => \N__41868\,
            I => \N__41865\
        );

    \I__8550\ : Span4Mux_v
    port map (
            O => \N__41865\,
            I => \N__41862\
        );

    \I__8549\ : Odrv4
    port map (
            O => \N__41862\,
            I => n3_adj_621
        );

    \I__8548\ : InMux
    port map (
            O => \N__41859\,
            I => \N__41856\
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__41856\,
            I => n2566
        );

    \I__8546\ : CascadeMux
    port map (
            O => \N__41853\,
            I => \N__41850\
        );

    \I__8545\ : InMux
    port map (
            O => \N__41850\,
            I => \N__41847\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__41847\,
            I => \N__41843\
        );

    \I__8543\ : InMux
    port map (
            O => \N__41846\,
            I => \N__41840\
        );

    \I__8542\ : Span4Mux_h
    port map (
            O => \N__41843\,
            I => \N__41835\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__41840\,
            I => \N__41835\
        );

    \I__8540\ : Odrv4
    port map (
            O => \N__41835\,
            I => n7
        );

    \I__8539\ : CascadeMux
    port map (
            O => \N__41832\,
            I => \n13662_cascade_\
        );

    \I__8538\ : CascadeMux
    port map (
            O => \N__41829\,
            I => \N__41825\
        );

    \I__8537\ : CascadeMux
    port map (
            O => \N__41828\,
            I => \N__41822\
        );

    \I__8536\ : InMux
    port map (
            O => \N__41825\,
            I => \N__41818\
        );

    \I__8535\ : InMux
    port map (
            O => \N__41822\,
            I => \N__41814\
        );

    \I__8534\ : InMux
    port map (
            O => \N__41821\,
            I => \N__41811\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__41818\,
            I => \N__41808\
        );

    \I__8532\ : InMux
    port map (
            O => \N__41817\,
            I => \N__41805\
        );

    \I__8531\ : LocalMux
    port map (
            O => \N__41814\,
            I => encoder0_position_26
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__41811\,
            I => encoder0_position_26
        );

    \I__8529\ : Odrv4
    port map (
            O => \N__41808\,
            I => encoder0_position_26
        );

    \I__8528\ : LocalMux
    port map (
            O => \N__41805\,
            I => encoder0_position_26
        );

    \I__8527\ : CascadeMux
    port map (
            O => \N__41796\,
            I => \N__41793\
        );

    \I__8526\ : InMux
    port map (
            O => \N__41793\,
            I => \N__41790\
        );

    \I__8525\ : LocalMux
    port map (
            O => \N__41790\,
            I => n2565
        );

    \I__8524\ : InMux
    port map (
            O => \N__41787\,
            I => \N__41781\
        );

    \I__8523\ : InMux
    port map (
            O => \N__41786\,
            I => \N__41778\
        );

    \I__8522\ : InMux
    port map (
            O => \N__41785\,
            I => \N__41775\
        );

    \I__8521\ : InMux
    port map (
            O => \N__41784\,
            I => \N__41772\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__41781\,
            I => \N__41767\
        );

    \I__8519\ : LocalMux
    port map (
            O => \N__41778\,
            I => \N__41767\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__41775\,
            I => encoder0_position_27
        );

    \I__8517\ : LocalMux
    port map (
            O => \N__41772\,
            I => encoder0_position_27
        );

    \I__8516\ : Odrv4
    port map (
            O => \N__41767\,
            I => encoder0_position_27
        );

    \I__8515\ : CascadeMux
    port map (
            O => \N__41760\,
            I => \n13660_cascade_\
        );

    \I__8514\ : CascadeMux
    port map (
            O => \N__41757\,
            I => \N__41754\
        );

    \I__8513\ : InMux
    port map (
            O => \N__41754\,
            I => \N__41751\
        );

    \I__8512\ : LocalMux
    port map (
            O => \N__41751\,
            I => \N__41748\
        );

    \I__8511\ : Odrv4
    port map (
            O => \N__41748\,
            I => n1895
        );

    \I__8510\ : CascadeMux
    port map (
            O => \N__41745\,
            I => \N__41741\
        );

    \I__8509\ : CascadeMux
    port map (
            O => \N__41744\,
            I => \N__41738\
        );

    \I__8508\ : InMux
    port map (
            O => \N__41741\,
            I => \N__41735\
        );

    \I__8507\ : InMux
    port map (
            O => \N__41738\,
            I => \N__41732\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__41735\,
            I => \N__41729\
        );

    \I__8505\ : LocalMux
    port map (
            O => \N__41732\,
            I => \N__41726\
        );

    \I__8504\ : Span4Mux_h
    port map (
            O => \N__41729\,
            I => \N__41720\
        );

    \I__8503\ : Span4Mux_v
    port map (
            O => \N__41726\,
            I => \N__41720\
        );

    \I__8502\ : InMux
    port map (
            O => \N__41725\,
            I => \N__41717\
        );

    \I__8501\ : Odrv4
    port map (
            O => \N__41720\,
            I => n1927
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__41717\,
            I => n1927
        );

    \I__8499\ : InMux
    port map (
            O => \N__41712\,
            I => \N__41709\
        );

    \I__8498\ : LocalMux
    port map (
            O => \N__41709\,
            I => \N__41706\
        );

    \I__8497\ : Odrv4
    port map (
            O => \N__41706\,
            I => n1894
        );

    \I__8496\ : CascadeMux
    port map (
            O => \N__41703\,
            I => \N__41699\
        );

    \I__8495\ : CascadeMux
    port map (
            O => \N__41702\,
            I => \N__41696\
        );

    \I__8494\ : InMux
    port map (
            O => \N__41699\,
            I => \N__41693\
        );

    \I__8493\ : InMux
    port map (
            O => \N__41696\,
            I => \N__41690\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__41693\,
            I => \N__41687\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__41690\,
            I => \N__41684\
        );

    \I__8490\ : Span4Mux_h
    port map (
            O => \N__41687\,
            I => \N__41680\
        );

    \I__8489\ : Span4Mux_h
    port map (
            O => \N__41684\,
            I => \N__41677\
        );

    \I__8488\ : InMux
    port map (
            O => \N__41683\,
            I => \N__41674\
        );

    \I__8487\ : Odrv4
    port map (
            O => \N__41680\,
            I => n1926
        );

    \I__8486\ : Odrv4
    port map (
            O => \N__41677\,
            I => n1926
        );

    \I__8485\ : LocalMux
    port map (
            O => \N__41674\,
            I => n1926
        );

    \I__8484\ : CascadeMux
    port map (
            O => \N__41667\,
            I => \N__41662\
        );

    \I__8483\ : InMux
    port map (
            O => \N__41666\,
            I => \N__41657\
        );

    \I__8482\ : InMux
    port map (
            O => \N__41665\,
            I => \N__41657\
        );

    \I__8481\ : InMux
    port map (
            O => \N__41662\,
            I => \N__41654\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__41657\,
            I => \N__41649\
        );

    \I__8479\ : LocalMux
    port map (
            O => \N__41654\,
            I => \N__41649\
        );

    \I__8478\ : Odrv4
    port map (
            O => \N__41649\,
            I => n1829
        );

    \I__8477\ : CascadeMux
    port map (
            O => \N__41646\,
            I => \N__41643\
        );

    \I__8476\ : InMux
    port map (
            O => \N__41643\,
            I => \N__41640\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__41640\,
            I => n1885
        );

    \I__8474\ : InMux
    port map (
            O => \N__41637\,
            I => \N__41633\
        );

    \I__8473\ : InMux
    port map (
            O => \N__41636\,
            I => \N__41630\
        );

    \I__8472\ : LocalMux
    port map (
            O => \N__41633\,
            I => \N__41627\
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__41630\,
            I => \N__41624\
        );

    \I__8470\ : Span4Mux_v
    port map (
            O => \N__41627\,
            I => \N__41621\
        );

    \I__8469\ : Span4Mux_v
    port map (
            O => \N__41624\,
            I => \N__41618\
        );

    \I__8468\ : Odrv4
    port map (
            O => \N__41621\,
            I => n1917
        );

    \I__8467\ : Odrv4
    port map (
            O => \N__41618\,
            I => n1917
        );

    \I__8466\ : InMux
    port map (
            O => \N__41613\,
            I => \N__41610\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__41610\,
            I => \N__41607\
        );

    \I__8464\ : Span4Mux_v
    port map (
            O => \N__41607\,
            I => \N__41604\
        );

    \I__8463\ : Odrv4
    port map (
            O => \N__41604\,
            I => n30
        );

    \I__8462\ : CascadeMux
    port map (
            O => \N__41601\,
            I => \N__41597\
        );

    \I__8461\ : CascadeMux
    port map (
            O => \N__41600\,
            I => \N__41593\
        );

    \I__8460\ : InMux
    port map (
            O => \N__41597\,
            I => \N__41590\
        );

    \I__8459\ : InMux
    port map (
            O => \N__41596\,
            I => \N__41587\
        );

    \I__8458\ : InMux
    port map (
            O => \N__41593\,
            I => \N__41584\
        );

    \I__8457\ : LocalMux
    port map (
            O => \N__41590\,
            I => \N__41581\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__41587\,
            I => \N__41578\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__41584\,
            I => encoder0_position_3
        );

    \I__8454\ : Odrv4
    port map (
            O => \N__41581\,
            I => encoder0_position_3
        );

    \I__8453\ : Odrv4
    port map (
            O => \N__41578\,
            I => encoder0_position_3
        );

    \I__8452\ : InMux
    port map (
            O => \N__41571\,
            I => \N__41567\
        );

    \I__8451\ : InMux
    port map (
            O => \N__41570\,
            I => \N__41564\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__41567\,
            I => \N__41560\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__41564\,
            I => \N__41557\
        );

    \I__8448\ : InMux
    port map (
            O => \N__41563\,
            I => \N__41554\
        );

    \I__8447\ : Span4Mux_v
    port map (
            O => \N__41560\,
            I => \N__41551\
        );

    \I__8446\ : Span4Mux_s3_h
    port map (
            O => \N__41557\,
            I => \N__41546\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__41554\,
            I => \N__41546\
        );

    \I__8444\ : Span4Mux_h
    port map (
            O => \N__41551\,
            I => \N__41541\
        );

    \I__8443\ : Span4Mux_h
    port map (
            O => \N__41546\,
            I => \N__41541\
        );

    \I__8442\ : Span4Mux_v
    port map (
            O => \N__41541\,
            I => \N__41538\
        );

    \I__8441\ : Span4Mux_v
    port map (
            O => \N__41538\,
            I => \N__41535\
        );

    \I__8440\ : Odrv4
    port map (
            O => \N__41535\,
            I => n316
        );

    \I__8439\ : InMux
    port map (
            O => \N__41532\,
            I => \N__41529\
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__41529\,
            I => \N__41526\
        );

    \I__8437\ : Odrv4
    port map (
            O => \N__41526\,
            I => n1888
        );

    \I__8436\ : InMux
    port map (
            O => \N__41523\,
            I => \N__41520\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__41520\,
            I => \N__41516\
        );

    \I__8434\ : InMux
    port map (
            O => \N__41519\,
            I => \N__41509\
        );

    \I__8433\ : Span4Mux_v
    port map (
            O => \N__41516\,
            I => \N__41506\
        );

    \I__8432\ : InMux
    port map (
            O => \N__41515\,
            I => \N__41498\
        );

    \I__8431\ : CascadeMux
    port map (
            O => \N__41514\,
            I => \N__41491\
        );

    \I__8430\ : CascadeMux
    port map (
            O => \N__41513\,
            I => \N__41486\
        );

    \I__8429\ : CascadeMux
    port map (
            O => \N__41512\,
            I => \N__41483\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__41509\,
            I => \N__41477\
        );

    \I__8427\ : Span4Mux_v
    port map (
            O => \N__41506\,
            I => \N__41477\
        );

    \I__8426\ : InMux
    port map (
            O => \N__41505\,
            I => \N__41472\
        );

    \I__8425\ : InMux
    port map (
            O => \N__41504\,
            I => \N__41472\
        );

    \I__8424\ : InMux
    port map (
            O => \N__41503\,
            I => \N__41465\
        );

    \I__8423\ : InMux
    port map (
            O => \N__41502\,
            I => \N__41465\
        );

    \I__8422\ : InMux
    port map (
            O => \N__41501\,
            I => \N__41465\
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__41498\,
            I => \N__41462\
        );

    \I__8420\ : InMux
    port map (
            O => \N__41497\,
            I => \N__41455\
        );

    \I__8419\ : InMux
    port map (
            O => \N__41496\,
            I => \N__41455\
        );

    \I__8418\ : InMux
    port map (
            O => \N__41495\,
            I => \N__41455\
        );

    \I__8417\ : InMux
    port map (
            O => \N__41494\,
            I => \N__41446\
        );

    \I__8416\ : InMux
    port map (
            O => \N__41491\,
            I => \N__41446\
        );

    \I__8415\ : InMux
    port map (
            O => \N__41490\,
            I => \N__41446\
        );

    \I__8414\ : InMux
    port map (
            O => \N__41489\,
            I => \N__41446\
        );

    \I__8413\ : InMux
    port map (
            O => \N__41486\,
            I => \N__41439\
        );

    \I__8412\ : InMux
    port map (
            O => \N__41483\,
            I => \N__41439\
        );

    \I__8411\ : InMux
    port map (
            O => \N__41482\,
            I => \N__41439\
        );

    \I__8410\ : Span4Mux_h
    port map (
            O => \N__41477\,
            I => \N__41432\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__41472\,
            I => \N__41432\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__41465\,
            I => \N__41432\
        );

    \I__8407\ : Odrv4
    port map (
            O => \N__41462\,
            I => n1851
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__41455\,
            I => n1851
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__41446\,
            I => n1851
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__41439\,
            I => n1851
        );

    \I__8403\ : Odrv4
    port map (
            O => \N__41432\,
            I => n1851
        );

    \I__8402\ : InMux
    port map (
            O => \N__41421\,
            I => \N__41417\
        );

    \I__8401\ : InMux
    port map (
            O => \N__41420\,
            I => \N__41414\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__41417\,
            I => \N__41411\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__41414\,
            I => \N__41408\
        );

    \I__8398\ : Span4Mux_h
    port map (
            O => \N__41411\,
            I => \N__41405\
        );

    \I__8397\ : Span4Mux_h
    port map (
            O => \N__41408\,
            I => \N__41402\
        );

    \I__8396\ : Odrv4
    port map (
            O => \N__41405\,
            I => n1920
        );

    \I__8395\ : Odrv4
    port map (
            O => \N__41402\,
            I => n1920
        );

    \I__8394\ : InMux
    port map (
            O => \N__41397\,
            I => \N__41394\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__41394\,
            I => \N__41391\
        );

    \I__8392\ : Span4Mux_h
    port map (
            O => \N__41391\,
            I => \N__41388\
        );

    \I__8391\ : Odrv4
    port map (
            O => \N__41388\,
            I => n1987
        );

    \I__8390\ : CascadeMux
    port map (
            O => \N__41385\,
            I => \n1920_cascade_\
        );

    \I__8389\ : InMux
    port map (
            O => \N__41382\,
            I => \N__41379\
        );

    \I__8388\ : LocalMux
    port map (
            O => \N__41379\,
            I => \N__41375\
        );

    \I__8387\ : InMux
    port map (
            O => \N__41378\,
            I => \N__41371\
        );

    \I__8386\ : Span4Mux_v
    port map (
            O => \N__41375\,
            I => \N__41363\
        );

    \I__8385\ : InMux
    port map (
            O => \N__41374\,
            I => \N__41360\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__41371\,
            I => \N__41353\
        );

    \I__8383\ : InMux
    port map (
            O => \N__41370\,
            I => \N__41350\
        );

    \I__8382\ : CascadeMux
    port map (
            O => \N__41369\,
            I => \N__41347\
        );

    \I__8381\ : CascadeMux
    port map (
            O => \N__41368\,
            I => \N__41344\
        );

    \I__8380\ : CascadeMux
    port map (
            O => \N__41367\,
            I => \N__41337\
        );

    \I__8379\ : CascadeMux
    port map (
            O => \N__41366\,
            I => \N__41334\
        );

    \I__8378\ : Span4Mux_v
    port map (
            O => \N__41363\,
            I => \N__41327\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__41360\,
            I => \N__41327\
        );

    \I__8376\ : InMux
    port map (
            O => \N__41359\,
            I => \N__41324\
        );

    \I__8375\ : InMux
    port map (
            O => \N__41358\,
            I => \N__41317\
        );

    \I__8374\ : InMux
    port map (
            O => \N__41357\,
            I => \N__41317\
        );

    \I__8373\ : InMux
    port map (
            O => \N__41356\,
            I => \N__41317\
        );

    \I__8372\ : Span4Mux_h
    port map (
            O => \N__41353\,
            I => \N__41314\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__41350\,
            I => \N__41311\
        );

    \I__8370\ : InMux
    port map (
            O => \N__41347\,
            I => \N__41298\
        );

    \I__8369\ : InMux
    port map (
            O => \N__41344\,
            I => \N__41298\
        );

    \I__8368\ : InMux
    port map (
            O => \N__41343\,
            I => \N__41298\
        );

    \I__8367\ : InMux
    port map (
            O => \N__41342\,
            I => \N__41298\
        );

    \I__8366\ : InMux
    port map (
            O => \N__41341\,
            I => \N__41298\
        );

    \I__8365\ : InMux
    port map (
            O => \N__41340\,
            I => \N__41298\
        );

    \I__8364\ : InMux
    port map (
            O => \N__41337\,
            I => \N__41289\
        );

    \I__8363\ : InMux
    port map (
            O => \N__41334\,
            I => \N__41289\
        );

    \I__8362\ : InMux
    port map (
            O => \N__41333\,
            I => \N__41289\
        );

    \I__8361\ : InMux
    port map (
            O => \N__41332\,
            I => \N__41289\
        );

    \I__8360\ : Odrv4
    port map (
            O => \N__41327\,
            I => n1950
        );

    \I__8359\ : LocalMux
    port map (
            O => \N__41324\,
            I => n1950
        );

    \I__8358\ : LocalMux
    port map (
            O => \N__41317\,
            I => n1950
        );

    \I__8357\ : Odrv4
    port map (
            O => \N__41314\,
            I => n1950
        );

    \I__8356\ : Odrv4
    port map (
            O => \N__41311\,
            I => n1950
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__41298\,
            I => n1950
        );

    \I__8354\ : LocalMux
    port map (
            O => \N__41289\,
            I => n1950
        );

    \I__8353\ : CascadeMux
    port map (
            O => \N__41274\,
            I => \N__41269\
        );

    \I__8352\ : CascadeMux
    port map (
            O => \N__41273\,
            I => \N__41266\
        );

    \I__8351\ : CascadeMux
    port map (
            O => \N__41272\,
            I => \N__41263\
        );

    \I__8350\ : InMux
    port map (
            O => \N__41269\,
            I => \N__41260\
        );

    \I__8349\ : InMux
    port map (
            O => \N__41266\,
            I => \N__41257\
        );

    \I__8348\ : InMux
    port map (
            O => \N__41263\,
            I => \N__41254\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__41260\,
            I => \N__41251\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__41257\,
            I => \N__41248\
        );

    \I__8345\ : LocalMux
    port map (
            O => \N__41254\,
            I => \N__41245\
        );

    \I__8344\ : Span4Mux_v
    port map (
            O => \N__41251\,
            I => \N__41240\
        );

    \I__8343\ : Span4Mux_h
    port map (
            O => \N__41248\,
            I => \N__41240\
        );

    \I__8342\ : Span4Mux_h
    port map (
            O => \N__41245\,
            I => \N__41237\
        );

    \I__8341\ : Span4Mux_h
    port map (
            O => \N__41240\,
            I => \N__41234\
        );

    \I__8340\ : Odrv4
    port map (
            O => \N__41237\,
            I => n2019
        );

    \I__8339\ : Odrv4
    port map (
            O => \N__41234\,
            I => n2019
        );

    \I__8338\ : InMux
    port map (
            O => \N__41229\,
            I => \N__41224\
        );

    \I__8337\ : CascadeMux
    port map (
            O => \N__41228\,
            I => \N__41221\
        );

    \I__8336\ : InMux
    port map (
            O => \N__41227\,
            I => \N__41218\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__41224\,
            I => \N__41215\
        );

    \I__8334\ : InMux
    port map (
            O => \N__41221\,
            I => \N__41212\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__41218\,
            I => \N__41209\
        );

    \I__8332\ : Span4Mux_h
    port map (
            O => \N__41215\,
            I => \N__41206\
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__41212\,
            I => \N__41203\
        );

    \I__8330\ : Span4Mux_h
    port map (
            O => \N__41209\,
            I => \N__41200\
        );

    \I__8329\ : Odrv4
    port map (
            O => \N__41206\,
            I => n1819
        );

    \I__8328\ : Odrv4
    port map (
            O => \N__41203\,
            I => n1819
        );

    \I__8327\ : Odrv4
    port map (
            O => \N__41200\,
            I => n1819
        );

    \I__8326\ : CascadeMux
    port map (
            O => \N__41193\,
            I => \N__41190\
        );

    \I__8325\ : InMux
    port map (
            O => \N__41190\,
            I => \N__41187\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__41187\,
            I => \N__41184\
        );

    \I__8323\ : Odrv4
    port map (
            O => \N__41184\,
            I => n1889
        );

    \I__8322\ : InMux
    port map (
            O => \N__41181\,
            I => n12617
        );

    \I__8321\ : InMux
    port map (
            O => \N__41178\,
            I => n12618
        );

    \I__8320\ : CascadeMux
    port map (
            O => \N__41175\,
            I => \N__41172\
        );

    \I__8319\ : InMux
    port map (
            O => \N__41172\,
            I => \N__41169\
        );

    \I__8318\ : LocalMux
    port map (
            O => \N__41169\,
            I => \N__41166\
        );

    \I__8317\ : Odrv4
    port map (
            O => \N__41166\,
            I => n1887
        );

    \I__8316\ : InMux
    port map (
            O => \N__41163\,
            I => n12619
        );

    \I__8315\ : CascadeMux
    port map (
            O => \N__41160\,
            I => \N__41157\
        );

    \I__8314\ : InMux
    port map (
            O => \N__41157\,
            I => \N__41154\
        );

    \I__8313\ : LocalMux
    port map (
            O => \N__41154\,
            I => \N__41151\
        );

    \I__8312\ : Odrv4
    port map (
            O => \N__41151\,
            I => n1886
        );

    \I__8311\ : InMux
    port map (
            O => \N__41148\,
            I => n12620
        );

    \I__8310\ : InMux
    port map (
            O => \N__41145\,
            I => \bfn_11_19_0_\
        );

    \I__8309\ : CascadeMux
    port map (
            O => \N__41142\,
            I => \N__41139\
        );

    \I__8308\ : InMux
    port map (
            O => \N__41139\,
            I => \N__41136\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__41136\,
            I => n1892
        );

    \I__8306\ : CascadeMux
    port map (
            O => \N__41133\,
            I => \N__41129\
        );

    \I__8305\ : CascadeMux
    port map (
            O => \N__41132\,
            I => \N__41126\
        );

    \I__8304\ : InMux
    port map (
            O => \N__41129\,
            I => \N__41123\
        );

    \I__8303\ : InMux
    port map (
            O => \N__41126\,
            I => \N__41120\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__41123\,
            I => \N__41117\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__41120\,
            I => \N__41114\
        );

    \I__8300\ : Span4Mux_h
    port map (
            O => \N__41117\,
            I => \N__41111\
        );

    \I__8299\ : Odrv12
    port map (
            O => \N__41114\,
            I => n1924
        );

    \I__8298\ : Odrv4
    port map (
            O => \N__41111\,
            I => n1924
        );

    \I__8297\ : CascadeMux
    port map (
            O => \N__41106\,
            I => \n1924_cascade_\
        );

    \I__8296\ : InMux
    port map (
            O => \N__41103\,
            I => \N__41100\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__41100\,
            I => \N__41097\
        );

    \I__8294\ : Span4Mux_h
    port map (
            O => \N__41097\,
            I => \N__41094\
        );

    \I__8293\ : Odrv4
    port map (
            O => \N__41094\,
            I => n14438
        );

    \I__8292\ : InMux
    port map (
            O => \N__41091\,
            I => \N__41088\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__41088\,
            I => \N__41084\
        );

    \I__8290\ : CascadeMux
    port map (
            O => \N__41087\,
            I => \N__41081\
        );

    \I__8289\ : Span4Mux_h
    port map (
            O => \N__41084\,
            I => \N__41078\
        );

    \I__8288\ : InMux
    port map (
            O => \N__41081\,
            I => \N__41075\
        );

    \I__8287\ : Odrv4
    port map (
            O => \N__41078\,
            I => n1822
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__41075\,
            I => n1822
        );

    \I__8285\ : CascadeMux
    port map (
            O => \N__41070\,
            I => \n1822_cascade_\
        );

    \I__8284\ : InMux
    port map (
            O => \N__41067\,
            I => \N__41064\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__41064\,
            I => \N__41061\
        );

    \I__8282\ : Odrv4
    port map (
            O => \N__41061\,
            I => n14534
        );

    \I__8281\ : InMux
    port map (
            O => \N__41058\,
            I => n12608
        );

    \I__8280\ : InMux
    port map (
            O => \N__41055\,
            I => \N__41052\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__41052\,
            I => n1897
        );

    \I__8278\ : InMux
    port map (
            O => \N__41049\,
            I => n12609
        );

    \I__8277\ : InMux
    port map (
            O => \N__41046\,
            I => \N__41043\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__41043\,
            I => n1896
        );

    \I__8275\ : InMux
    port map (
            O => \N__41040\,
            I => n12610
        );

    \I__8274\ : InMux
    port map (
            O => \N__41037\,
            I => n12611
        );

    \I__8273\ : InMux
    port map (
            O => \N__41034\,
            I => n12612
        );

    \I__8272\ : InMux
    port map (
            O => \N__41031\,
            I => \N__41028\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__41028\,
            I => n1893
        );

    \I__8270\ : InMux
    port map (
            O => \N__41025\,
            I => \bfn_11_18_0_\
        );

    \I__8269\ : InMux
    port map (
            O => \N__41022\,
            I => n12614
        );

    \I__8268\ : CascadeMux
    port map (
            O => \N__41019\,
            I => \N__41016\
        );

    \I__8267\ : InMux
    port map (
            O => \N__41016\,
            I => \N__41013\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__41013\,
            I => n1891
        );

    \I__8265\ : InMux
    port map (
            O => \N__41010\,
            I => n12615
        );

    \I__8264\ : InMux
    port map (
            O => \N__41007\,
            I => \N__41004\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__41004\,
            I => \N__41001\
        );

    \I__8262\ : Span4Mux_v
    port map (
            O => \N__41001\,
            I => \N__40998\
        );

    \I__8261\ : Odrv4
    port map (
            O => \N__40998\,
            I => n1890
        );

    \I__8260\ : InMux
    port map (
            O => \N__40995\,
            I => n12616
        );

    \I__8259\ : InMux
    port map (
            O => \N__40992\,
            I => \N__40985\
        );

    \I__8258\ : InMux
    port map (
            O => \N__40991\,
            I => \N__40985\
        );

    \I__8257\ : InMux
    port map (
            O => \N__40990\,
            I => \N__40982\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__40985\,
            I => blink_counter_24
        );

    \I__8255\ : LocalMux
    port map (
            O => \N__40982\,
            I => blink_counter_24
        );

    \I__8254\ : InMux
    port map (
            O => \N__40977\,
            I => \bfn_10_32_0_\
        );

    \I__8253\ : InMux
    port map (
            O => \N__40974\,
            I => n13094
        );

    \I__8252\ : InMux
    port map (
            O => \N__40971\,
            I => \N__40967\
        );

    \I__8251\ : InMux
    port map (
            O => \N__40970\,
            I => \N__40964\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__40967\,
            I => blink_counter_25
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__40964\,
            I => blink_counter_25
        );

    \I__8248\ : CascadeMux
    port map (
            O => \N__40959\,
            I => \n1833_cascade_\
        );

    \I__8247\ : InMux
    port map (
            O => \N__40956\,
            I => \N__40953\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__40953\,
            I => n11989
        );

    \I__8245\ : InMux
    port map (
            O => \N__40950\,
            I => \N__40945\
        );

    \I__8244\ : InMux
    port map (
            O => \N__40949\,
            I => \N__40942\
        );

    \I__8243\ : InMux
    port map (
            O => \N__40948\,
            I => \N__40939\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__40945\,
            I => \N__40934\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__40942\,
            I => \N__40934\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__40939\,
            I => \N__40931\
        );

    \I__8239\ : Span4Mux_h
    port map (
            O => \N__40934\,
            I => \N__40928\
        );

    \I__8238\ : Span4Mux_h
    port map (
            O => \N__40931\,
            I => \N__40925\
        );

    \I__8237\ : Odrv4
    port map (
            O => \N__40928\,
            I => n304
        );

    \I__8236\ : Odrv4
    port map (
            O => \N__40925\,
            I => n304
        );

    \I__8235\ : InMux
    port map (
            O => \N__40920\,
            I => \N__40917\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__40917\,
            I => n1901
        );

    \I__8233\ : InMux
    port map (
            O => \N__40914\,
            I => \bfn_11_17_0_\
        );

    \I__8232\ : InMux
    port map (
            O => \N__40911\,
            I => \N__40907\
        );

    \I__8231\ : CascadeMux
    port map (
            O => \N__40910\,
            I => \N__40904\
        );

    \I__8230\ : LocalMux
    port map (
            O => \N__40907\,
            I => \N__40901\
        );

    \I__8229\ : InMux
    port map (
            O => \N__40904\,
            I => \N__40898\
        );

    \I__8228\ : Odrv4
    port map (
            O => \N__40901\,
            I => n1833
        );

    \I__8227\ : LocalMux
    port map (
            O => \N__40898\,
            I => n1833
        );

    \I__8226\ : InMux
    port map (
            O => \N__40893\,
            I => \N__40890\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__40890\,
            I => n1900
        );

    \I__8224\ : InMux
    port map (
            O => \N__40887\,
            I => n12606
        );

    \I__8223\ : CascadeMux
    port map (
            O => \N__40884\,
            I => \N__40880\
        );

    \I__8222\ : InMux
    port map (
            O => \N__40883\,
            I => \N__40876\
        );

    \I__8221\ : InMux
    port map (
            O => \N__40880\,
            I => \N__40873\
        );

    \I__8220\ : InMux
    port map (
            O => \N__40879\,
            I => \N__40870\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__40876\,
            I => n1832
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__40873\,
            I => n1832
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__40870\,
            I => n1832
        );

    \I__8216\ : CascadeMux
    port map (
            O => \N__40863\,
            I => \N__40860\
        );

    \I__8215\ : InMux
    port map (
            O => \N__40860\,
            I => \N__40857\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__40857\,
            I => n1899
        );

    \I__8213\ : InMux
    port map (
            O => \N__40854\,
            I => n12607
        );

    \I__8212\ : CascadeMux
    port map (
            O => \N__40851\,
            I => \N__40848\
        );

    \I__8211\ : InMux
    port map (
            O => \N__40848\,
            I => \N__40844\
        );

    \I__8210\ : InMux
    port map (
            O => \N__40847\,
            I => \N__40841\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__40844\,
            I => n1831
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__40841\,
            I => n1831
        );

    \I__8207\ : InMux
    port map (
            O => \N__40836\,
            I => \N__40833\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__40833\,
            I => n1898
        );

    \I__8205\ : InMux
    port map (
            O => \N__40830\,
            I => \N__40827\
        );

    \I__8204\ : LocalMux
    port map (
            O => \N__40827\,
            I => n10_adj_687
        );

    \I__8203\ : InMux
    port map (
            O => \N__40824\,
            I => \bfn_10_31_0_\
        );

    \I__8202\ : InMux
    port map (
            O => \N__40821\,
            I => \N__40818\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__40818\,
            I => n9_adj_686
        );

    \I__8200\ : InMux
    port map (
            O => \N__40815\,
            I => n13086
        );

    \I__8199\ : InMux
    port map (
            O => \N__40812\,
            I => \N__40809\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__40809\,
            I => n8_adj_685
        );

    \I__8197\ : InMux
    port map (
            O => \N__40806\,
            I => n13087
        );

    \I__8196\ : InMux
    port map (
            O => \N__40803\,
            I => \N__40800\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__40800\,
            I => n7_adj_684
        );

    \I__8194\ : InMux
    port map (
            O => \N__40797\,
            I => n13088
        );

    \I__8193\ : InMux
    port map (
            O => \N__40794\,
            I => \N__40791\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__40791\,
            I => n6_adj_683
        );

    \I__8191\ : InMux
    port map (
            O => \N__40788\,
            I => n13089
        );

    \I__8190\ : CascadeMux
    port map (
            O => \N__40785\,
            I => \N__40781\
        );

    \I__8189\ : InMux
    port map (
            O => \N__40784\,
            I => \N__40775\
        );

    \I__8188\ : InMux
    port map (
            O => \N__40781\,
            I => \N__40775\
        );

    \I__8187\ : InMux
    port map (
            O => \N__40780\,
            I => \N__40772\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__40775\,
            I => blink_counter_21
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__40772\,
            I => blink_counter_21
        );

    \I__8184\ : InMux
    port map (
            O => \N__40767\,
            I => n13090
        );

    \I__8183\ : InMux
    port map (
            O => \N__40764\,
            I => \N__40757\
        );

    \I__8182\ : InMux
    port map (
            O => \N__40763\,
            I => \N__40757\
        );

    \I__8181\ : InMux
    port map (
            O => \N__40762\,
            I => \N__40754\
        );

    \I__8180\ : LocalMux
    port map (
            O => \N__40757\,
            I => blink_counter_22
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__40754\,
            I => blink_counter_22
        );

    \I__8178\ : InMux
    port map (
            O => \N__40749\,
            I => n13091
        );

    \I__8177\ : CascadeMux
    port map (
            O => \N__40746\,
            I => \N__40743\
        );

    \I__8176\ : InMux
    port map (
            O => \N__40743\,
            I => \N__40736\
        );

    \I__8175\ : InMux
    port map (
            O => \N__40742\,
            I => \N__40736\
        );

    \I__8174\ : InMux
    port map (
            O => \N__40741\,
            I => \N__40733\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__40736\,
            I => blink_counter_23
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__40733\,
            I => blink_counter_23
        );

    \I__8171\ : InMux
    port map (
            O => \N__40728\,
            I => n13092
        );

    \I__8170\ : InMux
    port map (
            O => \N__40725\,
            I => \N__40722\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__40722\,
            I => n19_adj_696
        );

    \I__8168\ : InMux
    port map (
            O => \N__40719\,
            I => n13076
        );

    \I__8167\ : InMux
    port map (
            O => \N__40716\,
            I => \N__40713\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__40713\,
            I => n18_adj_695
        );

    \I__8165\ : InMux
    port map (
            O => \N__40710\,
            I => \bfn_10_30_0_\
        );

    \I__8164\ : InMux
    port map (
            O => \N__40707\,
            I => \N__40704\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__40704\,
            I => n17_adj_694
        );

    \I__8162\ : InMux
    port map (
            O => \N__40701\,
            I => n13078
        );

    \I__8161\ : InMux
    port map (
            O => \N__40698\,
            I => \N__40695\
        );

    \I__8160\ : LocalMux
    port map (
            O => \N__40695\,
            I => n16_adj_693
        );

    \I__8159\ : InMux
    port map (
            O => \N__40692\,
            I => n13079
        );

    \I__8158\ : InMux
    port map (
            O => \N__40689\,
            I => \N__40686\
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__40686\,
            I => n15_adj_692
        );

    \I__8156\ : InMux
    port map (
            O => \N__40683\,
            I => n13080
        );

    \I__8155\ : InMux
    port map (
            O => \N__40680\,
            I => \N__40677\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__40677\,
            I => n14_adj_691
        );

    \I__8153\ : InMux
    port map (
            O => \N__40674\,
            I => n13081
        );

    \I__8152\ : InMux
    port map (
            O => \N__40671\,
            I => \N__40668\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__40668\,
            I => n13_adj_690
        );

    \I__8150\ : InMux
    port map (
            O => \N__40665\,
            I => n13082
        );

    \I__8149\ : InMux
    port map (
            O => \N__40662\,
            I => \N__40659\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__40659\,
            I => n12_adj_689
        );

    \I__8147\ : InMux
    port map (
            O => \N__40656\,
            I => n13083
        );

    \I__8146\ : InMux
    port map (
            O => \N__40653\,
            I => \N__40650\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__40650\,
            I => n11_adj_688
        );

    \I__8144\ : InMux
    port map (
            O => \N__40647\,
            I => n13084
        );

    \I__8143\ : InMux
    port map (
            O => \N__40644\,
            I => \N__40641\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__40641\,
            I => n26_adj_703
        );

    \I__8141\ : InMux
    port map (
            O => \N__40638\,
            I => \bfn_10_29_0_\
        );

    \I__8140\ : InMux
    port map (
            O => \N__40635\,
            I => \N__40632\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__40632\,
            I => n25_adj_702
        );

    \I__8138\ : InMux
    port map (
            O => \N__40629\,
            I => n13070
        );

    \I__8137\ : InMux
    port map (
            O => \N__40626\,
            I => \N__40623\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__40623\,
            I => n24_adj_701
        );

    \I__8135\ : InMux
    port map (
            O => \N__40620\,
            I => n13071
        );

    \I__8134\ : InMux
    port map (
            O => \N__40617\,
            I => \N__40614\
        );

    \I__8133\ : LocalMux
    port map (
            O => \N__40614\,
            I => n23_adj_700
        );

    \I__8132\ : InMux
    port map (
            O => \N__40611\,
            I => n13072
        );

    \I__8131\ : InMux
    port map (
            O => \N__40608\,
            I => \N__40605\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__40605\,
            I => n22_adj_699
        );

    \I__8129\ : InMux
    port map (
            O => \N__40602\,
            I => n13073
        );

    \I__8128\ : InMux
    port map (
            O => \N__40599\,
            I => \N__40596\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__40596\,
            I => n21_adj_698
        );

    \I__8126\ : InMux
    port map (
            O => \N__40593\,
            I => n13074
        );

    \I__8125\ : InMux
    port map (
            O => \N__40590\,
            I => \N__40587\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__40587\,
            I => n20_adj_697
        );

    \I__8123\ : InMux
    port map (
            O => \N__40584\,
            I => n13075
        );

    \I__8122\ : InMux
    port map (
            O => \N__40581\,
            I => \N__40578\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__40578\,
            I => \N__40575\
        );

    \I__8120\ : Odrv12
    port map (
            O => \N__40575\,
            I => encoder0_position_scaled_21
        );

    \I__8119\ : InMux
    port map (
            O => \N__40572\,
            I => \N__40569\
        );

    \I__8118\ : LocalMux
    port map (
            O => \N__40569\,
            I => \N__40566\
        );

    \I__8117\ : Odrv4
    port map (
            O => \N__40566\,
            I => encoder0_position_scaled_19
        );

    \I__8116\ : InMux
    port map (
            O => \N__40563\,
            I => \N__40559\
        );

    \I__8115\ : InMux
    port map (
            O => \N__40562\,
            I => \N__40556\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__40559\,
            I => pwm_setpoint_4
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__40556\,
            I => pwm_setpoint_4
        );

    \I__8112\ : InMux
    port map (
            O => \N__40551\,
            I => \N__40548\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__40548\,
            I => \N__40545\
        );

    \I__8110\ : Odrv12
    port map (
            O => \N__40545\,
            I => encoder0_position_scaled_22
        );

    \I__8109\ : InMux
    port map (
            O => \N__40542\,
            I => \N__40538\
        );

    \I__8108\ : InMux
    port map (
            O => \N__40541\,
            I => \N__40535\
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__40538\,
            I => \N__40532\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__40535\,
            I => \quad_counter0.a_prev\
        );

    \I__8105\ : Odrv4
    port map (
            O => \N__40532\,
            I => \quad_counter0.a_prev\
        );

    \I__8104\ : CascadeMux
    port map (
            O => \N__40527\,
            I => \N__40509\
        );

    \I__8103\ : CascadeMux
    port map (
            O => \N__40526\,
            I => \N__40505\
        );

    \I__8102\ : CascadeMux
    port map (
            O => \N__40525\,
            I => \N__40501\
        );

    \I__8101\ : CascadeMux
    port map (
            O => \N__40524\,
            I => \N__40497\
        );

    \I__8100\ : CascadeMux
    port map (
            O => \N__40523\,
            I => \N__40493\
        );

    \I__8099\ : CascadeMux
    port map (
            O => \N__40522\,
            I => \N__40489\
        );

    \I__8098\ : CascadeMux
    port map (
            O => \N__40521\,
            I => \N__40485\
        );

    \I__8097\ : CascadeMux
    port map (
            O => \N__40520\,
            I => \N__40481\
        );

    \I__8096\ : CascadeMux
    port map (
            O => \N__40519\,
            I => \N__40477\
        );

    \I__8095\ : CascadeMux
    port map (
            O => \N__40518\,
            I => \N__40473\
        );

    \I__8094\ : CascadeMux
    port map (
            O => \N__40517\,
            I => \N__40469\
        );

    \I__8093\ : CascadeMux
    port map (
            O => \N__40516\,
            I => \N__40464\
        );

    \I__8092\ : CascadeMux
    port map (
            O => \N__40515\,
            I => \N__40460\
        );

    \I__8091\ : CascadeMux
    port map (
            O => \N__40514\,
            I => \N__40456\
        );

    \I__8090\ : InMux
    port map (
            O => \N__40513\,
            I => \N__40438\
        );

    \I__8089\ : InMux
    port map (
            O => \N__40512\,
            I => \N__40438\
        );

    \I__8088\ : InMux
    port map (
            O => \N__40509\,
            I => \N__40438\
        );

    \I__8087\ : InMux
    port map (
            O => \N__40508\,
            I => \N__40438\
        );

    \I__8086\ : InMux
    port map (
            O => \N__40505\,
            I => \N__40438\
        );

    \I__8085\ : InMux
    port map (
            O => \N__40504\,
            I => \N__40438\
        );

    \I__8084\ : InMux
    port map (
            O => \N__40501\,
            I => \N__40438\
        );

    \I__8083\ : InMux
    port map (
            O => \N__40500\,
            I => \N__40438\
        );

    \I__8082\ : InMux
    port map (
            O => \N__40497\,
            I => \N__40421\
        );

    \I__8081\ : InMux
    port map (
            O => \N__40496\,
            I => \N__40421\
        );

    \I__8080\ : InMux
    port map (
            O => \N__40493\,
            I => \N__40421\
        );

    \I__8079\ : InMux
    port map (
            O => \N__40492\,
            I => \N__40421\
        );

    \I__8078\ : InMux
    port map (
            O => \N__40489\,
            I => \N__40421\
        );

    \I__8077\ : InMux
    port map (
            O => \N__40488\,
            I => \N__40421\
        );

    \I__8076\ : InMux
    port map (
            O => \N__40485\,
            I => \N__40421\
        );

    \I__8075\ : InMux
    port map (
            O => \N__40484\,
            I => \N__40421\
        );

    \I__8074\ : InMux
    port map (
            O => \N__40481\,
            I => \N__40404\
        );

    \I__8073\ : InMux
    port map (
            O => \N__40480\,
            I => \N__40404\
        );

    \I__8072\ : InMux
    port map (
            O => \N__40477\,
            I => \N__40404\
        );

    \I__8071\ : InMux
    port map (
            O => \N__40476\,
            I => \N__40404\
        );

    \I__8070\ : InMux
    port map (
            O => \N__40473\,
            I => \N__40404\
        );

    \I__8069\ : InMux
    port map (
            O => \N__40472\,
            I => \N__40404\
        );

    \I__8068\ : InMux
    port map (
            O => \N__40469\,
            I => \N__40404\
        );

    \I__8067\ : InMux
    port map (
            O => \N__40468\,
            I => \N__40404\
        );

    \I__8066\ : InMux
    port map (
            O => \N__40467\,
            I => \N__40389\
        );

    \I__8065\ : InMux
    port map (
            O => \N__40464\,
            I => \N__40389\
        );

    \I__8064\ : InMux
    port map (
            O => \N__40463\,
            I => \N__40389\
        );

    \I__8063\ : InMux
    port map (
            O => \N__40460\,
            I => \N__40389\
        );

    \I__8062\ : InMux
    port map (
            O => \N__40459\,
            I => \N__40389\
        );

    \I__8061\ : InMux
    port map (
            O => \N__40456\,
            I => \N__40389\
        );

    \I__8060\ : InMux
    port map (
            O => \N__40455\,
            I => \N__40389\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__40438\,
            I => \N__40386\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__40421\,
            I => \N__40379\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__40404\,
            I => \N__40379\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__40389\,
            I => \N__40379\
        );

    \I__8055\ : Sp12to4
    port map (
            O => \N__40386\,
            I => \N__40374\
        );

    \I__8054\ : Span12Mux_v
    port map (
            O => \N__40379\,
            I => \N__40374\
        );

    \I__8053\ : Odrv12
    port map (
            O => \N__40374\,
            I => \quad_counter0.direction_N_536\
        );

    \I__8052\ : InMux
    port map (
            O => \N__40371\,
            I => \N__40368\
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__40368\,
            I => \N__40365\
        );

    \I__8050\ : Odrv4
    port map (
            O => \N__40365\,
            I => encoder0_position_scaled_1
        );

    \I__8049\ : InMux
    port map (
            O => \N__40362\,
            I => \N__40359\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__40359\,
            I => \quad_counter0.direction_N_540\
        );

    \I__8047\ : InMux
    port map (
            O => \N__40356\,
            I => \N__40353\
        );

    \I__8046\ : LocalMux
    port map (
            O => \N__40353\,
            I => \N__40350\
        );

    \I__8045\ : Odrv4
    port map (
            O => \N__40350\,
            I => encoder0_position_scaled_9
        );

    \I__8044\ : InMux
    port map (
            O => \N__40347\,
            I => \N__40344\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__40344\,
            I => \N__40341\
        );

    \I__8042\ : Span4Mux_h
    port map (
            O => \N__40341\,
            I => \N__40338\
        );

    \I__8041\ : Odrv4
    port map (
            O => \N__40338\,
            I => encoder0_position_scaled_20
        );

    \I__8040\ : InMux
    port map (
            O => \N__40335\,
            I => \N__40332\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__40332\,
            I => \N__40329\
        );

    \I__8038\ : Odrv12
    port map (
            O => \N__40329\,
            I => encoder0_position_scaled_11
        );

    \I__8037\ : CascadeMux
    port map (
            O => \N__40326\,
            I => \N__40323\
        );

    \I__8036\ : InMux
    port map (
            O => \N__40323\,
            I => \N__40320\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__40320\,
            I => n15_adj_633
        );

    \I__8034\ : CascadeMux
    port map (
            O => \N__40317\,
            I => \N__40314\
        );

    \I__8033\ : InMux
    port map (
            O => \N__40314\,
            I => \N__40311\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__40311\,
            I => n6_adj_624
        );

    \I__8031\ : CEMux
    port map (
            O => \N__40308\,
            I => \N__40305\
        );

    \I__8030\ : LocalMux
    port map (
            O => \N__40305\,
            I => \N__40299\
        );

    \I__8029\ : CEMux
    port map (
            O => \N__40304\,
            I => \N__40296\
        );

    \I__8028\ : CEMux
    port map (
            O => \N__40303\,
            I => \N__40293\
        );

    \I__8027\ : CEMux
    port map (
            O => \N__40302\,
            I => \N__40290\
        );

    \I__8026\ : Span4Mux_v
    port map (
            O => \N__40299\,
            I => \N__40287\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__40296\,
            I => \N__40284\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__40293\,
            I => \N__40281\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__40290\,
            I => \N__40278\
        );

    \I__8022\ : Span4Mux_v
    port map (
            O => \N__40287\,
            I => \N__40275\
        );

    \I__8021\ : Span12Mux_v
    port map (
            O => \N__40284\,
            I => \N__40272\
        );

    \I__8020\ : Span4Mux_v
    port map (
            O => \N__40281\,
            I => \N__40267\
        );

    \I__8019\ : Span4Mux_h
    port map (
            O => \N__40278\,
            I => \N__40267\
        );

    \I__8018\ : Odrv4
    port map (
            O => \N__40275\,
            I => \direction_N_537\
        );

    \I__8017\ : Odrv12
    port map (
            O => \N__40272\,
            I => \direction_N_537\
        );

    \I__8016\ : Odrv4
    port map (
            O => \N__40267\,
            I => \direction_N_537\
        );

    \I__8015\ : CascadeMux
    port map (
            O => \N__40260\,
            I => \direction_N_537_cascade_\
        );

    \I__8014\ : InMux
    port map (
            O => \N__40257\,
            I => \N__40254\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__40254\,
            I => n1302
        );

    \I__8012\ : CascadeMux
    port map (
            O => \N__40251\,
            I => \N__40248\
        );

    \I__8011\ : InMux
    port map (
            O => \N__40248\,
            I => \N__40245\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__40245\,
            I => n8_adj_626
        );

    \I__8009\ : CascadeMux
    port map (
            O => \N__40242\,
            I => \N__40239\
        );

    \I__8008\ : InMux
    port map (
            O => \N__40239\,
            I => \N__40236\
        );

    \I__8007\ : LocalMux
    port map (
            O => \N__40236\,
            I => n5_adj_623
        );

    \I__8006\ : CascadeMux
    port map (
            O => \N__40233\,
            I => \N__40217\
        );

    \I__8005\ : CascadeMux
    port map (
            O => \N__40232\,
            I => \N__40214\
        );

    \I__8004\ : CascadeMux
    port map (
            O => \N__40231\,
            I => \N__40211\
        );

    \I__8003\ : CascadeMux
    port map (
            O => \N__40230\,
            I => \N__40207\
        );

    \I__8002\ : CascadeMux
    port map (
            O => \N__40229\,
            I => \N__40203\
        );

    \I__8001\ : CascadeMux
    port map (
            O => \N__40228\,
            I => \N__40200\
        );

    \I__8000\ : CascadeMux
    port map (
            O => \N__40227\,
            I => \N__40197\
        );

    \I__7999\ : CascadeMux
    port map (
            O => \N__40226\,
            I => \N__40194\
        );

    \I__7998\ : CascadeMux
    port map (
            O => \N__40225\,
            I => \N__40191\
        );

    \I__7997\ : CascadeMux
    port map (
            O => \N__40224\,
            I => \N__40188\
        );

    \I__7996\ : CascadeMux
    port map (
            O => \N__40223\,
            I => \N__40185\
        );

    \I__7995\ : CascadeMux
    port map (
            O => \N__40222\,
            I => \N__40182\
        );

    \I__7994\ : CascadeMux
    port map (
            O => \N__40221\,
            I => \N__40179\
        );

    \I__7993\ : CascadeMux
    port map (
            O => \N__40220\,
            I => \N__40176\
        );

    \I__7992\ : InMux
    port map (
            O => \N__40217\,
            I => \N__40164\
        );

    \I__7991\ : InMux
    port map (
            O => \N__40214\,
            I => \N__40164\
        );

    \I__7990\ : InMux
    port map (
            O => \N__40211\,
            I => \N__40151\
        );

    \I__7989\ : InMux
    port map (
            O => \N__40210\,
            I => \N__40151\
        );

    \I__7988\ : InMux
    port map (
            O => \N__40207\,
            I => \N__40151\
        );

    \I__7987\ : InMux
    port map (
            O => \N__40206\,
            I => \N__40151\
        );

    \I__7986\ : InMux
    port map (
            O => \N__40203\,
            I => \N__40151\
        );

    \I__7985\ : InMux
    port map (
            O => \N__40200\,
            I => \N__40151\
        );

    \I__7984\ : InMux
    port map (
            O => \N__40197\,
            I => \N__40142\
        );

    \I__7983\ : InMux
    port map (
            O => \N__40194\,
            I => \N__40142\
        );

    \I__7982\ : InMux
    port map (
            O => \N__40191\,
            I => \N__40142\
        );

    \I__7981\ : InMux
    port map (
            O => \N__40188\,
            I => \N__40142\
        );

    \I__7980\ : InMux
    port map (
            O => \N__40185\,
            I => \N__40133\
        );

    \I__7979\ : InMux
    port map (
            O => \N__40182\,
            I => \N__40133\
        );

    \I__7978\ : InMux
    port map (
            O => \N__40179\,
            I => \N__40133\
        );

    \I__7977\ : InMux
    port map (
            O => \N__40176\,
            I => \N__40133\
        );

    \I__7976\ : CascadeMux
    port map (
            O => \N__40175\,
            I => \N__40130\
        );

    \I__7975\ : CascadeMux
    port map (
            O => \N__40174\,
            I => \N__40127\
        );

    \I__7974\ : CascadeMux
    port map (
            O => \N__40173\,
            I => \N__40124\
        );

    \I__7973\ : CascadeMux
    port map (
            O => \N__40172\,
            I => \N__40121\
        );

    \I__7972\ : CascadeMux
    port map (
            O => \N__40171\,
            I => \N__40118\
        );

    \I__7971\ : CascadeMux
    port map (
            O => \N__40170\,
            I => \N__40115\
        );

    \I__7970\ : CascadeMux
    port map (
            O => \N__40169\,
            I => \N__40112\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__40164\,
            I => \N__40102\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__40151\,
            I => \N__40102\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__40142\,
            I => \N__40102\
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__40133\,
            I => \N__40102\
        );

    \I__7965\ : InMux
    port map (
            O => \N__40130\,
            I => \N__40095\
        );

    \I__7964\ : InMux
    port map (
            O => \N__40127\,
            I => \N__40095\
        );

    \I__7963\ : InMux
    port map (
            O => \N__40124\,
            I => \N__40095\
        );

    \I__7962\ : InMux
    port map (
            O => \N__40121\,
            I => \N__40084\
        );

    \I__7961\ : InMux
    port map (
            O => \N__40118\,
            I => \N__40084\
        );

    \I__7960\ : InMux
    port map (
            O => \N__40115\,
            I => \N__40084\
        );

    \I__7959\ : InMux
    port map (
            O => \N__40112\,
            I => \N__40084\
        );

    \I__7958\ : InMux
    port map (
            O => \N__40111\,
            I => \N__40084\
        );

    \I__7957\ : Span4Mux_v
    port map (
            O => \N__40102\,
            I => \N__40080\
        );

    \I__7956\ : LocalMux
    port map (
            O => \N__40095\,
            I => \N__40075\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__40084\,
            I => \N__40075\
        );

    \I__7954\ : InMux
    port map (
            O => \N__40083\,
            I => \N__40072\
        );

    \I__7953\ : Odrv4
    port map (
            O => \N__40080\,
            I => n2_adj_620
        );

    \I__7952\ : Odrv12
    port map (
            O => \N__40075\,
            I => n2_adj_620
        );

    \I__7951\ : LocalMux
    port map (
            O => \N__40072\,
            I => n2_adj_620
        );

    \I__7950\ : CascadeMux
    port map (
            O => \N__40065\,
            I => \N__40062\
        );

    \I__7949\ : InMux
    port map (
            O => \N__40062\,
            I => \N__40059\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__40059\,
            I => n9_adj_627
        );

    \I__7947\ : InMux
    port map (
            O => \N__40056\,
            I => \N__40053\
        );

    \I__7946\ : LocalMux
    port map (
            O => \N__40053\,
            I => \N__40050\
        );

    \I__7945\ : Odrv4
    port map (
            O => \N__40050\,
            I => encoder0_position_scaled_5
        );

    \I__7944\ : CascadeMux
    port map (
            O => \N__40047\,
            I => \N__40044\
        );

    \I__7943\ : InMux
    port map (
            O => \N__40044\,
            I => \N__40041\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__40041\,
            I => n38
        );

    \I__7941\ : CascadeMux
    port map (
            O => \N__40038\,
            I => \N__40035\
        );

    \I__7940\ : InMux
    port map (
            O => \N__40035\,
            I => \N__40032\
        );

    \I__7939\ : LocalMux
    port map (
            O => \N__40032\,
            I => n402
        );

    \I__7938\ : CascadeMux
    port map (
            O => \N__40029\,
            I => \N__40026\
        );

    \I__7937\ : InMux
    port map (
            O => \N__40026\,
            I => \N__40023\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__40023\,
            I => n39
        );

    \I__7935\ : InMux
    port map (
            O => \N__40020\,
            I => \N__40017\
        );

    \I__7934\ : LocalMux
    port map (
            O => \N__40017\,
            I => n2562
        );

    \I__7933\ : CEMux
    port map (
            O => \N__40014\,
            I => \N__40011\
        );

    \I__7932\ : LocalMux
    port map (
            O => \N__40011\,
            I => \N__40008\
        );

    \I__7931\ : Span4Mux_h
    port map (
            O => \N__40008\,
            I => \N__40005\
        );

    \I__7930\ : Odrv4
    port map (
            O => \N__40005\,
            I => n5187
        );

    \I__7929\ : InMux
    port map (
            O => \N__40002\,
            I => \N__39997\
        );

    \I__7928\ : InMux
    port map (
            O => \N__40001\,
            I => \N__39994\
        );

    \I__7927\ : InMux
    port map (
            O => \N__40000\,
            I => \N__39991\
        );

    \I__7926\ : LocalMux
    port map (
            O => \N__39997\,
            I => \N__39988\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__39994\,
            I => encoder0_position_11
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__39991\,
            I => encoder0_position_11
        );

    \I__7923\ : Odrv12
    port map (
            O => \N__39988\,
            I => encoder0_position_11
        );

    \I__7922\ : CascadeMux
    port map (
            O => \N__39981\,
            I => \N__39978\
        );

    \I__7921\ : InMux
    port map (
            O => \N__39978\,
            I => \N__39975\
        );

    \I__7920\ : LocalMux
    port map (
            O => \N__39975\,
            I => n22_adj_640
        );

    \I__7919\ : InMux
    port map (
            O => \N__39972\,
            I => \N__39967\
        );

    \I__7918\ : InMux
    port map (
            O => \N__39971\,
            I => \N__39964\
        );

    \I__7917\ : CascadeMux
    port map (
            O => \N__39970\,
            I => \N__39961\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__39967\,
            I => \N__39958\
        );

    \I__7915\ : LocalMux
    port map (
            O => \N__39964\,
            I => \N__39955\
        );

    \I__7914\ : InMux
    port map (
            O => \N__39961\,
            I => \N__39952\
        );

    \I__7913\ : Span4Mux_h
    port map (
            O => \N__39958\,
            I => \N__39949\
        );

    \I__7912\ : Span4Mux_v
    port map (
            O => \N__39955\,
            I => \N__39946\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__39952\,
            I => encoder0_position_12
        );

    \I__7910\ : Odrv4
    port map (
            O => \N__39949\,
            I => encoder0_position_12
        );

    \I__7909\ : Odrv4
    port map (
            O => \N__39946\,
            I => encoder0_position_12
        );

    \I__7908\ : CascadeMux
    port map (
            O => \N__39939\,
            I => \N__39936\
        );

    \I__7907\ : InMux
    port map (
            O => \N__39936\,
            I => \N__39933\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__39933\,
            I => n21_adj_639
        );

    \I__7905\ : InMux
    port map (
            O => \N__39930\,
            I => \N__39925\
        );

    \I__7904\ : InMux
    port map (
            O => \N__39929\,
            I => \N__39922\
        );

    \I__7903\ : InMux
    port map (
            O => \N__39928\,
            I => \N__39919\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__39925\,
            I => \N__39916\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__39922\,
            I => encoder0_position_13
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__39919\,
            I => encoder0_position_13
        );

    \I__7899\ : Odrv12
    port map (
            O => \N__39916\,
            I => encoder0_position_13
        );

    \I__7898\ : CascadeMux
    port map (
            O => \N__39909\,
            I => \N__39906\
        );

    \I__7897\ : InMux
    port map (
            O => \N__39906\,
            I => \N__39903\
        );

    \I__7896\ : LocalMux
    port map (
            O => \N__39903\,
            I => n20_adj_638
        );

    \I__7895\ : InMux
    port map (
            O => \N__39900\,
            I => n12496
        );

    \I__7894\ : InMux
    port map (
            O => \N__39897\,
            I => n12497
        );

    \I__7893\ : InMux
    port map (
            O => \N__39894\,
            I => n12498
        );

    \I__7892\ : InMux
    port map (
            O => \N__39891\,
            I => n12499
        );

    \I__7891\ : InMux
    port map (
            O => \N__39888\,
            I => n12500
        );

    \I__7890\ : InMux
    port map (
            O => \N__39885\,
            I => \N__39882\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__39882\,
            I => n2563
        );

    \I__7888\ : InMux
    port map (
            O => \N__39879\,
            I => \N__39876\
        );

    \I__7887\ : LocalMux
    port map (
            O => \N__39876\,
            I => n13656
        );

    \I__7886\ : CascadeMux
    port map (
            O => \N__39873\,
            I => \N__39870\
        );

    \I__7885\ : InMux
    port map (
            O => \N__39870\,
            I => \N__39867\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__39867\,
            I => n403
        );

    \I__7883\ : CascadeMux
    port map (
            O => \N__39864\,
            I => \N__39861\
        );

    \I__7882\ : InMux
    port map (
            O => \N__39861\,
            I => \N__39858\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__39858\,
            I => n13_adj_631
        );

    \I__7880\ : InMux
    port map (
            O => \N__39855\,
            I => \bfn_10_21_0_\
        );

    \I__7879\ : InMux
    port map (
            O => \N__39852\,
            I => \quad_counter0.n13119\
        );

    \I__7878\ : InMux
    port map (
            O => \N__39849\,
            I => \quad_counter0.n13120\
        );

    \I__7877\ : InMux
    port map (
            O => \N__39846\,
            I => \quad_counter0.n13121\
        );

    \I__7876\ : InMux
    port map (
            O => \N__39843\,
            I => \quad_counter0.n13122\
        );

    \I__7875\ : InMux
    port map (
            O => \N__39840\,
            I => \quad_counter0.n13123\
        );

    \I__7874\ : InMux
    port map (
            O => \N__39837\,
            I => \quad_counter0.n13124\
        );

    \I__7873\ : InMux
    port map (
            O => \N__39834\,
            I => \quad_counter0.n13125\
        );

    \I__7872\ : InMux
    port map (
            O => \N__39831\,
            I => \bfn_10_22_0_\
        );

    \I__7871\ : InMux
    port map (
            O => \N__39828\,
            I => \N__39823\
        );

    \I__7870\ : InMux
    port map (
            O => \N__39827\,
            I => \N__39818\
        );

    \I__7869\ : InMux
    port map (
            O => \N__39826\,
            I => \N__39818\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__39823\,
            I => encoder0_position_15
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__39818\,
            I => encoder0_position_15
        );

    \I__7866\ : InMux
    port map (
            O => \N__39813\,
            I => \quad_counter0.n13109\
        );

    \I__7865\ : InMux
    port map (
            O => \N__39810\,
            I => \bfn_10_20_0_\
        );

    \I__7864\ : InMux
    port map (
            O => \N__39807\,
            I => \quad_counter0.n13111\
        );

    \I__7863\ : InMux
    port map (
            O => \N__39804\,
            I => \quad_counter0.n13112\
        );

    \I__7862\ : CascadeMux
    port map (
            O => \N__39801\,
            I => \N__39796\
        );

    \I__7861\ : InMux
    port map (
            O => \N__39800\,
            I => \N__39793\
        );

    \I__7860\ : InMux
    port map (
            O => \N__39799\,
            I => \N__39790\
        );

    \I__7859\ : InMux
    port map (
            O => \N__39796\,
            I => \N__39787\
        );

    \I__7858\ : LocalMux
    port map (
            O => \N__39793\,
            I => encoder0_position_19
        );

    \I__7857\ : LocalMux
    port map (
            O => \N__39790\,
            I => encoder0_position_19
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__39787\,
            I => encoder0_position_19
        );

    \I__7855\ : InMux
    port map (
            O => \N__39780\,
            I => \quad_counter0.n13113\
        );

    \I__7854\ : InMux
    port map (
            O => \N__39777\,
            I => \quad_counter0.n13114\
        );

    \I__7853\ : InMux
    port map (
            O => \N__39774\,
            I => \quad_counter0.n13115\
        );

    \I__7852\ : InMux
    port map (
            O => \N__39771\,
            I => \quad_counter0.n13116\
        );

    \I__7851\ : InMux
    port map (
            O => \N__39768\,
            I => \quad_counter0.n13117\
        );

    \I__7850\ : InMux
    port map (
            O => \N__39765\,
            I => \N__39761\
        );

    \I__7849\ : CascadeMux
    port map (
            O => \N__39764\,
            I => \N__39757\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__39761\,
            I => \N__39754\
        );

    \I__7847\ : InMux
    port map (
            O => \N__39760\,
            I => \N__39751\
        );

    \I__7846\ : InMux
    port map (
            O => \N__39757\,
            I => \N__39748\
        );

    \I__7845\ : Span4Mux_h
    port map (
            O => \N__39754\,
            I => \N__39743\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__39751\,
            I => \N__39743\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__39748\,
            I => encoder0_position_7
        );

    \I__7842\ : Odrv4
    port map (
            O => \N__39743\,
            I => encoder0_position_7
        );

    \I__7841\ : InMux
    port map (
            O => \N__39738\,
            I => \quad_counter0.n13101\
        );

    \I__7840\ : InMux
    port map (
            O => \N__39735\,
            I => \N__39732\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__39732\,
            I => \N__39728\
        );

    \I__7838\ : CascadeMux
    port map (
            O => \N__39731\,
            I => \N__39724\
        );

    \I__7837\ : Span4Mux_h
    port map (
            O => \N__39728\,
            I => \N__39721\
        );

    \I__7836\ : CascadeMux
    port map (
            O => \N__39727\,
            I => \N__39718\
        );

    \I__7835\ : InMux
    port map (
            O => \N__39724\,
            I => \N__39715\
        );

    \I__7834\ : Span4Mux_v
    port map (
            O => \N__39721\,
            I => \N__39712\
        );

    \I__7833\ : InMux
    port map (
            O => \N__39718\,
            I => \N__39709\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__39715\,
            I => encoder0_position_8
        );

    \I__7831\ : Odrv4
    port map (
            O => \N__39712\,
            I => encoder0_position_8
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__39709\,
            I => encoder0_position_8
        );

    \I__7829\ : InMux
    port map (
            O => \N__39702\,
            I => \bfn_10_19_0_\
        );

    \I__7828\ : InMux
    port map (
            O => \N__39699\,
            I => \N__39696\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__39696\,
            I => \N__39692\
        );

    \I__7826\ : InMux
    port map (
            O => \N__39695\,
            I => \N__39688\
        );

    \I__7825\ : Span4Mux_h
    port map (
            O => \N__39692\,
            I => \N__39685\
        );

    \I__7824\ : InMux
    port map (
            O => \N__39691\,
            I => \N__39682\
        );

    \I__7823\ : LocalMux
    port map (
            O => \N__39688\,
            I => encoder0_position_9
        );

    \I__7822\ : Odrv4
    port map (
            O => \N__39685\,
            I => encoder0_position_9
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__39682\,
            I => encoder0_position_9
        );

    \I__7820\ : InMux
    port map (
            O => \N__39675\,
            I => \quad_counter0.n13103\
        );

    \I__7819\ : CascadeMux
    port map (
            O => \N__39672\,
            I => \N__39668\
        );

    \I__7818\ : InMux
    port map (
            O => \N__39671\,
            I => \N__39665\
        );

    \I__7817\ : InMux
    port map (
            O => \N__39668\,
            I => \N__39661\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__39665\,
            I => \N__39658\
        );

    \I__7815\ : InMux
    port map (
            O => \N__39664\,
            I => \N__39655\
        );

    \I__7814\ : LocalMux
    port map (
            O => \N__39661\,
            I => encoder0_position_10
        );

    \I__7813\ : Odrv4
    port map (
            O => \N__39658\,
            I => encoder0_position_10
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__39655\,
            I => encoder0_position_10
        );

    \I__7811\ : InMux
    port map (
            O => \N__39648\,
            I => \quad_counter0.n13104\
        );

    \I__7810\ : InMux
    port map (
            O => \N__39645\,
            I => \quad_counter0.n13105\
        );

    \I__7809\ : InMux
    port map (
            O => \N__39642\,
            I => \quad_counter0.n13106\
        );

    \I__7808\ : InMux
    port map (
            O => \N__39639\,
            I => \quad_counter0.n13107\
        );

    \I__7807\ : CascadeMux
    port map (
            O => \N__39636\,
            I => \N__39633\
        );

    \I__7806\ : InMux
    port map (
            O => \N__39633\,
            I => \N__39628\
        );

    \I__7805\ : InMux
    port map (
            O => \N__39632\,
            I => \N__39625\
        );

    \I__7804\ : InMux
    port map (
            O => \N__39631\,
            I => \N__39622\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__39628\,
            I => encoder0_position_14
        );

    \I__7802\ : LocalMux
    port map (
            O => \N__39625\,
            I => encoder0_position_14
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__39622\,
            I => encoder0_position_14
        );

    \I__7800\ : InMux
    port map (
            O => \N__39615\,
            I => \quad_counter0.n13108\
        );

    \I__7799\ : InMux
    port map (
            O => \N__39612\,
            I => \N__39609\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__39609\,
            I => \N__39605\
        );

    \I__7797\ : CascadeMux
    port map (
            O => \N__39608\,
            I => \N__39602\
        );

    \I__7796\ : Span4Mux_h
    port map (
            O => \N__39605\,
            I => \N__39598\
        );

    \I__7795\ : InMux
    port map (
            O => \N__39602\,
            I => \N__39595\
        );

    \I__7794\ : InMux
    port map (
            O => \N__39601\,
            I => \N__39592\
        );

    \I__7793\ : Odrv4
    port map (
            O => \N__39598\,
            I => n1925
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__39595\,
            I => n1925
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__39592\,
            I => n1925
        );

    \I__7790\ : CascadeMux
    port map (
            O => \N__39585\,
            I => \n1928_cascade_\
        );

    \I__7789\ : InMux
    port map (
            O => \N__39582\,
            I => \N__39579\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__39579\,
            I => \N__39575\
        );

    \I__7787\ : CascadeMux
    port map (
            O => \N__39578\,
            I => \N__39572\
        );

    \I__7786\ : Span4Mux_h
    port map (
            O => \N__39575\,
            I => \N__39568\
        );

    \I__7785\ : InMux
    port map (
            O => \N__39572\,
            I => \N__39565\
        );

    \I__7784\ : InMux
    port map (
            O => \N__39571\,
            I => \N__39562\
        );

    \I__7783\ : Odrv4
    port map (
            O => \N__39568\,
            I => n1923
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__39565\,
            I => n1923
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__39562\,
            I => n1923
        );

    \I__7780\ : CascadeMux
    port map (
            O => \N__39555\,
            I => \N__39552\
        );

    \I__7779\ : InMux
    port map (
            O => \N__39552\,
            I => \N__39549\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__39549\,
            I => \N__39546\
        );

    \I__7777\ : Span4Mux_h
    port map (
            O => \N__39546\,
            I => \N__39543\
        );

    \I__7776\ : Odrv4
    port map (
            O => \N__39543\,
            I => n14440
        );

    \I__7775\ : InMux
    port map (
            O => \N__39540\,
            I => \N__39537\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__39537\,
            I => \N__39532\
        );

    \I__7773\ : InMux
    port map (
            O => \N__39536\,
            I => \N__39529\
        );

    \I__7772\ : CascadeMux
    port map (
            O => \N__39535\,
            I => \N__39526\
        );

    \I__7771\ : Span4Mux_v
    port map (
            O => \N__39532\,
            I => \N__39521\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__39529\,
            I => \N__39521\
        );

    \I__7769\ : InMux
    port map (
            O => \N__39526\,
            I => \N__39518\
        );

    \I__7768\ : Odrv4
    port map (
            O => \N__39521\,
            I => n1932
        );

    \I__7767\ : LocalMux
    port map (
            O => \N__39518\,
            I => n1932
        );

    \I__7766\ : InMux
    port map (
            O => \N__39513\,
            I => \N__39510\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__39510\,
            I => \N__39507\
        );

    \I__7764\ : Span4Mux_h
    port map (
            O => \N__39507\,
            I => \N__39502\
        );

    \I__7763\ : CascadeMux
    port map (
            O => \N__39506\,
            I => \N__39499\
        );

    \I__7762\ : InMux
    port map (
            O => \N__39505\,
            I => \N__39496\
        );

    \I__7761\ : Span4Mux_v
    port map (
            O => \N__39502\,
            I => \N__39493\
        );

    \I__7760\ : InMux
    port map (
            O => \N__39499\,
            I => \N__39490\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__39496\,
            I => encoder0_position_0
        );

    \I__7758\ : Odrv4
    port map (
            O => \N__39493\,
            I => encoder0_position_0
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__39490\,
            I => encoder0_position_0
        );

    \I__7756\ : InMux
    port map (
            O => \N__39483\,
            I => \bfn_10_18_0_\
        );

    \I__7755\ : InMux
    port map (
            O => \N__39480\,
            I => \quad_counter0.n13095\
        );

    \I__7754\ : InMux
    port map (
            O => \N__39477\,
            I => \N__39474\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__39474\,
            I => \N__39470\
        );

    \I__7752\ : InMux
    port map (
            O => \N__39473\,
            I => \N__39466\
        );

    \I__7751\ : Span4Mux_v
    port map (
            O => \N__39470\,
            I => \N__39463\
        );

    \I__7750\ : InMux
    port map (
            O => \N__39469\,
            I => \N__39460\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__39466\,
            I => encoder0_position_2
        );

    \I__7748\ : Odrv4
    port map (
            O => \N__39463\,
            I => encoder0_position_2
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__39460\,
            I => encoder0_position_2
        );

    \I__7746\ : InMux
    port map (
            O => \N__39453\,
            I => \quad_counter0.n13096\
        );

    \I__7745\ : InMux
    port map (
            O => \N__39450\,
            I => \quad_counter0.n13097\
        );

    \I__7744\ : InMux
    port map (
            O => \N__39447\,
            I => \N__39444\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__39444\,
            I => \N__39441\
        );

    \I__7742\ : Span4Mux_h
    port map (
            O => \N__39441\,
            I => \N__39436\
        );

    \I__7741\ : InMux
    port map (
            O => \N__39440\,
            I => \N__39433\
        );

    \I__7740\ : InMux
    port map (
            O => \N__39439\,
            I => \N__39430\
        );

    \I__7739\ : Span4Mux_v
    port map (
            O => \N__39436\,
            I => \N__39427\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__39433\,
            I => \N__39424\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__39430\,
            I => encoder0_position_4
        );

    \I__7736\ : Odrv4
    port map (
            O => \N__39427\,
            I => encoder0_position_4
        );

    \I__7735\ : Odrv4
    port map (
            O => \N__39424\,
            I => encoder0_position_4
        );

    \I__7734\ : InMux
    port map (
            O => \N__39417\,
            I => \quad_counter0.n13098\
        );

    \I__7733\ : InMux
    port map (
            O => \N__39414\,
            I => \N__39410\
        );

    \I__7732\ : CascadeMux
    port map (
            O => \N__39413\,
            I => \N__39407\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__39410\,
            I => \N__39404\
        );

    \I__7730\ : InMux
    port map (
            O => \N__39407\,
            I => \N__39400\
        );

    \I__7729\ : Span4Mux_v
    port map (
            O => \N__39404\,
            I => \N__39397\
        );

    \I__7728\ : InMux
    port map (
            O => \N__39403\,
            I => \N__39394\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__39400\,
            I => encoder0_position_5
        );

    \I__7726\ : Odrv4
    port map (
            O => \N__39397\,
            I => encoder0_position_5
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__39394\,
            I => encoder0_position_5
        );

    \I__7724\ : InMux
    port map (
            O => \N__39387\,
            I => \quad_counter0.n13099\
        );

    \I__7723\ : InMux
    port map (
            O => \N__39384\,
            I => \N__39381\
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__39381\,
            I => \N__39376\
        );

    \I__7721\ : InMux
    port map (
            O => \N__39380\,
            I => \N__39373\
        );

    \I__7720\ : InMux
    port map (
            O => \N__39379\,
            I => \N__39370\
        );

    \I__7719\ : Span4Mux_v
    port map (
            O => \N__39376\,
            I => \N__39367\
        );

    \I__7718\ : LocalMux
    port map (
            O => \N__39373\,
            I => \N__39364\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__39370\,
            I => encoder0_position_6
        );

    \I__7716\ : Odrv4
    port map (
            O => \N__39367\,
            I => encoder0_position_6
        );

    \I__7715\ : Odrv4
    port map (
            O => \N__39364\,
            I => encoder0_position_6
        );

    \I__7714\ : InMux
    port map (
            O => \N__39357\,
            I => \quad_counter0.n13100\
        );

    \I__7713\ : CascadeMux
    port map (
            O => \N__39354\,
            I => \N__39350\
        );

    \I__7712\ : InMux
    port map (
            O => \N__39353\,
            I => \N__39346\
        );

    \I__7711\ : InMux
    port map (
            O => \N__39350\,
            I => \N__39343\
        );

    \I__7710\ : CascadeMux
    port map (
            O => \N__39349\,
            I => \N__39340\
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__39346\,
            I => \N__39337\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__39343\,
            I => \N__39334\
        );

    \I__7707\ : InMux
    port map (
            O => \N__39340\,
            I => \N__39331\
        );

    \I__7706\ : Span4Mux_v
    port map (
            O => \N__39337\,
            I => \N__39328\
        );

    \I__7705\ : Odrv4
    port map (
            O => \N__39334\,
            I => n1931
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__39331\,
            I => n1931
        );

    \I__7703\ : Odrv4
    port map (
            O => \N__39328\,
            I => n1931
        );

    \I__7702\ : CascadeMux
    port map (
            O => \N__39321\,
            I => \N__39317\
        );

    \I__7701\ : InMux
    port map (
            O => \N__39320\,
            I => \N__39314\
        );

    \I__7700\ : InMux
    port map (
            O => \N__39317\,
            I => \N__39310\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__39314\,
            I => \N__39307\
        );

    \I__7698\ : CascadeMux
    port map (
            O => \N__39313\,
            I => \N__39304\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__39310\,
            I => \N__39301\
        );

    \I__7696\ : Span4Mux_h
    port map (
            O => \N__39307\,
            I => \N__39298\
        );

    \I__7695\ : InMux
    port map (
            O => \N__39304\,
            I => \N__39295\
        );

    \I__7694\ : Span4Mux_h
    port map (
            O => \N__39301\,
            I => \N__39292\
        );

    \I__7693\ : Odrv4
    port map (
            O => \N__39298\,
            I => n1933
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__39295\,
            I => n1933
        );

    \I__7691\ : Odrv4
    port map (
            O => \N__39292\,
            I => n1933
        );

    \I__7690\ : InMux
    port map (
            O => \N__39285\,
            I => \N__39282\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__39282\,
            I => \N__39277\
        );

    \I__7688\ : CascadeMux
    port map (
            O => \N__39281\,
            I => \N__39274\
        );

    \I__7687\ : InMux
    port map (
            O => \N__39280\,
            I => \N__39271\
        );

    \I__7686\ : Span4Mux_h
    port map (
            O => \N__39277\,
            I => \N__39268\
        );

    \I__7685\ : InMux
    port map (
            O => \N__39274\,
            I => \N__39265\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__39271\,
            I => \N__39262\
        );

    \I__7683\ : Odrv4
    port map (
            O => \N__39268\,
            I => n1929
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__39265\,
            I => n1929
        );

    \I__7681\ : Odrv4
    port map (
            O => \N__39262\,
            I => n1929
        );

    \I__7680\ : CascadeMux
    port map (
            O => \N__39255\,
            I => \n14524_cascade_\
        );

    \I__7679\ : CascadeMux
    port map (
            O => \N__39252\,
            I => \n14526_cascade_\
        );

    \I__7678\ : CascadeMux
    port map (
            O => \N__39249\,
            I => \n1851_cascade_\
        );

    \I__7677\ : InMux
    port map (
            O => \N__39246\,
            I => \N__39243\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__39243\,
            I => \N__39239\
        );

    \I__7675\ : CascadeMux
    port map (
            O => \N__39242\,
            I => \N__39236\
        );

    \I__7674\ : Span4Mux_v
    port map (
            O => \N__39239\,
            I => \N__39233\
        );

    \I__7673\ : InMux
    port map (
            O => \N__39236\,
            I => \N__39230\
        );

    \I__7672\ : Odrv4
    port map (
            O => \N__39233\,
            I => n1928
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__39230\,
            I => n1928
        );

    \I__7670\ : CascadeMux
    port map (
            O => \N__39225\,
            I => \N__39221\
        );

    \I__7669\ : CascadeMux
    port map (
            O => \N__39224\,
            I => \N__39218\
        );

    \I__7668\ : InMux
    port map (
            O => \N__39221\,
            I => \N__39215\
        );

    \I__7667\ : InMux
    port map (
            O => \N__39218\,
            I => \N__39211\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__39215\,
            I => \N__39208\
        );

    \I__7665\ : InMux
    port map (
            O => \N__39214\,
            I => \N__39205\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__39211\,
            I => dti_counter_1
        );

    \I__7663\ : Odrv4
    port map (
            O => \N__39208\,
            I => dti_counter_1
        );

    \I__7662\ : LocalMux
    port map (
            O => \N__39205\,
            I => dti_counter_1
        );

    \I__7661\ : InMux
    port map (
            O => \N__39198\,
            I => \N__39195\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__39195\,
            I => \N__39192\
        );

    \I__7659\ : Odrv4
    port map (
            O => \N__39192\,
            I => n15076
        );

    \I__7658\ : InMux
    port map (
            O => \N__39189\,
            I => \N__39176\
        );

    \I__7657\ : InMux
    port map (
            O => \N__39188\,
            I => \N__39176\
        );

    \I__7656\ : InMux
    port map (
            O => \N__39187\,
            I => \N__39165\
        );

    \I__7655\ : InMux
    port map (
            O => \N__39186\,
            I => \N__39165\
        );

    \I__7654\ : InMux
    port map (
            O => \N__39185\,
            I => \N__39165\
        );

    \I__7653\ : InMux
    port map (
            O => \N__39184\,
            I => \N__39165\
        );

    \I__7652\ : InMux
    port map (
            O => \N__39183\,
            I => \N__39165\
        );

    \I__7651\ : InMux
    port map (
            O => \N__39182\,
            I => \N__39160\
        );

    \I__7650\ : InMux
    port map (
            O => \N__39181\,
            I => \N__39160\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__39176\,
            I => \N__39157\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__39165\,
            I => commutation_state_prev_0
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__39160\,
            I => commutation_state_prev_0
        );

    \I__7646\ : Odrv12
    port map (
            O => \N__39157\,
            I => commutation_state_prev_0
        );

    \I__7645\ : InMux
    port map (
            O => \N__39150\,
            I => \N__39147\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__39147\,
            I => n14929
        );

    \I__7643\ : InMux
    port map (
            O => \N__39144\,
            I => \N__39141\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__39141\,
            I => n14928
        );

    \I__7641\ : IoInMux
    port map (
            O => \N__39138\,
            I => \N__39135\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__39135\,
            I => \N__39132\
        );

    \I__7639\ : IoSpan4Mux
    port map (
            O => \N__39132\,
            I => \N__39129\
        );

    \I__7638\ : Odrv4
    port map (
            O => \N__39129\,
            I => \LED_c\
        );

    \I__7637\ : CascadeMux
    port map (
            O => \N__39126\,
            I => \n1831_cascade_\
        );

    \I__7636\ : InMux
    port map (
            O => \N__39123\,
            I => \N__39119\
        );

    \I__7635\ : CascadeMux
    port map (
            O => \N__39122\,
            I => \N__39115\
        );

    \I__7634\ : LocalMux
    port map (
            O => \N__39119\,
            I => \N__39112\
        );

    \I__7633\ : CascadeMux
    port map (
            O => \N__39118\,
            I => \N__39109\
        );

    \I__7632\ : InMux
    port map (
            O => \N__39115\,
            I => \N__39106\
        );

    \I__7631\ : Span4Mux_h
    port map (
            O => \N__39112\,
            I => \N__39103\
        );

    \I__7630\ : InMux
    port map (
            O => \N__39109\,
            I => \N__39100\
        );

    \I__7629\ : LocalMux
    port map (
            O => \N__39106\,
            I => \N__39097\
        );

    \I__7628\ : Odrv4
    port map (
            O => \N__39103\,
            I => n1930
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__39100\,
            I => n1930
        );

    \I__7626\ : Odrv4
    port map (
            O => \N__39097\,
            I => n1930
        );

    \I__7625\ : InMux
    port map (
            O => \N__39090\,
            I => \N__39087\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__39087\,
            I => n15075
        );

    \I__7623\ : InMux
    port map (
            O => \N__39084\,
            I => \N__39081\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__39081\,
            I => n15071
        );

    \I__7621\ : CascadeMux
    port map (
            O => \N__39078\,
            I => \N__39074\
        );

    \I__7620\ : CascadeMux
    port map (
            O => \N__39077\,
            I => \N__39071\
        );

    \I__7619\ : InMux
    port map (
            O => \N__39074\,
            I => \N__39067\
        );

    \I__7618\ : InMux
    port map (
            O => \N__39071\,
            I => \N__39064\
        );

    \I__7617\ : InMux
    port map (
            O => \N__39070\,
            I => \N__39061\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__39067\,
            I => dti_counter_5
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__39064\,
            I => dti_counter_5
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__39061\,
            I => dti_counter_5
        );

    \I__7613\ : CascadeMux
    port map (
            O => \N__39054\,
            I => \N__39049\
        );

    \I__7612\ : CascadeMux
    port map (
            O => \N__39053\,
            I => \N__39046\
        );

    \I__7611\ : InMux
    port map (
            O => \N__39052\,
            I => \N__39043\
        );

    \I__7610\ : InMux
    port map (
            O => \N__39049\,
            I => \N__39040\
        );

    \I__7609\ : InMux
    port map (
            O => \N__39046\,
            I => \N__39037\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__39043\,
            I => dti_counter_6
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__39040\,
            I => dti_counter_6
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__39037\,
            I => dti_counter_6
        );

    \I__7605\ : CascadeMux
    port map (
            O => \N__39030\,
            I => \n14_adj_705_cascade_\
        );

    \I__7604\ : InMux
    port map (
            O => \N__39027\,
            I => \N__39022\
        );

    \I__7603\ : InMux
    port map (
            O => \N__39026\,
            I => \N__39017\
        );

    \I__7602\ : InMux
    port map (
            O => \N__39025\,
            I => \N__39017\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__39022\,
            I => dti_counter_2
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__39017\,
            I => dti_counter_2
        );

    \I__7599\ : InMux
    port map (
            O => \N__39012\,
            I => \N__39009\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__39009\,
            I => n10_adj_706
        );

    \I__7597\ : CascadeMux
    port map (
            O => \N__39006\,
            I => \N__39003\
        );

    \I__7596\ : InMux
    port map (
            O => \N__39003\,
            I => \N__38998\
        );

    \I__7595\ : InMux
    port map (
            O => \N__39002\,
            I => \N__38995\
        );

    \I__7594\ : InMux
    port map (
            O => \N__39001\,
            I => \N__38992\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__38998\,
            I => dti_counter_0
        );

    \I__7592\ : LocalMux
    port map (
            O => \N__38995\,
            I => dti_counter_0
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__38992\,
            I => dti_counter_0
        );

    \I__7590\ : InMux
    port map (
            O => \N__38985\,
            I => \N__38982\
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__38982\,
            I => n15081
        );

    \I__7588\ : CascadeMux
    port map (
            O => \N__38979\,
            I => \N__38976\
        );

    \I__7587\ : InMux
    port map (
            O => \N__38976\,
            I => \N__38971\
        );

    \I__7586\ : InMux
    port map (
            O => \N__38975\,
            I => \N__38966\
        );

    \I__7585\ : InMux
    port map (
            O => \N__38974\,
            I => \N__38966\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__38971\,
            I => dti_counter_3
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__38966\,
            I => dti_counter_3
        );

    \I__7582\ : InMux
    port map (
            O => \N__38961\,
            I => \N__38958\
        );

    \I__7581\ : LocalMux
    port map (
            O => \N__38958\,
            I => n15074
        );

    \I__7580\ : CascadeMux
    port map (
            O => \N__38955\,
            I => \N__38951\
        );

    \I__7579\ : InMux
    port map (
            O => \N__38954\,
            I => \N__38947\
        );

    \I__7578\ : InMux
    port map (
            O => \N__38951\,
            I => \N__38942\
        );

    \I__7577\ : InMux
    port map (
            O => \N__38950\,
            I => \N__38942\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__38947\,
            I => dti_counter_4
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__38942\,
            I => dti_counter_4
        );

    \I__7574\ : InMux
    port map (
            O => \N__38937\,
            I => \N__38934\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__38934\,
            I => n15073
        );

    \I__7572\ : CascadeMux
    port map (
            O => \N__38931\,
            I => \N__38928\
        );

    \I__7571\ : InMux
    port map (
            O => \N__38928\,
            I => \N__38924\
        );

    \I__7570\ : InMux
    port map (
            O => \N__38927\,
            I => \N__38920\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__38924\,
            I => \N__38917\
        );

    \I__7568\ : InMux
    port map (
            O => \N__38923\,
            I => \N__38914\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__38920\,
            I => dti_counter_7
        );

    \I__7566\ : Odrv4
    port map (
            O => \N__38917\,
            I => dti_counter_7
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__38914\,
            I => dti_counter_7
        );

    \I__7564\ : CascadeMux
    port map (
            O => \N__38907\,
            I => \N__38904\
        );

    \I__7563\ : InMux
    port map (
            O => \N__38904\,
            I => \N__38901\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__38901\,
            I => \N__38898\
        );

    \I__7561\ : Odrv4
    port map (
            O => \N__38898\,
            I => n15070
        );

    \I__7560\ : InMux
    port map (
            O => \N__38895\,
            I => \N__38892\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__38892\,
            I => \N__38889\
        );

    \I__7558\ : Span4Mux_v
    port map (
            O => \N__38889\,
            I => \N__38886\
        );

    \I__7557\ : Sp12to4
    port map (
            O => \N__38886\,
            I => \N__38882\
        );

    \I__7556\ : InMux
    port map (
            O => \N__38885\,
            I => \N__38879\
        );

    \I__7555\ : Odrv12
    port map (
            O => \N__38882\,
            I => \reg_B_1\
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__38879\,
            I => \reg_B_1\
        );

    \I__7553\ : InMux
    port map (
            O => \N__38874\,
            I => \N__38871\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__38871\,
            I => \N__38867\
        );

    \I__7551\ : InMux
    port map (
            O => \N__38870\,
            I => \N__38864\
        );

    \I__7550\ : Span4Mux_h
    port map (
            O => \N__38867\,
            I => \N__38861\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__38864\,
            I => \N__38858\
        );

    \I__7548\ : Span4Mux_h
    port map (
            O => \N__38861\,
            I => \N__38854\
        );

    \I__7547\ : Span4Mux_v
    port map (
            O => \N__38858\,
            I => \N__38851\
        );

    \I__7546\ : InMux
    port map (
            O => \N__38857\,
            I => \N__38848\
        );

    \I__7545\ : Odrv4
    port map (
            O => \N__38854\,
            I => n14129
        );

    \I__7544\ : Odrv4
    port map (
            O => \N__38851\,
            I => n14129
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__38848\,
            I => n14129
        );

    \I__7542\ : CascadeMux
    port map (
            O => \N__38841\,
            I => \N__38838\
        );

    \I__7541\ : InMux
    port map (
            O => \N__38838\,
            I => \N__38835\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__38835\,
            I => \N__38832\
        );

    \I__7539\ : Odrv4
    port map (
            O => \N__38832\,
            I => n1377
        );

    \I__7538\ : InMux
    port map (
            O => \N__38829\,
            I => \bfn_9_29_0_\
        );

    \I__7537\ : InMux
    port map (
            O => \N__38826\,
            I => n13006
        );

    \I__7536\ : InMux
    port map (
            O => \N__38823\,
            I => n13007
        );

    \I__7535\ : InMux
    port map (
            O => \N__38820\,
            I => n13008
        );

    \I__7534\ : InMux
    port map (
            O => \N__38817\,
            I => n13009
        );

    \I__7533\ : InMux
    port map (
            O => \N__38814\,
            I => \N__38811\
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__38811\,
            I => n15072
        );

    \I__7531\ : InMux
    port map (
            O => \N__38808\,
            I => n13010
        );

    \I__7530\ : InMux
    port map (
            O => \N__38805\,
            I => n13011
        );

    \I__7529\ : CascadeMux
    port map (
            O => \N__38802\,
            I => \N__38796\
        );

    \I__7528\ : CascadeMux
    port map (
            O => \N__38801\,
            I => \N__38792\
        );

    \I__7527\ : CascadeMux
    port map (
            O => \N__38800\,
            I => \N__38788\
        );

    \I__7526\ : InMux
    port map (
            O => \N__38799\,
            I => \N__38772\
        );

    \I__7525\ : InMux
    port map (
            O => \N__38796\,
            I => \N__38772\
        );

    \I__7524\ : InMux
    port map (
            O => \N__38795\,
            I => \N__38772\
        );

    \I__7523\ : InMux
    port map (
            O => \N__38792\,
            I => \N__38772\
        );

    \I__7522\ : InMux
    port map (
            O => \N__38791\,
            I => \N__38772\
        );

    \I__7521\ : InMux
    port map (
            O => \N__38788\,
            I => \N__38772\
        );

    \I__7520\ : InMux
    port map (
            O => \N__38787\,
            I => \N__38772\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__38772\,
            I => \N__38769\
        );

    \I__7518\ : Odrv4
    port map (
            O => \N__38769\,
            I => n11526
        );

    \I__7517\ : InMux
    port map (
            O => \N__38766\,
            I => n13012
        );

    \I__7516\ : InMux
    port map (
            O => \N__38763\,
            I => \N__38760\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__38760\,
            I => \N__38757\
        );

    \I__7514\ : Odrv4
    port map (
            O => \N__38757\,
            I => encoder0_position_scaled_18
        );

    \I__7513\ : InMux
    port map (
            O => \N__38754\,
            I => \N__38751\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__38751\,
            I => \N__38748\
        );

    \I__7511\ : Odrv4
    port map (
            O => \N__38748\,
            I => encoder0_position_scaled_23
        );

    \I__7510\ : InMux
    port map (
            O => \N__38745\,
            I => \N__38742\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__38742\,
            I => \N__38739\
        );

    \I__7508\ : Odrv4
    port map (
            O => \N__38739\,
            I => encoder0_position_scaled_17
        );

    \I__7507\ : CascadeMux
    port map (
            O => \N__38736\,
            I => \dti_N_333_cascade_\
        );

    \I__7506\ : InMux
    port map (
            O => \N__38733\,
            I => n13004
        );

    \I__7505\ : InMux
    port map (
            O => \N__38730\,
            I => n13005
        );

    \I__7504\ : InMux
    port map (
            O => \N__38727\,
            I => \N__38724\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__38724\,
            I => \N__38721\
        );

    \I__7502\ : Odrv4
    port map (
            O => \N__38721\,
            I => encoder0_position_scaled_8
        );

    \I__7501\ : InMux
    port map (
            O => \N__38718\,
            I => \N__38715\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__38715\,
            I => \N__38712\
        );

    \I__7499\ : Odrv4
    port map (
            O => \N__38712\,
            I => encoder0_position_scaled_14
        );

    \I__7498\ : InMux
    port map (
            O => \N__38709\,
            I => \N__38706\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__38706\,
            I => \N__38703\
        );

    \I__7496\ : Odrv4
    port map (
            O => \N__38703\,
            I => encoder0_position_scaled_10
        );

    \I__7495\ : InMux
    port map (
            O => \N__38700\,
            I => \N__38697\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__38697\,
            I => \N__38694\
        );

    \I__7493\ : Odrv4
    port map (
            O => \N__38694\,
            I => encoder0_position_scaled_12
        );

    \I__7492\ : InMux
    port map (
            O => \N__38691\,
            I => \N__38688\
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__38688\,
            I => \N__38685\
        );

    \I__7490\ : Odrv4
    port map (
            O => \N__38685\,
            I => encoder0_position_scaled_13
        );

    \I__7489\ : InMux
    port map (
            O => \N__38682\,
            I => \N__38679\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__38679\,
            I => \N__38676\
        );

    \I__7487\ : Odrv4
    port map (
            O => \N__38676\,
            I => encoder0_position_scaled_15
        );

    \I__7486\ : InMux
    port map (
            O => \N__38673\,
            I => \N__38670\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__38670\,
            I => \N__38667\
        );

    \I__7484\ : Odrv4
    port map (
            O => \N__38667\,
            I => n15508
        );

    \I__7483\ : InMux
    port map (
            O => \N__38664\,
            I => n12995
        );

    \I__7482\ : InMux
    port map (
            O => \N__38661\,
            I => n12996
        );

    \I__7481\ : InMux
    port map (
            O => \N__38658\,
            I => n12997
        );

    \I__7480\ : InMux
    port map (
            O => \N__38655\,
            I => \bfn_9_25_0_\
        );

    \I__7479\ : InMux
    port map (
            O => \N__38652\,
            I => n12999
        );

    \I__7478\ : InMux
    port map (
            O => \N__38649\,
            I => n13000
        );

    \I__7477\ : InMux
    port map (
            O => \N__38646\,
            I => n13001
        );

    \I__7476\ : InMux
    port map (
            O => \N__38643\,
            I => n13002
        );

    \I__7475\ : InMux
    port map (
            O => \N__38640\,
            I => \N__38637\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__38637\,
            I => \N__38634\
        );

    \I__7473\ : Span4Mux_v
    port map (
            O => \N__38634\,
            I => \N__38631\
        );

    \I__7472\ : Odrv4
    port map (
            O => \N__38631\,
            I => n4_adj_622
        );

    \I__7471\ : InMux
    port map (
            O => \N__38628\,
            I => n13003
        );

    \I__7470\ : InMux
    port map (
            O => \N__38625\,
            I => \N__38622\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__38622\,
            I => \N__38619\
        );

    \I__7468\ : Span4Mux_h
    port map (
            O => \N__38619\,
            I => \N__38616\
        );

    \I__7467\ : Odrv4
    port map (
            O => \N__38616\,
            I => n20
        );

    \I__7466\ : InMux
    port map (
            O => \N__38613\,
            I => n12987
        );

    \I__7465\ : CascadeMux
    port map (
            O => \N__38610\,
            I => \N__38607\
        );

    \I__7464\ : InMux
    port map (
            O => \N__38607\,
            I => \N__38604\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__38604\,
            I => \N__38601\
        );

    \I__7462\ : Odrv4
    port map (
            O => \N__38601\,
            I => n19_adj_637
        );

    \I__7461\ : InMux
    port map (
            O => \N__38598\,
            I => \N__38595\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__38595\,
            I => \N__38592\
        );

    \I__7459\ : Odrv12
    port map (
            O => \N__38592\,
            I => n19
        );

    \I__7458\ : InMux
    port map (
            O => \N__38589\,
            I => n12988
        );

    \I__7457\ : CascadeMux
    port map (
            O => \N__38586\,
            I => \N__38583\
        );

    \I__7456\ : InMux
    port map (
            O => \N__38583\,
            I => \N__38580\
        );

    \I__7455\ : LocalMux
    port map (
            O => \N__38580\,
            I => \N__38577\
        );

    \I__7454\ : Odrv4
    port map (
            O => \N__38577\,
            I => n18_adj_636
        );

    \I__7453\ : InMux
    port map (
            O => \N__38574\,
            I => \N__38571\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__38571\,
            I => \N__38568\
        );

    \I__7451\ : Span4Mux_h
    port map (
            O => \N__38568\,
            I => \N__38565\
        );

    \I__7450\ : Odrv4
    port map (
            O => \N__38565\,
            I => n18
        );

    \I__7449\ : InMux
    port map (
            O => \N__38562\,
            I => n12989
        );

    \I__7448\ : InMux
    port map (
            O => \N__38559\,
            I => \bfn_9_24_0_\
        );

    \I__7447\ : InMux
    port map (
            O => \N__38556\,
            I => n12991
        );

    \I__7446\ : InMux
    port map (
            O => \N__38553\,
            I => n12992
        );

    \I__7445\ : CascadeMux
    port map (
            O => \N__38550\,
            I => \N__38547\
        );

    \I__7444\ : InMux
    port map (
            O => \N__38547\,
            I => \N__38544\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__38544\,
            I => \N__38541\
        );

    \I__7442\ : Odrv12
    port map (
            O => \N__38541\,
            I => n14_adj_632
        );

    \I__7441\ : InMux
    port map (
            O => \N__38538\,
            I => \N__38535\
        );

    \I__7440\ : LocalMux
    port map (
            O => \N__38535\,
            I => \N__38532\
        );

    \I__7439\ : Odrv12
    port map (
            O => \N__38532\,
            I => n14
        );

    \I__7438\ : InMux
    port map (
            O => \N__38529\,
            I => n12993
        );

    \I__7437\ : InMux
    port map (
            O => \N__38526\,
            I => n12994
        );

    \I__7436\ : CascadeMux
    port map (
            O => \N__38523\,
            I => \N__38520\
        );

    \I__7435\ : InMux
    port map (
            O => \N__38520\,
            I => \N__38517\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__38517\,
            I => \N__38514\
        );

    \I__7433\ : Odrv12
    port map (
            O => \N__38514\,
            I => n28_adj_646
        );

    \I__7432\ : InMux
    port map (
            O => \N__38511\,
            I => \N__38508\
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__38508\,
            I => \N__38505\
        );

    \I__7430\ : Odrv4
    port map (
            O => \N__38505\,
            I => n28
        );

    \I__7429\ : InMux
    port map (
            O => \N__38502\,
            I => n12979
        );

    \I__7428\ : CascadeMux
    port map (
            O => \N__38499\,
            I => \N__38496\
        );

    \I__7427\ : InMux
    port map (
            O => \N__38496\,
            I => \N__38493\
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__38493\,
            I => n27_adj_645
        );

    \I__7425\ : InMux
    port map (
            O => \N__38490\,
            I => \N__38487\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__38487\,
            I => \N__38484\
        );

    \I__7423\ : Odrv4
    port map (
            O => \N__38484\,
            I => n27
        );

    \I__7422\ : InMux
    port map (
            O => \N__38481\,
            I => n12980
        );

    \I__7421\ : CascadeMux
    port map (
            O => \N__38478\,
            I => \N__38475\
        );

    \I__7420\ : InMux
    port map (
            O => \N__38475\,
            I => \N__38472\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__38472\,
            I => n26_adj_644
        );

    \I__7418\ : InMux
    port map (
            O => \N__38469\,
            I => \N__38466\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__38466\,
            I => \N__38463\
        );

    \I__7416\ : Span4Mux_h
    port map (
            O => \N__38463\,
            I => \N__38460\
        );

    \I__7415\ : Odrv4
    port map (
            O => \N__38460\,
            I => n26
        );

    \I__7414\ : InMux
    port map (
            O => \N__38457\,
            I => n12981
        );

    \I__7413\ : CascadeMux
    port map (
            O => \N__38454\,
            I => \N__38451\
        );

    \I__7412\ : InMux
    port map (
            O => \N__38451\,
            I => \N__38448\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__38448\,
            I => \N__38445\
        );

    \I__7410\ : Odrv4
    port map (
            O => \N__38445\,
            I => n25_adj_643
        );

    \I__7409\ : InMux
    port map (
            O => \N__38442\,
            I => \N__38439\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__38439\,
            I => \N__38436\
        );

    \I__7407\ : Span4Mux_h
    port map (
            O => \N__38436\,
            I => \N__38433\
        );

    \I__7406\ : Odrv4
    port map (
            O => \N__38433\,
            I => n25
        );

    \I__7405\ : InMux
    port map (
            O => \N__38430\,
            I => \bfn_9_23_0_\
        );

    \I__7404\ : CascadeMux
    port map (
            O => \N__38427\,
            I => \N__38424\
        );

    \I__7403\ : InMux
    port map (
            O => \N__38424\,
            I => \N__38421\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__38421\,
            I => \N__38418\
        );

    \I__7401\ : Odrv4
    port map (
            O => \N__38418\,
            I => n24_adj_642
        );

    \I__7400\ : InMux
    port map (
            O => \N__38415\,
            I => \N__38412\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__38412\,
            I => \N__38409\
        );

    \I__7398\ : Span4Mux_v
    port map (
            O => \N__38409\,
            I => \N__38406\
        );

    \I__7397\ : Odrv4
    port map (
            O => \N__38406\,
            I => n24
        );

    \I__7396\ : InMux
    port map (
            O => \N__38403\,
            I => n12983
        );

    \I__7395\ : CascadeMux
    port map (
            O => \N__38400\,
            I => \N__38397\
        );

    \I__7394\ : InMux
    port map (
            O => \N__38397\,
            I => \N__38394\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__38394\,
            I => \N__38391\
        );

    \I__7392\ : Odrv4
    port map (
            O => \N__38391\,
            I => n23_adj_641
        );

    \I__7391\ : InMux
    port map (
            O => \N__38388\,
            I => \N__38385\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__38385\,
            I => \N__38382\
        );

    \I__7389\ : Odrv4
    port map (
            O => \N__38382\,
            I => n23
        );

    \I__7388\ : InMux
    port map (
            O => \N__38379\,
            I => n12984
        );

    \I__7387\ : InMux
    port map (
            O => \N__38376\,
            I => \N__38373\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__38373\,
            I => \N__38370\
        );

    \I__7385\ : Odrv4
    port map (
            O => \N__38370\,
            I => n22
        );

    \I__7384\ : InMux
    port map (
            O => \N__38367\,
            I => n12985
        );

    \I__7383\ : InMux
    port map (
            O => \N__38364\,
            I => \N__38361\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__38361\,
            I => \N__38358\
        );

    \I__7381\ : Span4Mux_h
    port map (
            O => \N__38358\,
            I => \N__38355\
        );

    \I__7380\ : Odrv4
    port map (
            O => \N__38355\,
            I => n21
        );

    \I__7379\ : InMux
    port map (
            O => \N__38352\,
            I => n12986
        );

    \I__7378\ : InMux
    port map (
            O => \N__38349\,
            I => \N__38346\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__38346\,
            I => \N__38341\
        );

    \I__7376\ : InMux
    port map (
            O => \N__38345\,
            I => \N__38338\
        );

    \I__7375\ : InMux
    port map (
            O => \N__38344\,
            I => \N__38335\
        );

    \I__7374\ : Span4Mux_v
    port map (
            O => \N__38341\,
            I => \N__38330\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__38338\,
            I => \N__38330\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__38335\,
            I => \N__38327\
        );

    \I__7371\ : Span4Mux_h
    port map (
            O => \N__38330\,
            I => \N__38324\
        );

    \I__7370\ : Span4Mux_h
    port map (
            O => \N__38327\,
            I => \N__38321\
        );

    \I__7369\ : Span4Mux_h
    port map (
            O => \N__38324\,
            I => \N__38318\
        );

    \I__7368\ : Odrv4
    port map (
            O => \N__38321\,
            I => n309
        );

    \I__7367\ : Odrv4
    port map (
            O => \N__38318\,
            I => n309
        );

    \I__7366\ : CascadeMux
    port map (
            O => \N__38313\,
            I => \N__38310\
        );

    \I__7365\ : InMux
    port map (
            O => \N__38310\,
            I => \N__38307\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__38307\,
            I => \N__38304\
        );

    \I__7363\ : Odrv4
    port map (
            O => \N__38304\,
            I => n33_adj_651
        );

    \I__7362\ : InMux
    port map (
            O => \N__38301\,
            I => \N__38298\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__38298\,
            I => \N__38295\
        );

    \I__7360\ : Span4Mux_h
    port map (
            O => \N__38295\,
            I => \N__38292\
        );

    \I__7359\ : Odrv4
    port map (
            O => \N__38292\,
            I => n33
        );

    \I__7358\ : InMux
    port map (
            O => \N__38289\,
            I => \bfn_9_22_0_\
        );

    \I__7357\ : InMux
    port map (
            O => \N__38286\,
            I => \N__38283\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__38283\,
            I => \N__38280\
        );

    \I__7355\ : Odrv12
    port map (
            O => \N__38280\,
            I => n32
        );

    \I__7354\ : InMux
    port map (
            O => \N__38277\,
            I => n12975
        );

    \I__7353\ : CascadeMux
    port map (
            O => \N__38274\,
            I => \N__38271\
        );

    \I__7352\ : InMux
    port map (
            O => \N__38271\,
            I => \N__38268\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__38268\,
            I => \N__38265\
        );

    \I__7350\ : Odrv12
    port map (
            O => \N__38265\,
            I => n31_adj_649
        );

    \I__7349\ : InMux
    port map (
            O => \N__38262\,
            I => \N__38259\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__38259\,
            I => \N__38256\
        );

    \I__7347\ : Span4Mux_h
    port map (
            O => \N__38256\,
            I => \N__38253\
        );

    \I__7346\ : Odrv4
    port map (
            O => \N__38253\,
            I => n31
        );

    \I__7345\ : InMux
    port map (
            O => \N__38250\,
            I => n12976
        );

    \I__7344\ : CascadeMux
    port map (
            O => \N__38247\,
            I => \N__38244\
        );

    \I__7343\ : InMux
    port map (
            O => \N__38244\,
            I => \N__38241\
        );

    \I__7342\ : LocalMux
    port map (
            O => \N__38241\,
            I => n30_adj_648
        );

    \I__7341\ : InMux
    port map (
            O => \N__38238\,
            I => n12977
        );

    \I__7340\ : CascadeMux
    port map (
            O => \N__38235\,
            I => \N__38232\
        );

    \I__7339\ : InMux
    port map (
            O => \N__38232\,
            I => \N__38229\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__38229\,
            I => n29_adj_647
        );

    \I__7337\ : InMux
    port map (
            O => \N__38226\,
            I => \N__38223\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__38223\,
            I => \N__38220\
        );

    \I__7335\ : Span4Mux_h
    port map (
            O => \N__38220\,
            I => \N__38217\
        );

    \I__7334\ : Odrv4
    port map (
            O => \N__38217\,
            I => n29
        );

    \I__7333\ : InMux
    port map (
            O => \N__38214\,
            I => n12978
        );

    \I__7332\ : InMux
    port map (
            O => \N__38211\,
            I => \N__38207\
        );

    \I__7331\ : InMux
    port map (
            O => \N__38210\,
            I => \N__38203\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__38207\,
            I => \N__38200\
        );

    \I__7329\ : InMux
    port map (
            O => \N__38206\,
            I => \N__38197\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__38203\,
            I => \N__38194\
        );

    \I__7327\ : Span4Mux_h
    port map (
            O => \N__38200\,
            I => \N__38191\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__38197\,
            I => \N__38188\
        );

    \I__7325\ : Span4Mux_h
    port map (
            O => \N__38194\,
            I => \N__38185\
        );

    \I__7324\ : Span4Mux_h
    port map (
            O => \N__38191\,
            I => \N__38182\
        );

    \I__7323\ : Span12Mux_s8_h
    port map (
            O => \N__38188\,
            I => \N__38179\
        );

    \I__7322\ : Span4Mux_v
    port map (
            O => \N__38185\,
            I => \N__38176\
        );

    \I__7321\ : Odrv4
    port map (
            O => \N__38182\,
            I => n308
        );

    \I__7320\ : Odrv12
    port map (
            O => \N__38179\,
            I => n308
        );

    \I__7319\ : Odrv4
    port map (
            O => \N__38176\,
            I => n308
        );

    \I__7318\ : InMux
    port map (
            O => \N__38169\,
            I => \N__38166\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__38166\,
            I => \N__38163\
        );

    \I__7316\ : Odrv4
    port map (
            O => \N__38163\,
            I => n14530
        );

    \I__7315\ : InMux
    port map (
            O => \N__38160\,
            I => \N__38153\
        );

    \I__7314\ : InMux
    port map (
            O => \N__38159\,
            I => \N__38153\
        );

    \I__7313\ : InMux
    port map (
            O => \N__38158\,
            I => \N__38150\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__38153\,
            I => \N__38147\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__38150\,
            I => n1918
        );

    \I__7310\ : Odrv4
    port map (
            O => \N__38147\,
            I => n1918
        );

    \I__7309\ : InMux
    port map (
            O => \N__38142\,
            I => \N__38139\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__38139\,
            I => \N__38134\
        );

    \I__7307\ : InMux
    port map (
            O => \N__38138\,
            I => \N__38131\
        );

    \I__7306\ : InMux
    port map (
            O => \N__38137\,
            I => \N__38128\
        );

    \I__7305\ : Span4Mux_v
    port map (
            O => \N__38134\,
            I => \N__38123\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__38131\,
            I => \N__38123\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__38128\,
            I => n1919
        );

    \I__7302\ : Odrv4
    port map (
            O => \N__38123\,
            I => n1919
        );

    \I__7301\ : InMux
    port map (
            O => \N__38118\,
            I => \N__38114\
        );

    \I__7300\ : InMux
    port map (
            O => \N__38117\,
            I => \N__38111\
        );

    \I__7299\ : LocalMux
    port map (
            O => \N__38114\,
            I => \N__38108\
        );

    \I__7298\ : LocalMux
    port map (
            O => \N__38111\,
            I => \N__38102\
        );

    \I__7297\ : Span4Mux_v
    port map (
            O => \N__38108\,
            I => \N__38102\
        );

    \I__7296\ : InMux
    port map (
            O => \N__38107\,
            I => \N__38099\
        );

    \I__7295\ : Span4Mux_h
    port map (
            O => \N__38102\,
            I => \N__38096\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__38099\,
            I => \N__38093\
        );

    \I__7293\ : Odrv4
    port map (
            O => \N__38096\,
            I => n305
        );

    \I__7292\ : Odrv4
    port map (
            O => \N__38093\,
            I => n305
        );

    \I__7291\ : InMux
    port map (
            O => \N__38088\,
            I => \N__38084\
        );

    \I__7290\ : InMux
    port map (
            O => \N__38087\,
            I => \N__38081\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__38084\,
            I => \N__38075\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__38081\,
            I => \N__38075\
        );

    \I__7287\ : InMux
    port map (
            O => \N__38080\,
            I => \N__38072\
        );

    \I__7286\ : Span4Mux_v
    port map (
            O => \N__38075\,
            I => \N__38067\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__38072\,
            I => \N__38067\
        );

    \I__7284\ : Odrv4
    port map (
            O => \N__38067\,
            I => n306
        );

    \I__7283\ : InMux
    port map (
            O => \N__38064\,
            I => \N__38061\
        );

    \I__7282\ : LocalMux
    port map (
            O => \N__38061\,
            I => \N__38058\
        );

    \I__7281\ : Span4Mux_v
    port map (
            O => \N__38058\,
            I => \N__38055\
        );

    \I__7280\ : Odrv4
    port map (
            O => \N__38055\,
            I => n1991
        );

    \I__7279\ : InMux
    port map (
            O => \N__38052\,
            I => n12631
        );

    \I__7278\ : InMux
    port map (
            O => \N__38049\,
            I => \N__38046\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__38046\,
            I => \N__38043\
        );

    \I__7276\ : Span4Mux_v
    port map (
            O => \N__38043\,
            I => \N__38040\
        );

    \I__7275\ : Odrv4
    port map (
            O => \N__38040\,
            I => n1990
        );

    \I__7274\ : InMux
    port map (
            O => \N__38037\,
            I => n12632
        );

    \I__7273\ : CascadeMux
    port map (
            O => \N__38034\,
            I => \N__38031\
        );

    \I__7272\ : InMux
    port map (
            O => \N__38031\,
            I => \N__38028\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__38028\,
            I => \N__38024\
        );

    \I__7270\ : InMux
    port map (
            O => \N__38027\,
            I => \N__38021\
        );

    \I__7269\ : Odrv4
    port map (
            O => \N__38024\,
            I => n1922
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__38021\,
            I => n1922
        );

    \I__7267\ : InMux
    port map (
            O => \N__38016\,
            I => \N__38013\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__38013\,
            I => \N__38010\
        );

    \I__7265\ : Odrv4
    port map (
            O => \N__38010\,
            I => n1989
        );

    \I__7264\ : InMux
    port map (
            O => \N__38007\,
            I => n12633
        );

    \I__7263\ : CascadeMux
    port map (
            O => \N__38004\,
            I => \N__38001\
        );

    \I__7262\ : InMux
    port map (
            O => \N__38001\,
            I => \N__37998\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__37998\,
            I => \N__37995\
        );

    \I__7260\ : Odrv4
    port map (
            O => \N__37995\,
            I => n1988
        );

    \I__7259\ : InMux
    port map (
            O => \N__37992\,
            I => n12634
        );

    \I__7258\ : InMux
    port map (
            O => \N__37989\,
            I => n12635
        );

    \I__7257\ : CascadeMux
    port map (
            O => \N__37986\,
            I => \N__37983\
        );

    \I__7256\ : InMux
    port map (
            O => \N__37983\,
            I => \N__37980\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__37980\,
            I => \N__37977\
        );

    \I__7254\ : Span4Mux_h
    port map (
            O => \N__37977\,
            I => \N__37974\
        );

    \I__7253\ : Odrv4
    port map (
            O => \N__37974\,
            I => n1986
        );

    \I__7252\ : InMux
    port map (
            O => \N__37971\,
            I => n12636
        );

    \I__7251\ : InMux
    port map (
            O => \N__37968\,
            I => \N__37965\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__37965\,
            I => \N__37962\
        );

    \I__7249\ : Span4Mux_h
    port map (
            O => \N__37962\,
            I => \N__37959\
        );

    \I__7248\ : Odrv4
    port map (
            O => \N__37959\,
            I => n1985
        );

    \I__7247\ : InMux
    port map (
            O => \N__37956\,
            I => \bfn_9_18_0_\
        );

    \I__7246\ : CascadeMux
    port map (
            O => \N__37953\,
            I => \N__37949\
        );

    \I__7245\ : InMux
    port map (
            O => \N__37952\,
            I => \N__37946\
        );

    \I__7244\ : InMux
    port map (
            O => \N__37949\,
            I => \N__37943\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__37946\,
            I => \N__37940\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__37943\,
            I => \N__37937\
        );

    \I__7241\ : Odrv12
    port map (
            O => \N__37940\,
            I => n15674
        );

    \I__7240\ : Odrv4
    port map (
            O => \N__37937\,
            I => n15674
        );

    \I__7239\ : InMux
    port map (
            O => \N__37932\,
            I => n12638
        );

    \I__7238\ : CascadeMux
    port map (
            O => \N__37929\,
            I => \N__37926\
        );

    \I__7237\ : InMux
    port map (
            O => \N__37926\,
            I => \N__37920\
        );

    \I__7236\ : InMux
    port map (
            O => \N__37925\,
            I => \N__37920\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__37920\,
            I => \N__37917\
        );

    \I__7234\ : Span4Mux_h
    port map (
            O => \N__37917\,
            I => \N__37914\
        );

    \I__7233\ : Odrv4
    port map (
            O => \N__37914\,
            I => n2016
        );

    \I__7232\ : InMux
    port map (
            O => \N__37911\,
            I => \N__37908\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__37908\,
            I => \N__37903\
        );

    \I__7230\ : CascadeMux
    port map (
            O => \N__37907\,
            I => \N__37900\
        );

    \I__7229\ : InMux
    port map (
            O => \N__37906\,
            I => \N__37897\
        );

    \I__7228\ : Span4Mux_h
    port map (
            O => \N__37903\,
            I => \N__37894\
        );

    \I__7227\ : InMux
    port map (
            O => \N__37900\,
            I => \N__37891\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__37897\,
            I => \N__37888\
        );

    \I__7225\ : Odrv4
    port map (
            O => \N__37894\,
            I => n1921
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__37891\,
            I => n1921
        );

    \I__7223\ : Odrv4
    port map (
            O => \N__37888\,
            I => n1921
        );

    \I__7222\ : InMux
    port map (
            O => \N__37881\,
            I => \N__37878\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__37878\,
            I => \N__37875\
        );

    \I__7220\ : Span4Mux_v
    port map (
            O => \N__37875\,
            I => \N__37872\
        );

    \I__7219\ : Odrv4
    port map (
            O => \N__37872\,
            I => n1999
        );

    \I__7218\ : InMux
    port map (
            O => \N__37869\,
            I => n12623
        );

    \I__7217\ : InMux
    port map (
            O => \N__37866\,
            I => \N__37863\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__37863\,
            I => \N__37860\
        );

    \I__7215\ : Odrv4
    port map (
            O => \N__37860\,
            I => n1998
        );

    \I__7214\ : InMux
    port map (
            O => \N__37857\,
            I => n12624
        );

    \I__7213\ : CascadeMux
    port map (
            O => \N__37854\,
            I => \N__37851\
        );

    \I__7212\ : InMux
    port map (
            O => \N__37851\,
            I => \N__37848\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__37848\,
            I => \N__37845\
        );

    \I__7210\ : Span4Mux_v
    port map (
            O => \N__37845\,
            I => \N__37842\
        );

    \I__7209\ : Odrv4
    port map (
            O => \N__37842\,
            I => n1997
        );

    \I__7208\ : InMux
    port map (
            O => \N__37839\,
            I => n12625
        );

    \I__7207\ : CascadeMux
    port map (
            O => \N__37836\,
            I => \N__37833\
        );

    \I__7206\ : InMux
    port map (
            O => \N__37833\,
            I => \N__37830\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__37830\,
            I => \N__37827\
        );

    \I__7204\ : Span4Mux_h
    port map (
            O => \N__37827\,
            I => \N__37824\
        );

    \I__7203\ : Odrv4
    port map (
            O => \N__37824\,
            I => n1996
        );

    \I__7202\ : InMux
    port map (
            O => \N__37821\,
            I => n12626
        );

    \I__7201\ : CascadeMux
    port map (
            O => \N__37818\,
            I => \N__37815\
        );

    \I__7200\ : InMux
    port map (
            O => \N__37815\,
            I => \N__37812\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__37812\,
            I => \N__37809\
        );

    \I__7198\ : Span4Mux_h
    port map (
            O => \N__37809\,
            I => \N__37806\
        );

    \I__7197\ : Odrv4
    port map (
            O => \N__37806\,
            I => n1995
        );

    \I__7196\ : InMux
    port map (
            O => \N__37803\,
            I => n12627
        );

    \I__7195\ : InMux
    port map (
            O => \N__37800\,
            I => \N__37797\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__37797\,
            I => \N__37794\
        );

    \I__7193\ : Span4Mux_h
    port map (
            O => \N__37794\,
            I => \N__37791\
        );

    \I__7192\ : Odrv4
    port map (
            O => \N__37791\,
            I => n1994
        );

    \I__7191\ : InMux
    port map (
            O => \N__37788\,
            I => n12628
        );

    \I__7190\ : InMux
    port map (
            O => \N__37785\,
            I => \N__37782\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__37782\,
            I => \N__37779\
        );

    \I__7188\ : Span4Mux_h
    port map (
            O => \N__37779\,
            I => \N__37776\
        );

    \I__7187\ : Odrv4
    port map (
            O => \N__37776\,
            I => n1993
        );

    \I__7186\ : InMux
    port map (
            O => \N__37773\,
            I => \bfn_9_17_0_\
        );

    \I__7185\ : InMux
    port map (
            O => \N__37770\,
            I => \N__37767\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__37767\,
            I => \N__37764\
        );

    \I__7183\ : Span4Mux_h
    port map (
            O => \N__37764\,
            I => \N__37761\
        );

    \I__7182\ : Odrv4
    port map (
            O => \N__37761\,
            I => n1992
        );

    \I__7181\ : InMux
    port map (
            O => \N__37758\,
            I => n12630
        );

    \I__7180\ : InMux
    port map (
            O => \N__37755\,
            I => \N__37750\
        );

    \I__7179\ : InMux
    port map (
            O => \N__37754\,
            I => \N__37747\
        );

    \I__7178\ : InMux
    port map (
            O => \N__37753\,
            I => \N__37744\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__37750\,
            I => \N__37741\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__37747\,
            I => \N__37736\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__37744\,
            I => \N__37736\
        );

    \I__7174\ : Odrv4
    port map (
            O => \N__37741\,
            I => n3209
        );

    \I__7173\ : Odrv4
    port map (
            O => \N__37736\,
            I => n3209
        );

    \I__7172\ : CascadeMux
    port map (
            O => \N__37731\,
            I => \N__37728\
        );

    \I__7171\ : InMux
    port map (
            O => \N__37728\,
            I => \N__37725\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__37725\,
            I => \N__37722\
        );

    \I__7169\ : Odrv4
    port map (
            O => \N__37722\,
            I => n3276
        );

    \I__7168\ : InMux
    port map (
            O => \N__37719\,
            I => n12946
        );

    \I__7167\ : CascadeMux
    port map (
            O => \N__37716\,
            I => \N__37711\
        );

    \I__7166\ : InMux
    port map (
            O => \N__37715\,
            I => \N__37708\
        );

    \I__7165\ : InMux
    port map (
            O => \N__37714\,
            I => \N__37705\
        );

    \I__7164\ : InMux
    port map (
            O => \N__37711\,
            I => \N__37702\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__37708\,
            I => \N__37699\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__37705\,
            I => \N__37694\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__37702\,
            I => \N__37694\
        );

    \I__7160\ : Odrv4
    port map (
            O => \N__37699\,
            I => n3208
        );

    \I__7159\ : Odrv4
    port map (
            O => \N__37694\,
            I => n3208
        );

    \I__7158\ : InMux
    port map (
            O => \N__37689\,
            I => \N__37686\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__37686\,
            I => \N__37683\
        );

    \I__7156\ : Odrv4
    port map (
            O => \N__37683\,
            I => n3275
        );

    \I__7155\ : InMux
    port map (
            O => \N__37680\,
            I => n12947
        );

    \I__7154\ : InMux
    port map (
            O => \N__37677\,
            I => \N__37674\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__37674\,
            I => \N__37669\
        );

    \I__7152\ : InMux
    port map (
            O => \N__37673\,
            I => \N__37664\
        );

    \I__7151\ : InMux
    port map (
            O => \N__37672\,
            I => \N__37664\
        );

    \I__7150\ : Span4Mux_s2_v
    port map (
            O => \N__37669\,
            I => \N__37659\
        );

    \I__7149\ : LocalMux
    port map (
            O => \N__37664\,
            I => \N__37659\
        );

    \I__7148\ : Span4Mux_h
    port map (
            O => \N__37659\,
            I => \N__37656\
        );

    \I__7147\ : Odrv4
    port map (
            O => \N__37656\,
            I => n3207
        );

    \I__7146\ : InMux
    port map (
            O => \N__37653\,
            I => \N__37650\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__37650\,
            I => \N__37647\
        );

    \I__7144\ : Odrv4
    port map (
            O => \N__37647\,
            I => n3274
        );

    \I__7143\ : InMux
    port map (
            O => \N__37644\,
            I => n12948
        );

    \I__7142\ : InMux
    port map (
            O => \N__37641\,
            I => \N__37636\
        );

    \I__7141\ : InMux
    port map (
            O => \N__37640\,
            I => \N__37633\
        );

    \I__7140\ : InMux
    port map (
            O => \N__37639\,
            I => \N__37630\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__37636\,
            I => \N__37627\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__37633\,
            I => \N__37624\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__37630\,
            I => \N__37621\
        );

    \I__7136\ : Span4Mux_v
    port map (
            O => \N__37627\,
            I => \N__37614\
        );

    \I__7135\ : Span4Mux_h
    port map (
            O => \N__37624\,
            I => \N__37614\
        );

    \I__7134\ : Span4Mux_v
    port map (
            O => \N__37621\,
            I => \N__37614\
        );

    \I__7133\ : Odrv4
    port map (
            O => \N__37614\,
            I => n3206
        );

    \I__7132\ : InMux
    port map (
            O => \N__37611\,
            I => \N__37608\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__37608\,
            I => \N__37605\
        );

    \I__7130\ : Odrv4
    port map (
            O => \N__37605\,
            I => n3273
        );

    \I__7129\ : InMux
    port map (
            O => \N__37602\,
            I => n12949
        );

    \I__7128\ : InMux
    port map (
            O => \N__37599\,
            I => \N__37595\
        );

    \I__7127\ : InMux
    port map (
            O => \N__37598\,
            I => \N__37591\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__37595\,
            I => \N__37588\
        );

    \I__7125\ : InMux
    port map (
            O => \N__37594\,
            I => \N__37585\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__37591\,
            I => \N__37582\
        );

    \I__7123\ : Span4Mux_v
    port map (
            O => \N__37588\,
            I => \N__37579\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__37585\,
            I => \N__37576\
        );

    \I__7121\ : Span4Mux_h
    port map (
            O => \N__37582\,
            I => \N__37573\
        );

    \I__7120\ : Odrv4
    port map (
            O => \N__37579\,
            I => n3205
        );

    \I__7119\ : Odrv12
    port map (
            O => \N__37576\,
            I => n3205
        );

    \I__7118\ : Odrv4
    port map (
            O => \N__37573\,
            I => n3205
        );

    \I__7117\ : InMux
    port map (
            O => \N__37566\,
            I => \N__37563\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__37563\,
            I => \N__37560\
        );

    \I__7115\ : Odrv4
    port map (
            O => \N__37560\,
            I => n3272
        );

    \I__7114\ : InMux
    port map (
            O => \N__37557\,
            I => n12950
        );

    \I__7113\ : InMux
    port map (
            O => \N__37554\,
            I => \N__37551\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__37551\,
            I => \N__37546\
        );

    \I__7111\ : InMux
    port map (
            O => \N__37550\,
            I => \N__37543\
        );

    \I__7110\ : InMux
    port map (
            O => \N__37549\,
            I => \N__37540\
        );

    \I__7109\ : Span4Mux_v
    port map (
            O => \N__37546\,
            I => \N__37535\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__37543\,
            I => \N__37535\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__37540\,
            I => \N__37532\
        );

    \I__7106\ : Span4Mux_h
    port map (
            O => \N__37535\,
            I => \N__37529\
        );

    \I__7105\ : Odrv12
    port map (
            O => \N__37532\,
            I => n3204
        );

    \I__7104\ : Odrv4
    port map (
            O => \N__37529\,
            I => n3204
        );

    \I__7103\ : InMux
    port map (
            O => \N__37524\,
            I => n12951
        );

    \I__7102\ : CascadeMux
    port map (
            O => \N__37521\,
            I => \N__37518\
        );

    \I__7101\ : InMux
    port map (
            O => \N__37518\,
            I => \N__37515\
        );

    \I__7100\ : LocalMux
    port map (
            O => \N__37515\,
            I => \N__37512\
        );

    \I__7099\ : Span4Mux_h
    port map (
            O => \N__37512\,
            I => \N__37509\
        );

    \I__7098\ : Odrv4
    port map (
            O => \N__37509\,
            I => n3271
        );

    \I__7097\ : InMux
    port map (
            O => \N__37506\,
            I => \N__37503\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__37503\,
            I => \N__37500\
        );

    \I__7095\ : Span4Mux_v
    port map (
            O => \N__37500\,
            I => \N__37497\
        );

    \I__7094\ : Odrv4
    port map (
            O => \N__37497\,
            I => n2001
        );

    \I__7093\ : InMux
    port map (
            O => \N__37494\,
            I => \bfn_9_16_0_\
        );

    \I__7092\ : CascadeMux
    port map (
            O => \N__37491\,
            I => \N__37488\
        );

    \I__7091\ : InMux
    port map (
            O => \N__37488\,
            I => \N__37485\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__37485\,
            I => \N__37482\
        );

    \I__7089\ : Span4Mux_v
    port map (
            O => \N__37482\,
            I => \N__37479\
        );

    \I__7088\ : Odrv4
    port map (
            O => \N__37479\,
            I => n2000
        );

    \I__7087\ : InMux
    port map (
            O => \N__37476\,
            I => n12622
        );

    \I__7086\ : InMux
    port map (
            O => \N__37473\,
            I => \N__37468\
        );

    \I__7085\ : CascadeMux
    port map (
            O => \N__37472\,
            I => \N__37465\
        );

    \I__7084\ : InMux
    port map (
            O => \N__37471\,
            I => \N__37462\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__37468\,
            I => \N__37459\
        );

    \I__7082\ : InMux
    port map (
            O => \N__37465\,
            I => \N__37456\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__37462\,
            I => n3217
        );

    \I__7080\ : Odrv4
    port map (
            O => \N__37459\,
            I => n3217
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__37456\,
            I => n3217
        );

    \I__7078\ : InMux
    port map (
            O => \N__37449\,
            I => \N__37446\
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__37446\,
            I => \N__37443\
        );

    \I__7076\ : Odrv4
    port map (
            O => \N__37443\,
            I => n3284
        );

    \I__7075\ : InMux
    port map (
            O => \N__37440\,
            I => n12938
        );

    \I__7074\ : InMux
    port map (
            O => \N__37437\,
            I => \N__37433\
        );

    \I__7073\ : InMux
    port map (
            O => \N__37436\,
            I => \N__37429\
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__37433\,
            I => \N__37426\
        );

    \I__7071\ : InMux
    port map (
            O => \N__37432\,
            I => \N__37423\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__37429\,
            I => n3216
        );

    \I__7069\ : Odrv12
    port map (
            O => \N__37426\,
            I => n3216
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__37423\,
            I => n3216
        );

    \I__7067\ : InMux
    port map (
            O => \N__37416\,
            I => \N__37413\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__37413\,
            I => \N__37410\
        );

    \I__7065\ : Odrv4
    port map (
            O => \N__37410\,
            I => n3283
        );

    \I__7064\ : InMux
    port map (
            O => \N__37407\,
            I => n12939
        );

    \I__7063\ : InMux
    port map (
            O => \N__37404\,
            I => \N__37400\
        );

    \I__7062\ : InMux
    port map (
            O => \N__37403\,
            I => \N__37396\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__37400\,
            I => \N__37393\
        );

    \I__7060\ : InMux
    port map (
            O => \N__37399\,
            I => \N__37390\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__37396\,
            I => n3215
        );

    \I__7058\ : Odrv4
    port map (
            O => \N__37393\,
            I => n3215
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__37390\,
            I => n3215
        );

    \I__7056\ : InMux
    port map (
            O => \N__37383\,
            I => \N__37380\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__37380\,
            I => n3282
        );

    \I__7054\ : InMux
    port map (
            O => \N__37377\,
            I => n12940
        );

    \I__7053\ : InMux
    port map (
            O => \N__37374\,
            I => \N__37370\
        );

    \I__7052\ : InMux
    port map (
            O => \N__37373\,
            I => \N__37367\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__37370\,
            I => \N__37361\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__37367\,
            I => \N__37361\
        );

    \I__7049\ : InMux
    port map (
            O => \N__37366\,
            I => \N__37358\
        );

    \I__7048\ : Span4Mux_h
    port map (
            O => \N__37361\,
            I => \N__37353\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__37358\,
            I => \N__37353\
        );

    \I__7046\ : Odrv4
    port map (
            O => \N__37353\,
            I => n3214
        );

    \I__7045\ : InMux
    port map (
            O => \N__37350\,
            I => \N__37347\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__37347\,
            I => n3281
        );

    \I__7043\ : InMux
    port map (
            O => \N__37344\,
            I => n12941
        );

    \I__7042\ : InMux
    port map (
            O => \N__37341\,
            I => \N__37337\
        );

    \I__7041\ : InMux
    port map (
            O => \N__37340\,
            I => \N__37334\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__37337\,
            I => \N__37328\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__37334\,
            I => \N__37328\
        );

    \I__7038\ : InMux
    port map (
            O => \N__37333\,
            I => \N__37325\
        );

    \I__7037\ : Odrv12
    port map (
            O => \N__37328\,
            I => n3213
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__37325\,
            I => n3213
        );

    \I__7035\ : CascadeMux
    port map (
            O => \N__37320\,
            I => \N__37317\
        );

    \I__7034\ : InMux
    port map (
            O => \N__37317\,
            I => \N__37314\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__37314\,
            I => n3280
        );

    \I__7032\ : InMux
    port map (
            O => \N__37311\,
            I => n12942
        );

    \I__7031\ : CascadeMux
    port map (
            O => \N__37308\,
            I => \N__37304\
        );

    \I__7030\ : InMux
    port map (
            O => \N__37307\,
            I => \N__37301\
        );

    \I__7029\ : InMux
    port map (
            O => \N__37304\,
            I => \N__37298\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__37301\,
            I => \N__37293\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__37298\,
            I => \N__37293\
        );

    \I__7026\ : Odrv4
    port map (
            O => \N__37293\,
            I => n3212
        );

    \I__7025\ : InMux
    port map (
            O => \N__37290\,
            I => \N__37287\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__37287\,
            I => n3279
        );

    \I__7023\ : InMux
    port map (
            O => \N__37284\,
            I => n12943
        );

    \I__7022\ : InMux
    port map (
            O => \N__37281\,
            I => \N__37278\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__37278\,
            I => \N__37274\
        );

    \I__7020\ : InMux
    port map (
            O => \N__37277\,
            I => \N__37270\
        );

    \I__7019\ : Span4Mux_s2_v
    port map (
            O => \N__37274\,
            I => \N__37267\
        );

    \I__7018\ : InMux
    port map (
            O => \N__37273\,
            I => \N__37264\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__37270\,
            I => n3211
        );

    \I__7016\ : Odrv4
    port map (
            O => \N__37267\,
            I => n3211
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__37264\,
            I => n3211
        );

    \I__7014\ : InMux
    port map (
            O => \N__37257\,
            I => \N__37254\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__37254\,
            I => n3278
        );

    \I__7012\ : InMux
    port map (
            O => \N__37251\,
            I => \bfn_7_32_0_\
        );

    \I__7011\ : InMux
    port map (
            O => \N__37248\,
            I => \N__37243\
        );

    \I__7010\ : InMux
    port map (
            O => \N__37247\,
            I => \N__37240\
        );

    \I__7009\ : InMux
    port map (
            O => \N__37246\,
            I => \N__37237\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__37243\,
            I => \N__37234\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__37240\,
            I => \N__37231\
        );

    \I__7006\ : LocalMux
    port map (
            O => \N__37237\,
            I => n3210
        );

    \I__7005\ : Odrv4
    port map (
            O => \N__37234\,
            I => n3210
        );

    \I__7004\ : Odrv4
    port map (
            O => \N__37231\,
            I => n3210
        );

    \I__7003\ : InMux
    port map (
            O => \N__37224\,
            I => \N__37221\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__37221\,
            I => \N__37218\
        );

    \I__7001\ : Odrv4
    port map (
            O => \N__37218\,
            I => n3277
        );

    \I__7000\ : InMux
    port map (
            O => \N__37215\,
            I => n12945
        );

    \I__6999\ : CascadeMux
    port map (
            O => \N__37212\,
            I => \N__37208\
        );

    \I__6998\ : CascadeMux
    port map (
            O => \N__37211\,
            I => \N__37204\
        );

    \I__6997\ : InMux
    port map (
            O => \N__37208\,
            I => \N__37201\
        );

    \I__6996\ : InMux
    port map (
            O => \N__37207\,
            I => \N__37198\
        );

    \I__6995\ : InMux
    port map (
            O => \N__37204\,
            I => \N__37195\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__37201\,
            I => \N__37192\
        );

    \I__6993\ : LocalMux
    port map (
            O => \N__37198\,
            I => n3225
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__37195\,
            I => n3225
        );

    \I__6991\ : Odrv4
    port map (
            O => \N__37192\,
            I => n3225
        );

    \I__6990\ : InMux
    port map (
            O => \N__37185\,
            I => \N__37182\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__37182\,
            I => n3292
        );

    \I__6988\ : InMux
    port map (
            O => \N__37179\,
            I => n12930
        );

    \I__6987\ : CascadeMux
    port map (
            O => \N__37176\,
            I => \N__37173\
        );

    \I__6986\ : InMux
    port map (
            O => \N__37173\,
            I => \N__37169\
        );

    \I__6985\ : CascadeMux
    port map (
            O => \N__37172\,
            I => \N__37166\
        );

    \I__6984\ : LocalMux
    port map (
            O => \N__37169\,
            I => \N__37162\
        );

    \I__6983\ : InMux
    port map (
            O => \N__37166\,
            I => \N__37157\
        );

    \I__6982\ : InMux
    port map (
            O => \N__37165\,
            I => \N__37157\
        );

    \I__6981\ : Odrv4
    port map (
            O => \N__37162\,
            I => n3224
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__37157\,
            I => n3224
        );

    \I__6979\ : InMux
    port map (
            O => \N__37152\,
            I => \N__37149\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__37149\,
            I => \N__37146\
        );

    \I__6977\ : Odrv4
    port map (
            O => \N__37146\,
            I => n3291
        );

    \I__6976\ : InMux
    port map (
            O => \N__37143\,
            I => n12931
        );

    \I__6975\ : CascadeMux
    port map (
            O => \N__37140\,
            I => \N__37136\
        );

    \I__6974\ : InMux
    port map (
            O => \N__37139\,
            I => \N__37133\
        );

    \I__6973\ : InMux
    port map (
            O => \N__37136\,
            I => \N__37130\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__37133\,
            I => \N__37126\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__37130\,
            I => \N__37123\
        );

    \I__6970\ : InMux
    port map (
            O => \N__37129\,
            I => \N__37120\
        );

    \I__6969\ : Odrv4
    port map (
            O => \N__37126\,
            I => n3223
        );

    \I__6968\ : Odrv4
    port map (
            O => \N__37123\,
            I => n3223
        );

    \I__6967\ : LocalMux
    port map (
            O => \N__37120\,
            I => n3223
        );

    \I__6966\ : InMux
    port map (
            O => \N__37113\,
            I => \N__37110\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__37110\,
            I => \N__37107\
        );

    \I__6964\ : Span4Mux_s2_v
    port map (
            O => \N__37107\,
            I => \N__37104\
        );

    \I__6963\ : Odrv4
    port map (
            O => \N__37104\,
            I => n3290
        );

    \I__6962\ : InMux
    port map (
            O => \N__37101\,
            I => n12932
        );

    \I__6961\ : CascadeMux
    port map (
            O => \N__37098\,
            I => \N__37095\
        );

    \I__6960\ : InMux
    port map (
            O => \N__37095\,
            I => \N__37091\
        );

    \I__6959\ : InMux
    port map (
            O => \N__37094\,
            I => \N__37087\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__37091\,
            I => \N__37084\
        );

    \I__6957\ : InMux
    port map (
            O => \N__37090\,
            I => \N__37081\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__37087\,
            I => n3222
        );

    \I__6955\ : Odrv4
    port map (
            O => \N__37084\,
            I => n3222
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__37081\,
            I => n3222
        );

    \I__6953\ : InMux
    port map (
            O => \N__37074\,
            I => \N__37071\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__37071\,
            I => \N__37068\
        );

    \I__6951\ : Span4Mux_s2_v
    port map (
            O => \N__37068\,
            I => \N__37065\
        );

    \I__6950\ : Odrv4
    port map (
            O => \N__37065\,
            I => n3289
        );

    \I__6949\ : InMux
    port map (
            O => \N__37062\,
            I => n12933
        );

    \I__6948\ : CascadeMux
    port map (
            O => \N__37059\,
            I => \N__37055\
        );

    \I__6947\ : CascadeMux
    port map (
            O => \N__37058\,
            I => \N__37052\
        );

    \I__6946\ : InMux
    port map (
            O => \N__37055\,
            I => \N__37049\
        );

    \I__6945\ : InMux
    port map (
            O => \N__37052\,
            I => \N__37045\
        );

    \I__6944\ : LocalMux
    port map (
            O => \N__37049\,
            I => \N__37042\
        );

    \I__6943\ : InMux
    port map (
            O => \N__37048\,
            I => \N__37039\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__37045\,
            I => n3221
        );

    \I__6941\ : Odrv4
    port map (
            O => \N__37042\,
            I => n3221
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__37039\,
            I => n3221
        );

    \I__6939\ : InMux
    port map (
            O => \N__37032\,
            I => \N__37029\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__37029\,
            I => n3288
        );

    \I__6937\ : InMux
    port map (
            O => \N__37026\,
            I => n12934
        );

    \I__6936\ : CascadeMux
    port map (
            O => \N__37023\,
            I => \N__37020\
        );

    \I__6935\ : InMux
    port map (
            O => \N__37020\,
            I => \N__37016\
        );

    \I__6934\ : InMux
    port map (
            O => \N__37019\,
            I => \N__37012\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__37016\,
            I => \N__37009\
        );

    \I__6932\ : InMux
    port map (
            O => \N__37015\,
            I => \N__37006\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__37012\,
            I => n3220
        );

    \I__6930\ : Odrv4
    port map (
            O => \N__37009\,
            I => n3220
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__37006\,
            I => n3220
        );

    \I__6928\ : InMux
    port map (
            O => \N__36999\,
            I => \N__36996\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__36996\,
            I => \N__36993\
        );

    \I__6926\ : Odrv12
    port map (
            O => \N__36993\,
            I => n3287
        );

    \I__6925\ : InMux
    port map (
            O => \N__36990\,
            I => n12935
        );

    \I__6924\ : CascadeMux
    port map (
            O => \N__36987\,
            I => \N__36983\
        );

    \I__6923\ : InMux
    port map (
            O => \N__36986\,
            I => \N__36980\
        );

    \I__6922\ : InMux
    port map (
            O => \N__36983\,
            I => \N__36977\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__36980\,
            I => \N__36973\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__36977\,
            I => \N__36970\
        );

    \I__6919\ : InMux
    port map (
            O => \N__36976\,
            I => \N__36967\
        );

    \I__6918\ : Span4Mux_s1_v
    port map (
            O => \N__36973\,
            I => \N__36960\
        );

    \I__6917\ : Span4Mux_h
    port map (
            O => \N__36970\,
            I => \N__36960\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__36967\,
            I => \N__36960\
        );

    \I__6915\ : Span4Mux_h
    port map (
            O => \N__36960\,
            I => \N__36957\
        );

    \I__6914\ : Odrv4
    port map (
            O => \N__36957\,
            I => n3219
        );

    \I__6913\ : CascadeMux
    port map (
            O => \N__36954\,
            I => \N__36951\
        );

    \I__6912\ : InMux
    port map (
            O => \N__36951\,
            I => \N__36948\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__36948\,
            I => \N__36945\
        );

    \I__6910\ : Span4Mux_s1_v
    port map (
            O => \N__36945\,
            I => \N__36942\
        );

    \I__6909\ : Odrv4
    port map (
            O => \N__36942\,
            I => n3286
        );

    \I__6908\ : InMux
    port map (
            O => \N__36939\,
            I => \bfn_7_31_0_\
        );

    \I__6907\ : CascadeMux
    port map (
            O => \N__36936\,
            I => \N__36933\
        );

    \I__6906\ : InMux
    port map (
            O => \N__36933\,
            I => \N__36929\
        );

    \I__6905\ : InMux
    port map (
            O => \N__36932\,
            I => \N__36926\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__36929\,
            I => \N__36923\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__36926\,
            I => n3218
        );

    \I__6902\ : Odrv4
    port map (
            O => \N__36923\,
            I => n3218
        );

    \I__6901\ : CascadeMux
    port map (
            O => \N__36918\,
            I => \N__36915\
        );

    \I__6900\ : InMux
    port map (
            O => \N__36915\,
            I => \N__36912\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__36912\,
            I => \N__36909\
        );

    \I__6898\ : Odrv4
    port map (
            O => \N__36909\,
            I => n3285
        );

    \I__6897\ : InMux
    port map (
            O => \N__36906\,
            I => n12937
        );

    \I__6896\ : CascadeMux
    port map (
            O => \N__36903\,
            I => \N__36900\
        );

    \I__6895\ : InMux
    port map (
            O => \N__36900\,
            I => \N__36896\
        );

    \I__6894\ : InMux
    port map (
            O => \N__36899\,
            I => \N__36892\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__36896\,
            I => \N__36889\
        );

    \I__6892\ : InMux
    port map (
            O => \N__36895\,
            I => \N__36886\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__36892\,
            I => n3232
        );

    \I__6890\ : Odrv4
    port map (
            O => \N__36889\,
            I => n3232
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__36886\,
            I => n3232
        );

    \I__6888\ : InMux
    port map (
            O => \N__36879\,
            I => \N__36876\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__36876\,
            I => n3299
        );

    \I__6886\ : InMux
    port map (
            O => \N__36873\,
            I => n12923
        );

    \I__6885\ : CascadeMux
    port map (
            O => \N__36870\,
            I => \N__36867\
        );

    \I__6884\ : InMux
    port map (
            O => \N__36867\,
            I => \N__36862\
        );

    \I__6883\ : InMux
    port map (
            O => \N__36866\,
            I => \N__36859\
        );

    \I__6882\ : InMux
    port map (
            O => \N__36865\,
            I => \N__36856\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__36862\,
            I => \N__36853\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__36859\,
            I => n3231
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__36856\,
            I => n3231
        );

    \I__6878\ : Odrv4
    port map (
            O => \N__36853\,
            I => n3231
        );

    \I__6877\ : InMux
    port map (
            O => \N__36846\,
            I => n12924
        );

    \I__6876\ : InMux
    port map (
            O => \N__36843\,
            I => \N__36840\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__36840\,
            I => n3298
        );

    \I__6874\ : CascadeMux
    port map (
            O => \N__36837\,
            I => \N__36834\
        );

    \I__6873\ : InMux
    port map (
            O => \N__36834\,
            I => \N__36829\
        );

    \I__6872\ : InMux
    port map (
            O => \N__36833\,
            I => \N__36826\
        );

    \I__6871\ : InMux
    port map (
            O => \N__36832\,
            I => \N__36823\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__36829\,
            I => \N__36820\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__36826\,
            I => n3230
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__36823\,
            I => n3230
        );

    \I__6867\ : Odrv4
    port map (
            O => \N__36820\,
            I => n3230
        );

    \I__6866\ : InMux
    port map (
            O => \N__36813\,
            I => \N__36810\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__36810\,
            I => \N__36807\
        );

    \I__6864\ : Odrv4
    port map (
            O => \N__36807\,
            I => n15079
        );

    \I__6863\ : InMux
    port map (
            O => \N__36804\,
            I => n12925
        );

    \I__6862\ : InMux
    port map (
            O => \N__36801\,
            I => \N__36797\
        );

    \I__6861\ : CascadeMux
    port map (
            O => \N__36800\,
            I => \N__36794\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__36797\,
            I => \N__36790\
        );

    \I__6859\ : InMux
    port map (
            O => \N__36794\,
            I => \N__36787\
        );

    \I__6858\ : InMux
    port map (
            O => \N__36793\,
            I => \N__36784\
        );

    \I__6857\ : Span4Mux_h
    port map (
            O => \N__36790\,
            I => \N__36779\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__36787\,
            I => \N__36779\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__36784\,
            I => n3229
        );

    \I__6854\ : Odrv4
    port map (
            O => \N__36779\,
            I => n3229
        );

    \I__6853\ : InMux
    port map (
            O => \N__36774\,
            I => \N__36771\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__36771\,
            I => \N__36768\
        );

    \I__6851\ : Span4Mux_s3_v
    port map (
            O => \N__36768\,
            I => \N__36765\
        );

    \I__6850\ : Odrv4
    port map (
            O => \N__36765\,
            I => n3296
        );

    \I__6849\ : InMux
    port map (
            O => \N__36762\,
            I => n12926
        );

    \I__6848\ : CascadeMux
    port map (
            O => \N__36759\,
            I => \N__36755\
        );

    \I__6847\ : InMux
    port map (
            O => \N__36758\,
            I => \N__36752\
        );

    \I__6846\ : InMux
    port map (
            O => \N__36755\,
            I => \N__36749\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__36752\,
            I => \N__36746\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__36749\,
            I => \N__36743\
        );

    \I__6843\ : Odrv4
    port map (
            O => \N__36746\,
            I => n3228
        );

    \I__6842\ : Odrv4
    port map (
            O => \N__36743\,
            I => n3228
        );

    \I__6841\ : InMux
    port map (
            O => \N__36738\,
            I => \N__36735\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__36735\,
            I => \N__36732\
        );

    \I__6839\ : Span4Mux_h
    port map (
            O => \N__36732\,
            I => \N__36729\
        );

    \I__6838\ : Odrv4
    port map (
            O => \N__36729\,
            I => n3295
        );

    \I__6837\ : InMux
    port map (
            O => \N__36726\,
            I => n12927
        );

    \I__6836\ : CascadeMux
    port map (
            O => \N__36723\,
            I => \N__36720\
        );

    \I__6835\ : InMux
    port map (
            O => \N__36720\,
            I => \N__36717\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__36717\,
            I => \N__36713\
        );

    \I__6833\ : InMux
    port map (
            O => \N__36716\,
            I => \N__36709\
        );

    \I__6832\ : Span4Mux_h
    port map (
            O => \N__36713\,
            I => \N__36706\
        );

    \I__6831\ : InMux
    port map (
            O => \N__36712\,
            I => \N__36703\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__36709\,
            I => n3227
        );

    \I__6829\ : Odrv4
    port map (
            O => \N__36706\,
            I => n3227
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__36703\,
            I => n3227
        );

    \I__6827\ : InMux
    port map (
            O => \N__36696\,
            I => \N__36693\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__36693\,
            I => \N__36690\
        );

    \I__6825\ : Span4Mux_s2_v
    port map (
            O => \N__36690\,
            I => \N__36687\
        );

    \I__6824\ : Odrv4
    port map (
            O => \N__36687\,
            I => n3294
        );

    \I__6823\ : InMux
    port map (
            O => \N__36684\,
            I => \bfn_7_30_0_\
        );

    \I__6822\ : CascadeMux
    port map (
            O => \N__36681\,
            I => \N__36678\
        );

    \I__6821\ : InMux
    port map (
            O => \N__36678\,
            I => \N__36674\
        );

    \I__6820\ : InMux
    port map (
            O => \N__36677\,
            I => \N__36671\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__36674\,
            I => \N__36668\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__36671\,
            I => n3226
        );

    \I__6817\ : Odrv12
    port map (
            O => \N__36668\,
            I => n3226
        );

    \I__6816\ : InMux
    port map (
            O => \N__36663\,
            I => \N__36660\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__36660\,
            I => \N__36657\
        );

    \I__6814\ : Odrv12
    port map (
            O => \N__36657\,
            I => n3293
        );

    \I__6813\ : InMux
    port map (
            O => \N__36654\,
            I => n12929
        );

    \I__6812\ : InMux
    port map (
            O => \N__36651\,
            I => n12974
        );

    \I__6811\ : CascadeMux
    port map (
            O => \N__36648\,
            I => \N__36645\
        );

    \I__6810\ : InMux
    port map (
            O => \N__36645\,
            I => \N__36642\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__36642\,
            I => \N__36638\
        );

    \I__6808\ : InMux
    port map (
            O => \N__36641\,
            I => \N__36635\
        );

    \I__6807\ : Span4Mux_v
    port map (
            O => \N__36638\,
            I => \N__36632\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__36635\,
            I => n12051
        );

    \I__6805\ : Odrv4
    port map (
            O => \N__36632\,
            I => n12051
        );

    \I__6804\ : InMux
    port map (
            O => \N__36627\,
            I => \N__36624\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__36624\,
            I => \N__36621\
        );

    \I__6802\ : Odrv4
    port map (
            O => \N__36621\,
            I => n15490
        );

    \I__6801\ : InMux
    port map (
            O => \N__36618\,
            I => \N__36614\
        );

    \I__6800\ : InMux
    port map (
            O => \N__36617\,
            I => \N__36611\
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__36614\,
            I => \N__36608\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__36611\,
            I => \N__36605\
        );

    \I__6797\ : Sp12to4
    port map (
            O => \N__36608\,
            I => \N__36602\
        );

    \I__6796\ : Span4Mux_v
    port map (
            O => \N__36605\,
            I => \N__36599\
        );

    \I__6795\ : Odrv12
    port map (
            O => \N__36602\,
            I => n319
        );

    \I__6794\ : Odrv4
    port map (
            O => \N__36599\,
            I => n319
        );

    \I__6793\ : InMux
    port map (
            O => \N__36594\,
            I => \N__36589\
        );

    \I__6792\ : InMux
    port map (
            O => \N__36593\,
            I => \N__36586\
        );

    \I__6791\ : InMux
    port map (
            O => \N__36592\,
            I => \N__36583\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__36589\,
            I => \N__36576\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__36586\,
            I => \N__36576\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__36583\,
            I => \N__36576\
        );

    \I__6787\ : Span4Mux_v
    port map (
            O => \N__36576\,
            I => \N__36573\
        );

    \I__6786\ : Odrv4
    port map (
            O => \N__36573\,
            I => n318
        );

    \I__6785\ : CascadeMux
    port map (
            O => \N__36570\,
            I => \N__36567\
        );

    \I__6784\ : InMux
    port map (
            O => \N__36567\,
            I => \N__36564\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__36564\,
            I => n3301
        );

    \I__6782\ : InMux
    port map (
            O => \N__36561\,
            I => n12921
        );

    \I__6781\ : CascadeMux
    port map (
            O => \N__36558\,
            I => \N__36554\
        );

    \I__6780\ : CascadeMux
    port map (
            O => \N__36557\,
            I => \N__36551\
        );

    \I__6779\ : InMux
    port map (
            O => \N__36554\,
            I => \N__36548\
        );

    \I__6778\ : InMux
    port map (
            O => \N__36551\,
            I => \N__36545\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__36548\,
            I => n3233
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__36545\,
            I => n3233
        );

    \I__6775\ : InMux
    port map (
            O => \N__36540\,
            I => \N__36537\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__36537\,
            I => n3300
        );

    \I__6773\ : InMux
    port map (
            O => \N__36534\,
            I => n12922
        );

    \I__6772\ : InMux
    port map (
            O => \N__36531\,
            I => n12965
        );

    \I__6771\ : InMux
    port map (
            O => \N__36528\,
            I => \N__36525\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__36525\,
            I => \N__36522\
        );

    \I__6769\ : Span4Mux_v
    port map (
            O => \N__36522\,
            I => \N__36519\
        );

    \I__6768\ : Odrv4
    port map (
            O => \N__36519\,
            I => n15652
        );

    \I__6767\ : InMux
    port map (
            O => \N__36516\,
            I => n12966
        );

    \I__6766\ : InMux
    port map (
            O => \N__36513\,
            I => \bfn_7_27_0_\
        );

    \I__6765\ : InMux
    port map (
            O => \N__36510\,
            I => n12968
        );

    \I__6764\ : InMux
    port map (
            O => \N__36507\,
            I => n12969
        );

    \I__6763\ : InMux
    port map (
            O => \N__36504\,
            I => n12970
        );

    \I__6762\ : InMux
    port map (
            O => \N__36501\,
            I => n12971
        );

    \I__6761\ : InMux
    port map (
            O => \N__36498\,
            I => n12972
        );

    \I__6760\ : InMux
    port map (
            O => \N__36495\,
            I => n12973
        );

    \I__6759\ : InMux
    port map (
            O => \N__36492\,
            I => \N__36488\
        );

    \I__6758\ : CascadeMux
    port map (
            O => \N__36491\,
            I => \N__36485\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__36488\,
            I => \N__36482\
        );

    \I__6756\ : InMux
    port map (
            O => \N__36485\,
            I => \N__36479\
        );

    \I__6755\ : Span4Mux_v
    port map (
            O => \N__36482\,
            I => \N__36476\
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__36479\,
            I => \N__36473\
        );

    \I__6753\ : Span4Mux_h
    port map (
            O => \N__36476\,
            I => \N__36468\
        );

    \I__6752\ : Span4Mux_s2_h
    port map (
            O => \N__36473\,
            I => \N__36468\
        );

    \I__6751\ : Odrv4
    port map (
            O => \N__36468\,
            I => n15322
        );

    \I__6750\ : InMux
    port map (
            O => \N__36465\,
            I => \N__36462\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__36462\,
            I => \N__36459\
        );

    \I__6748\ : Span4Mux_v
    port map (
            O => \N__36459\,
            I => \N__36450\
        );

    \I__6747\ : InMux
    port map (
            O => \N__36458\,
            I => \N__36447\
        );

    \I__6746\ : CascadeMux
    port map (
            O => \N__36457\,
            I => \N__36442\
        );

    \I__6745\ : CascadeMux
    port map (
            O => \N__36456\,
            I => \N__36439\
        );

    \I__6744\ : CascadeMux
    port map (
            O => \N__36455\,
            I => \N__36434\
        );

    \I__6743\ : CascadeMux
    port map (
            O => \N__36454\,
            I => \N__36431\
        );

    \I__6742\ : CascadeMux
    port map (
            O => \N__36453\,
            I => \N__36419\
        );

    \I__6741\ : Span4Mux_h
    port map (
            O => \N__36450\,
            I => \N__36412\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__36447\,
            I => \N__36412\
        );

    \I__6739\ : CascadeMux
    port map (
            O => \N__36446\,
            I => \N__36405\
        );

    \I__6738\ : CascadeMux
    port map (
            O => \N__36445\,
            I => \N__36402\
        );

    \I__6737\ : InMux
    port map (
            O => \N__36442\,
            I => \N__36393\
        );

    \I__6736\ : InMux
    port map (
            O => \N__36439\,
            I => \N__36393\
        );

    \I__6735\ : InMux
    port map (
            O => \N__36438\,
            I => \N__36393\
        );

    \I__6734\ : InMux
    port map (
            O => \N__36437\,
            I => \N__36393\
        );

    \I__6733\ : InMux
    port map (
            O => \N__36434\,
            I => \N__36380\
        );

    \I__6732\ : InMux
    port map (
            O => \N__36431\,
            I => \N__36380\
        );

    \I__6731\ : InMux
    port map (
            O => \N__36430\,
            I => \N__36380\
        );

    \I__6730\ : InMux
    port map (
            O => \N__36429\,
            I => \N__36380\
        );

    \I__6729\ : InMux
    port map (
            O => \N__36428\,
            I => \N__36380\
        );

    \I__6728\ : InMux
    port map (
            O => \N__36427\,
            I => \N__36380\
        );

    \I__6727\ : InMux
    port map (
            O => \N__36426\,
            I => \N__36375\
        );

    \I__6726\ : InMux
    port map (
            O => \N__36425\,
            I => \N__36375\
        );

    \I__6725\ : InMux
    port map (
            O => \N__36424\,
            I => \N__36370\
        );

    \I__6724\ : InMux
    port map (
            O => \N__36423\,
            I => \N__36370\
        );

    \I__6723\ : InMux
    port map (
            O => \N__36422\,
            I => \N__36363\
        );

    \I__6722\ : InMux
    port map (
            O => \N__36419\,
            I => \N__36363\
        );

    \I__6721\ : InMux
    port map (
            O => \N__36418\,
            I => \N__36363\
        );

    \I__6720\ : InMux
    port map (
            O => \N__36417\,
            I => \N__36360\
        );

    \I__6719\ : Span4Mux_v
    port map (
            O => \N__36412\,
            I => \N__36357\
        );

    \I__6718\ : InMux
    port map (
            O => \N__36411\,
            I => \N__36354\
        );

    \I__6717\ : InMux
    port map (
            O => \N__36410\,
            I => \N__36349\
        );

    \I__6716\ : InMux
    port map (
            O => \N__36409\,
            I => \N__36349\
        );

    \I__6715\ : InMux
    port map (
            O => \N__36408\,
            I => \N__36342\
        );

    \I__6714\ : InMux
    port map (
            O => \N__36405\,
            I => \N__36342\
        );

    \I__6713\ : InMux
    port map (
            O => \N__36402\,
            I => \N__36342\
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__36393\,
            I => \N__36335\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__36380\,
            I => \N__36335\
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__36375\,
            I => \N__36335\
        );

    \I__6709\ : LocalMux
    port map (
            O => \N__36370\,
            I => \N__36330\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__36363\,
            I => \N__36330\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__36360\,
            I => \N__36327\
        );

    \I__6706\ : Odrv4
    port map (
            O => \N__36357\,
            I => n2742
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__36354\,
            I => n2742
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__36349\,
            I => n2742
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__36342\,
            I => n2742
        );

    \I__6702\ : Odrv4
    port map (
            O => \N__36335\,
            I => n2742
        );

    \I__6701\ : Odrv4
    port map (
            O => \N__36330\,
            I => n2742
        );

    \I__6700\ : Odrv4
    port map (
            O => \N__36327\,
            I => n2742
        );

    \I__6699\ : InMux
    port map (
            O => \N__36312\,
            I => n12957
        );

    \I__6698\ : InMux
    port map (
            O => \N__36309\,
            I => \N__36306\
        );

    \I__6697\ : LocalMux
    port map (
            O => \N__36306\,
            I => \N__36303\
        );

    \I__6696\ : Span4Mux_h
    port map (
            O => \N__36303\,
            I => \N__36300\
        );

    \I__6695\ : Odrv4
    port map (
            O => \N__36300\,
            I => n15292
        );

    \I__6694\ : InMux
    port map (
            O => \N__36297\,
            I => \N__36289\
        );

    \I__6693\ : InMux
    port map (
            O => \N__36296\,
            I => \N__36286\
        );

    \I__6692\ : InMux
    port map (
            O => \N__36295\,
            I => \N__36283\
        );

    \I__6691\ : CascadeMux
    port map (
            O => \N__36294\,
            I => \N__36272\
        );

    \I__6690\ : CascadeMux
    port map (
            O => \N__36293\,
            I => \N__36269\
        );

    \I__6689\ : CascadeMux
    port map (
            O => \N__36292\,
            I => \N__36263\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__36289\,
            I => \N__36259\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__36286\,
            I => \N__36255\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__36283\,
            I => \N__36252\
        );

    \I__6685\ : CascadeMux
    port map (
            O => \N__36282\,
            I => \N__36249\
        );

    \I__6684\ : CascadeMux
    port map (
            O => \N__36281\,
            I => \N__36246\
        );

    \I__6683\ : CascadeMux
    port map (
            O => \N__36280\,
            I => \N__36242\
        );

    \I__6682\ : CascadeMux
    port map (
            O => \N__36279\,
            I => \N__36236\
        );

    \I__6681\ : CascadeMux
    port map (
            O => \N__36278\,
            I => \N__36231\
        );

    \I__6680\ : CascadeMux
    port map (
            O => \N__36277\,
            I => \N__36228\
        );

    \I__6679\ : CascadeMux
    port map (
            O => \N__36276\,
            I => \N__36225\
        );

    \I__6678\ : InMux
    port map (
            O => \N__36275\,
            I => \N__36217\
        );

    \I__6677\ : InMux
    port map (
            O => \N__36272\,
            I => \N__36217\
        );

    \I__6676\ : InMux
    port map (
            O => \N__36269\,
            I => \N__36217\
        );

    \I__6675\ : InMux
    port map (
            O => \N__36268\,
            I => \N__36212\
        );

    \I__6674\ : InMux
    port map (
            O => \N__36267\,
            I => \N__36212\
        );

    \I__6673\ : InMux
    port map (
            O => \N__36266\,
            I => \N__36205\
        );

    \I__6672\ : InMux
    port map (
            O => \N__36263\,
            I => \N__36205\
        );

    \I__6671\ : InMux
    port map (
            O => \N__36262\,
            I => \N__36205\
        );

    \I__6670\ : Span12Mux_s9_v
    port map (
            O => \N__36259\,
            I => \N__36202\
        );

    \I__6669\ : InMux
    port map (
            O => \N__36258\,
            I => \N__36199\
        );

    \I__6668\ : Span4Mux_h
    port map (
            O => \N__36255\,
            I => \N__36194\
        );

    \I__6667\ : Span4Mux_s3_h
    port map (
            O => \N__36252\,
            I => \N__36194\
        );

    \I__6666\ : InMux
    port map (
            O => \N__36249\,
            I => \N__36189\
        );

    \I__6665\ : InMux
    port map (
            O => \N__36246\,
            I => \N__36189\
        );

    \I__6664\ : InMux
    port map (
            O => \N__36245\,
            I => \N__36184\
        );

    \I__6663\ : InMux
    port map (
            O => \N__36242\,
            I => \N__36184\
        );

    \I__6662\ : InMux
    port map (
            O => \N__36241\,
            I => \N__36179\
        );

    \I__6661\ : InMux
    port map (
            O => \N__36240\,
            I => \N__36179\
        );

    \I__6660\ : InMux
    port map (
            O => \N__36239\,
            I => \N__36170\
        );

    \I__6659\ : InMux
    port map (
            O => \N__36236\,
            I => \N__36170\
        );

    \I__6658\ : InMux
    port map (
            O => \N__36235\,
            I => \N__36170\
        );

    \I__6657\ : InMux
    port map (
            O => \N__36234\,
            I => \N__36170\
        );

    \I__6656\ : InMux
    port map (
            O => \N__36231\,
            I => \N__36161\
        );

    \I__6655\ : InMux
    port map (
            O => \N__36228\,
            I => \N__36161\
        );

    \I__6654\ : InMux
    port map (
            O => \N__36225\,
            I => \N__36161\
        );

    \I__6653\ : InMux
    port map (
            O => \N__36224\,
            I => \N__36161\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__36217\,
            I => \N__36154\
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__36212\,
            I => \N__36154\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__36205\,
            I => \N__36154\
        );

    \I__6649\ : Odrv12
    port map (
            O => \N__36202\,
            I => n2643
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__36199\,
            I => n2643
        );

    \I__6647\ : Odrv4
    port map (
            O => \N__36194\,
            I => n2643
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__36189\,
            I => n2643
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__36184\,
            I => n2643
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__36179\,
            I => n2643
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__36170\,
            I => n2643
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__36161\,
            I => n2643
        );

    \I__6641\ : Odrv4
    port map (
            O => \N__36154\,
            I => n2643
        );

    \I__6640\ : InMux
    port map (
            O => \N__36135\,
            I => \N__36132\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__36132\,
            I => \N__36129\
        );

    \I__6638\ : Span4Mux_h
    port map (
            O => \N__36129\,
            I => \N__36126\
        );

    \I__6637\ : Odrv4
    port map (
            O => \N__36126\,
            I => encoder0_position_scaled_7
        );

    \I__6636\ : InMux
    port map (
            O => \N__36123\,
            I => n12958
        );

    \I__6635\ : InMux
    port map (
            O => \N__36120\,
            I => \N__36117\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__36117\,
            I => \N__36114\
        );

    \I__6633\ : Span4Mux_h
    port map (
            O => \N__36114\,
            I => \N__36110\
        );

    \I__6632\ : InMux
    port map (
            O => \N__36113\,
            I => \N__36107\
        );

    \I__6631\ : Odrv4
    port map (
            O => \N__36110\,
            I => n15830
        );

    \I__6630\ : LocalMux
    port map (
            O => \N__36107\,
            I => n15830
        );

    \I__6629\ : CascadeMux
    port map (
            O => \N__36102\,
            I => \N__36091\
        );

    \I__6628\ : InMux
    port map (
            O => \N__36101\,
            I => \N__36087\
        );

    \I__6627\ : CascadeMux
    port map (
            O => \N__36100\,
            I => \N__36082\
        );

    \I__6626\ : InMux
    port map (
            O => \N__36099\,
            I => \N__36077\
        );

    \I__6625\ : InMux
    port map (
            O => \N__36098\,
            I => \N__36077\
        );

    \I__6624\ : InMux
    port map (
            O => \N__36097\,
            I => \N__36074\
        );

    \I__6623\ : InMux
    port map (
            O => \N__36096\,
            I => \N__36071\
        );

    \I__6622\ : InMux
    port map (
            O => \N__36095\,
            I => \N__36065\
        );

    \I__6621\ : InMux
    port map (
            O => \N__36094\,
            I => \N__36058\
        );

    \I__6620\ : InMux
    port map (
            O => \N__36091\,
            I => \N__36058\
        );

    \I__6619\ : InMux
    port map (
            O => \N__36090\,
            I => \N__36058\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__36087\,
            I => \N__36054\
        );

    \I__6617\ : CascadeMux
    port map (
            O => \N__36086\,
            I => \N__36051\
        );

    \I__6616\ : CascadeMux
    port map (
            O => \N__36085\,
            I => \N__36045\
        );

    \I__6615\ : InMux
    port map (
            O => \N__36082\,
            I => \N__36041\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__36077\,
            I => \N__36038\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__36074\,
            I => \N__36035\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__36071\,
            I => \N__36032\
        );

    \I__6611\ : CascadeMux
    port map (
            O => \N__36070\,
            I => \N__36027\
        );

    \I__6610\ : CascadeMux
    port map (
            O => \N__36069\,
            I => \N__36024\
        );

    \I__6609\ : InMux
    port map (
            O => \N__36068\,
            I => \N__36020\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__36065\,
            I => \N__36015\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__36058\,
            I => \N__36015\
        );

    \I__6606\ : InMux
    port map (
            O => \N__36057\,
            I => \N__36012\
        );

    \I__6605\ : Span4Mux_v
    port map (
            O => \N__36054\,
            I => \N__36008\
        );

    \I__6604\ : InMux
    port map (
            O => \N__36051\,
            I => \N__35995\
        );

    \I__6603\ : InMux
    port map (
            O => \N__36050\,
            I => \N__35995\
        );

    \I__6602\ : InMux
    port map (
            O => \N__36049\,
            I => \N__35995\
        );

    \I__6601\ : InMux
    port map (
            O => \N__36048\,
            I => \N__35995\
        );

    \I__6600\ : InMux
    port map (
            O => \N__36045\,
            I => \N__35995\
        );

    \I__6599\ : InMux
    port map (
            O => \N__36044\,
            I => \N__35995\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__36041\,
            I => \N__35986\
        );

    \I__6597\ : Span4Mux_h
    port map (
            O => \N__36038\,
            I => \N__35986\
        );

    \I__6596\ : Span4Mux_v
    port map (
            O => \N__36035\,
            I => \N__35986\
        );

    \I__6595\ : Span4Mux_h
    port map (
            O => \N__36032\,
            I => \N__35986\
        );

    \I__6594\ : InMux
    port map (
            O => \N__36031\,
            I => \N__35975\
        );

    \I__6593\ : InMux
    port map (
            O => \N__36030\,
            I => \N__35975\
        );

    \I__6592\ : InMux
    port map (
            O => \N__36027\,
            I => \N__35975\
        );

    \I__6591\ : InMux
    port map (
            O => \N__36024\,
            I => \N__35975\
        );

    \I__6590\ : InMux
    port map (
            O => \N__36023\,
            I => \N__35975\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__36020\,
            I => \N__35968\
        );

    \I__6588\ : Span4Mux_h
    port map (
            O => \N__36015\,
            I => \N__35968\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__36012\,
            I => \N__35968\
        );

    \I__6586\ : InMux
    port map (
            O => \N__36011\,
            I => \N__35965\
        );

    \I__6585\ : Odrv4
    port map (
            O => \N__36008\,
            I => n2544
        );

    \I__6584\ : LocalMux
    port map (
            O => \N__35995\,
            I => n2544
        );

    \I__6583\ : Odrv4
    port map (
            O => \N__35986\,
            I => n2544
        );

    \I__6582\ : LocalMux
    port map (
            O => \N__35975\,
            I => n2544
        );

    \I__6581\ : Odrv4
    port map (
            O => \N__35968\,
            I => n2544
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__35965\,
            I => n2544
        );

    \I__6579\ : InMux
    port map (
            O => \N__35952\,
            I => \bfn_7_26_0_\
        );

    \I__6578\ : InMux
    port map (
            O => \N__35949\,
            I => \N__35945\
        );

    \I__6577\ : CascadeMux
    port map (
            O => \N__35948\,
            I => \N__35942\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__35945\,
            I => \N__35939\
        );

    \I__6575\ : InMux
    port map (
            O => \N__35942\,
            I => \N__35936\
        );

    \I__6574\ : Span4Mux_v
    port map (
            O => \N__35939\,
            I => \N__35933\
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__35936\,
            I => \N__35930\
        );

    \I__6572\ : Span4Mux_v
    port map (
            O => \N__35933\,
            I => \N__35927\
        );

    \I__6571\ : Span4Mux_v
    port map (
            O => \N__35930\,
            I => \N__35924\
        );

    \I__6570\ : Span4Mux_h
    port map (
            O => \N__35927\,
            I => \N__35921\
        );

    \I__6569\ : Span4Mux_h
    port map (
            O => \N__35924\,
            I => \N__35918\
        );

    \I__6568\ : Odrv4
    port map (
            O => \N__35921\,
            I => n15802
        );

    \I__6567\ : Odrv4
    port map (
            O => \N__35918\,
            I => n15802
        );

    \I__6566\ : InMux
    port map (
            O => \N__35913\,
            I => \N__35908\
        );

    \I__6565\ : CascadeMux
    port map (
            O => \N__35912\,
            I => \N__35905\
        );

    \I__6564\ : InMux
    port map (
            O => \N__35911\,
            I => \N__35893\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__35908\,
            I => \N__35890\
        );

    \I__6562\ : InMux
    port map (
            O => \N__35905\,
            I => \N__35881\
        );

    \I__6561\ : InMux
    port map (
            O => \N__35904\,
            I => \N__35881\
        );

    \I__6560\ : InMux
    port map (
            O => \N__35903\,
            I => \N__35881\
        );

    \I__6559\ : InMux
    port map (
            O => \N__35902\,
            I => \N__35881\
        );

    \I__6558\ : InMux
    port map (
            O => \N__35901\,
            I => \N__35878\
        );

    \I__6557\ : InMux
    port map (
            O => \N__35900\,
            I => \N__35875\
        );

    \I__6556\ : CascadeMux
    port map (
            O => \N__35899\,
            I => \N__35871\
        );

    \I__6555\ : CascadeMux
    port map (
            O => \N__35898\,
            I => \N__35863\
        );

    \I__6554\ : CascadeMux
    port map (
            O => \N__35897\,
            I => \N__35857\
        );

    \I__6553\ : InMux
    port map (
            O => \N__35896\,
            I => \N__35852\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__35893\,
            I => \N__35847\
        );

    \I__6551\ : Span4Mux_h
    port map (
            O => \N__35890\,
            I => \N__35847\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__35881\,
            I => \N__35844\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__35878\,
            I => \N__35839\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__35875\,
            I => \N__35839\
        );

    \I__6547\ : InMux
    port map (
            O => \N__35874\,
            I => \N__35832\
        );

    \I__6546\ : InMux
    port map (
            O => \N__35871\,
            I => \N__35832\
        );

    \I__6545\ : InMux
    port map (
            O => \N__35870\,
            I => \N__35832\
        );

    \I__6544\ : InMux
    port map (
            O => \N__35869\,
            I => \N__35829\
        );

    \I__6543\ : InMux
    port map (
            O => \N__35868\,
            I => \N__35822\
        );

    \I__6542\ : InMux
    port map (
            O => \N__35867\,
            I => \N__35822\
        );

    \I__6541\ : InMux
    port map (
            O => \N__35866\,
            I => \N__35822\
        );

    \I__6540\ : InMux
    port map (
            O => \N__35863\,
            I => \N__35813\
        );

    \I__6539\ : InMux
    port map (
            O => \N__35862\,
            I => \N__35813\
        );

    \I__6538\ : InMux
    port map (
            O => \N__35861\,
            I => \N__35813\
        );

    \I__6537\ : InMux
    port map (
            O => \N__35860\,
            I => \N__35813\
        );

    \I__6536\ : InMux
    port map (
            O => \N__35857\,
            I => \N__35806\
        );

    \I__6535\ : InMux
    port map (
            O => \N__35856\,
            I => \N__35806\
        );

    \I__6534\ : InMux
    port map (
            O => \N__35855\,
            I => \N__35806\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__35852\,
            I => \N__35801\
        );

    \I__6532\ : Span4Mux_v
    port map (
            O => \N__35847\,
            I => \N__35801\
        );

    \I__6531\ : Span4Mux_h
    port map (
            O => \N__35844\,
            I => \N__35796\
        );

    \I__6530\ : Span4Mux_v
    port map (
            O => \N__35839\,
            I => \N__35796\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__35832\,
            I => n2445
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__35829\,
            I => n2445
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__35822\,
            I => n2445
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__35813\,
            I => n2445
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__35806\,
            I => n2445
        );

    \I__6524\ : Odrv4
    port map (
            O => \N__35801\,
            I => n2445
        );

    \I__6523\ : Odrv4
    port map (
            O => \N__35796\,
            I => n2445
        );

    \I__6522\ : InMux
    port map (
            O => \N__35781\,
            I => n12960
        );

    \I__6521\ : InMux
    port map (
            O => \N__35778\,
            I => \N__35775\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__35775\,
            I => \N__35772\
        );

    \I__6519\ : Span4Mux_v
    port map (
            O => \N__35772\,
            I => \N__35769\
        );

    \I__6518\ : Span4Mux_h
    port map (
            O => \N__35769\,
            I => \N__35766\
        );

    \I__6517\ : Span4Mux_v
    port map (
            O => \N__35766\,
            I => \N__35762\
        );

    \I__6516\ : InMux
    port map (
            O => \N__35765\,
            I => \N__35759\
        );

    \I__6515\ : Odrv4
    port map (
            O => \N__35762\,
            I => n15775
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__35759\,
            I => n15775
        );

    \I__6513\ : InMux
    port map (
            O => \N__35754\,
            I => \N__35751\
        );

    \I__6512\ : LocalMux
    port map (
            O => \N__35751\,
            I => \N__35748\
        );

    \I__6511\ : Span4Mux_h
    port map (
            O => \N__35748\,
            I => \N__35735\
        );

    \I__6510\ : InMux
    port map (
            O => \N__35747\,
            I => \N__35730\
        );

    \I__6509\ : InMux
    port map (
            O => \N__35746\,
            I => \N__35730\
        );

    \I__6508\ : CascadeMux
    port map (
            O => \N__35745\,
            I => \N__35727\
        );

    \I__6507\ : InMux
    port map (
            O => \N__35744\,
            I => \N__35724\
        );

    \I__6506\ : CascadeMux
    port map (
            O => \N__35743\,
            I => \N__35719\
        );

    \I__6505\ : CascadeMux
    port map (
            O => \N__35742\,
            I => \N__35713\
        );

    \I__6504\ : CascadeMux
    port map (
            O => \N__35741\,
            I => \N__35710\
        );

    \I__6503\ : CascadeMux
    port map (
            O => \N__35740\,
            I => \N__35705\
        );

    \I__6502\ : CascadeMux
    port map (
            O => \N__35739\,
            I => \N__35699\
        );

    \I__6501\ : CascadeMux
    port map (
            O => \N__35738\,
            I => \N__35696\
        );

    \I__6500\ : Span4Mux_v
    port map (
            O => \N__35735\,
            I => \N__35690\
        );

    \I__6499\ : LocalMux
    port map (
            O => \N__35730\,
            I => \N__35690\
        );

    \I__6498\ : InMux
    port map (
            O => \N__35727\,
            I => \N__35687\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__35724\,
            I => \N__35684\
        );

    \I__6496\ : InMux
    port map (
            O => \N__35723\,
            I => \N__35675\
        );

    \I__6495\ : InMux
    port map (
            O => \N__35722\,
            I => \N__35675\
        );

    \I__6494\ : InMux
    port map (
            O => \N__35719\,
            I => \N__35675\
        );

    \I__6493\ : InMux
    port map (
            O => \N__35718\,
            I => \N__35675\
        );

    \I__6492\ : InMux
    port map (
            O => \N__35717\,
            I => \N__35670\
        );

    \I__6491\ : InMux
    port map (
            O => \N__35716\,
            I => \N__35670\
        );

    \I__6490\ : InMux
    port map (
            O => \N__35713\,
            I => \N__35663\
        );

    \I__6489\ : InMux
    port map (
            O => \N__35710\,
            I => \N__35663\
        );

    \I__6488\ : InMux
    port map (
            O => \N__35709\,
            I => \N__35663\
        );

    \I__6487\ : InMux
    port map (
            O => \N__35708\,
            I => \N__35656\
        );

    \I__6486\ : InMux
    port map (
            O => \N__35705\,
            I => \N__35656\
        );

    \I__6485\ : InMux
    port map (
            O => \N__35704\,
            I => \N__35656\
        );

    \I__6484\ : InMux
    port map (
            O => \N__35703\,
            I => \N__35645\
        );

    \I__6483\ : InMux
    port map (
            O => \N__35702\,
            I => \N__35645\
        );

    \I__6482\ : InMux
    port map (
            O => \N__35699\,
            I => \N__35645\
        );

    \I__6481\ : InMux
    port map (
            O => \N__35696\,
            I => \N__35645\
        );

    \I__6480\ : InMux
    port map (
            O => \N__35695\,
            I => \N__35645\
        );

    \I__6479\ : Odrv4
    port map (
            O => \N__35690\,
            I => n2346
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__35687\,
            I => n2346
        );

    \I__6477\ : Odrv4
    port map (
            O => \N__35684\,
            I => n2346
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__35675\,
            I => n2346
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__35670\,
            I => n2346
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__35663\,
            I => n2346
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__35656\,
            I => n2346
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__35645\,
            I => n2346
        );

    \I__6471\ : InMux
    port map (
            O => \N__35628\,
            I => n12961
        );

    \I__6470\ : InMux
    port map (
            O => \N__35625\,
            I => \N__35622\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__35622\,
            I => \N__35619\
        );

    \I__6468\ : Span4Mux_v
    port map (
            O => \N__35619\,
            I => \N__35616\
        );

    \I__6467\ : Span4Mux_v
    port map (
            O => \N__35616\,
            I => \N__35613\
        );

    \I__6466\ : Span4Mux_h
    port map (
            O => \N__35613\,
            I => \N__35609\
        );

    \I__6465\ : InMux
    port map (
            O => \N__35612\,
            I => \N__35606\
        );

    \I__6464\ : Odrv4
    port map (
            O => \N__35609\,
            I => n15748
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__35606\,
            I => n15748
        );

    \I__6462\ : InMux
    port map (
            O => \N__35601\,
            I => \N__35598\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__35598\,
            I => \N__35591\
        );

    \I__6460\ : InMux
    port map (
            O => \N__35597\,
            I => \N__35584\
        );

    \I__6459\ : CascadeMux
    port map (
            O => \N__35596\,
            I => \N__35581\
        );

    \I__6458\ : CascadeMux
    port map (
            O => \N__35595\,
            I => \N__35578\
        );

    \I__6457\ : CascadeMux
    port map (
            O => \N__35594\,
            I => \N__35575\
        );

    \I__6456\ : Span4Mux_v
    port map (
            O => \N__35591\,
            I => \N__35570\
        );

    \I__6455\ : CascadeMux
    port map (
            O => \N__35590\,
            I => \N__35567\
        );

    \I__6454\ : CascadeMux
    port map (
            O => \N__35589\,
            I => \N__35563\
        );

    \I__6453\ : CascadeMux
    port map (
            O => \N__35588\,
            I => \N__35558\
        );

    \I__6452\ : CascadeMux
    port map (
            O => \N__35587\,
            I => \N__35555\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__35584\,
            I => \N__35551\
        );

    \I__6450\ : InMux
    port map (
            O => \N__35581\,
            I => \N__35542\
        );

    \I__6449\ : InMux
    port map (
            O => \N__35578\,
            I => \N__35542\
        );

    \I__6448\ : InMux
    port map (
            O => \N__35575\,
            I => \N__35542\
        );

    \I__6447\ : InMux
    port map (
            O => \N__35574\,
            I => \N__35542\
        );

    \I__6446\ : CascadeMux
    port map (
            O => \N__35573\,
            I => \N__35534\
        );

    \I__6445\ : Span4Mux_h
    port map (
            O => \N__35570\,
            I => \N__35530\
        );

    \I__6444\ : InMux
    port map (
            O => \N__35567\,
            I => \N__35525\
        );

    \I__6443\ : InMux
    port map (
            O => \N__35566\,
            I => \N__35525\
        );

    \I__6442\ : InMux
    port map (
            O => \N__35563\,
            I => \N__35518\
        );

    \I__6441\ : InMux
    port map (
            O => \N__35562\,
            I => \N__35518\
        );

    \I__6440\ : InMux
    port map (
            O => \N__35561\,
            I => \N__35518\
        );

    \I__6439\ : InMux
    port map (
            O => \N__35558\,
            I => \N__35511\
        );

    \I__6438\ : InMux
    port map (
            O => \N__35555\,
            I => \N__35511\
        );

    \I__6437\ : InMux
    port map (
            O => \N__35554\,
            I => \N__35511\
        );

    \I__6436\ : Span4Mux_h
    port map (
            O => \N__35551\,
            I => \N__35506\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__35542\,
            I => \N__35506\
        );

    \I__6434\ : InMux
    port map (
            O => \N__35541\,
            I => \N__35501\
        );

    \I__6433\ : InMux
    port map (
            O => \N__35540\,
            I => \N__35501\
        );

    \I__6432\ : InMux
    port map (
            O => \N__35539\,
            I => \N__35490\
        );

    \I__6431\ : InMux
    port map (
            O => \N__35538\,
            I => \N__35490\
        );

    \I__6430\ : InMux
    port map (
            O => \N__35537\,
            I => \N__35490\
        );

    \I__6429\ : InMux
    port map (
            O => \N__35534\,
            I => \N__35490\
        );

    \I__6428\ : InMux
    port map (
            O => \N__35533\,
            I => \N__35490\
        );

    \I__6427\ : Odrv4
    port map (
            O => \N__35530\,
            I => n2247
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__35525\,
            I => n2247
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__35518\,
            I => n2247
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__35511\,
            I => n2247
        );

    \I__6423\ : Odrv4
    port map (
            O => \N__35506\,
            I => n2247
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__35501\,
            I => n2247
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__35490\,
            I => n2247
        );

    \I__6420\ : InMux
    port map (
            O => \N__35475\,
            I => n12962
        );

    \I__6419\ : InMux
    port map (
            O => \N__35472\,
            I => \N__35469\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__35469\,
            I => \N__35466\
        );

    \I__6417\ : Span4Mux_h
    port map (
            O => \N__35466\,
            I => \N__35463\
        );

    \I__6416\ : Span4Mux_v
    port map (
            O => \N__35463\,
            I => \N__35459\
        );

    \I__6415\ : InMux
    port map (
            O => \N__35462\,
            I => \N__35456\
        );

    \I__6414\ : Odrv4
    port map (
            O => \N__35459\,
            I => n15722
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__35456\,
            I => n15722
        );

    \I__6412\ : InMux
    port map (
            O => \N__35451\,
            I => \N__35448\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__35448\,
            I => \N__35438\
        );

    \I__6410\ : InMux
    port map (
            O => \N__35447\,
            I => \N__35433\
        );

    \I__6409\ : CascadeMux
    port map (
            O => \N__35446\,
            I => \N__35430\
        );

    \I__6408\ : CascadeMux
    port map (
            O => \N__35445\,
            I => \N__35427\
        );

    \I__6407\ : CascadeMux
    port map (
            O => \N__35444\,
            I => \N__35424\
        );

    \I__6406\ : CascadeMux
    port map (
            O => \N__35443\,
            I => \N__35421\
        );

    \I__6405\ : CascadeMux
    port map (
            O => \N__35442\,
            I => \N__35413\
        );

    \I__6404\ : CascadeMux
    port map (
            O => \N__35441\,
            I => \N__35410\
        );

    \I__6403\ : Span4Mux_v
    port map (
            O => \N__35438\,
            I => \N__35405\
        );

    \I__6402\ : InMux
    port map (
            O => \N__35437\,
            I => \N__35400\
        );

    \I__6401\ : InMux
    port map (
            O => \N__35436\,
            I => \N__35400\
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__35433\,
            I => \N__35396\
        );

    \I__6399\ : InMux
    port map (
            O => \N__35430\,
            I => \N__35391\
        );

    \I__6398\ : InMux
    port map (
            O => \N__35427\,
            I => \N__35391\
        );

    \I__6397\ : InMux
    port map (
            O => \N__35424\,
            I => \N__35380\
        );

    \I__6396\ : InMux
    port map (
            O => \N__35421\,
            I => \N__35380\
        );

    \I__6395\ : InMux
    port map (
            O => \N__35420\,
            I => \N__35380\
        );

    \I__6394\ : InMux
    port map (
            O => \N__35419\,
            I => \N__35380\
        );

    \I__6393\ : InMux
    port map (
            O => \N__35418\,
            I => \N__35380\
        );

    \I__6392\ : InMux
    port map (
            O => \N__35417\,
            I => \N__35373\
        );

    \I__6391\ : InMux
    port map (
            O => \N__35416\,
            I => \N__35373\
        );

    \I__6390\ : InMux
    port map (
            O => \N__35413\,
            I => \N__35364\
        );

    \I__6389\ : InMux
    port map (
            O => \N__35410\,
            I => \N__35364\
        );

    \I__6388\ : InMux
    port map (
            O => \N__35409\,
            I => \N__35364\
        );

    \I__6387\ : InMux
    port map (
            O => \N__35408\,
            I => \N__35364\
        );

    \I__6386\ : Span4Mux_v
    port map (
            O => \N__35405\,
            I => \N__35359\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__35400\,
            I => \N__35359\
        );

    \I__6384\ : InMux
    port map (
            O => \N__35399\,
            I => \N__35356\
        );

    \I__6383\ : Span4Mux_h
    port map (
            O => \N__35396\,
            I => \N__35353\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__35391\,
            I => \N__35348\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__35380\,
            I => \N__35348\
        );

    \I__6380\ : InMux
    port map (
            O => \N__35379\,
            I => \N__35343\
        );

    \I__6379\ : InMux
    port map (
            O => \N__35378\,
            I => \N__35343\
        );

    \I__6378\ : LocalMux
    port map (
            O => \N__35373\,
            I => n2148
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__35364\,
            I => n2148
        );

    \I__6376\ : Odrv4
    port map (
            O => \N__35359\,
            I => n2148
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__35356\,
            I => n2148
        );

    \I__6374\ : Odrv4
    port map (
            O => \N__35353\,
            I => n2148
        );

    \I__6373\ : Odrv4
    port map (
            O => \N__35348\,
            I => n2148
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__35343\,
            I => n2148
        );

    \I__6371\ : InMux
    port map (
            O => \N__35328\,
            I => n12963
        );

    \I__6370\ : InMux
    port map (
            O => \N__35325\,
            I => \N__35322\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__35322\,
            I => \N__35319\
        );

    \I__6368\ : Span4Mux_h
    port map (
            O => \N__35319\,
            I => \N__35316\
        );

    \I__6367\ : Span4Mux_v
    port map (
            O => \N__35316\,
            I => \N__35312\
        );

    \I__6366\ : InMux
    port map (
            O => \N__35315\,
            I => \N__35309\
        );

    \I__6365\ : Odrv4
    port map (
            O => \N__35312\,
            I => n15697
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__35309\,
            I => n15697
        );

    \I__6363\ : InMux
    port map (
            O => \N__35304\,
            I => \N__35299\
        );

    \I__6362\ : CascadeMux
    port map (
            O => \N__35303\,
            I => \N__35293\
        );

    \I__6361\ : CascadeMux
    port map (
            O => \N__35302\,
            I => \N__35289\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__35299\,
            I => \N__35285\
        );

    \I__6359\ : InMux
    port map (
            O => \N__35298\,
            I => \N__35282\
        );

    \I__6358\ : InMux
    port map (
            O => \N__35297\,
            I => \N__35271\
        );

    \I__6357\ : InMux
    port map (
            O => \N__35296\,
            I => \N__35271\
        );

    \I__6356\ : InMux
    port map (
            O => \N__35293\,
            I => \N__35266\
        );

    \I__6355\ : InMux
    port map (
            O => \N__35292\,
            I => \N__35266\
        );

    \I__6354\ : InMux
    port map (
            O => \N__35289\,
            I => \N__35263\
        );

    \I__6353\ : CascadeMux
    port map (
            O => \N__35288\,
            I => \N__35259\
        );

    \I__6352\ : Span4Mux_v
    port map (
            O => \N__35285\,
            I => \N__35254\
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__35282\,
            I => \N__35251\
        );

    \I__6350\ : CascadeMux
    port map (
            O => \N__35281\,
            I => \N__35248\
        );

    \I__6349\ : CascadeMux
    port map (
            O => \N__35280\,
            I => \N__35245\
        );

    \I__6348\ : InMux
    port map (
            O => \N__35279\,
            I => \N__35240\
        );

    \I__6347\ : InMux
    port map (
            O => \N__35278\,
            I => \N__35233\
        );

    \I__6346\ : InMux
    port map (
            O => \N__35277\,
            I => \N__35233\
        );

    \I__6345\ : InMux
    port map (
            O => \N__35276\,
            I => \N__35233\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__35271\,
            I => \N__35230\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__35266\,
            I => \N__35225\
        );

    \I__6342\ : LocalMux
    port map (
            O => \N__35263\,
            I => \N__35225\
        );

    \I__6341\ : InMux
    port map (
            O => \N__35262\,
            I => \N__35218\
        );

    \I__6340\ : InMux
    port map (
            O => \N__35259\,
            I => \N__35218\
        );

    \I__6339\ : InMux
    port map (
            O => \N__35258\,
            I => \N__35218\
        );

    \I__6338\ : InMux
    port map (
            O => \N__35257\,
            I => \N__35215\
        );

    \I__6337\ : Span4Mux_v
    port map (
            O => \N__35254\,
            I => \N__35210\
        );

    \I__6336\ : Span4Mux_v
    port map (
            O => \N__35251\,
            I => \N__35210\
        );

    \I__6335\ : InMux
    port map (
            O => \N__35248\,
            I => \N__35203\
        );

    \I__6334\ : InMux
    port map (
            O => \N__35245\,
            I => \N__35203\
        );

    \I__6333\ : InMux
    port map (
            O => \N__35244\,
            I => \N__35203\
        );

    \I__6332\ : InMux
    port map (
            O => \N__35243\,
            I => \N__35200\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__35240\,
            I => n2049
        );

    \I__6330\ : LocalMux
    port map (
            O => \N__35233\,
            I => n2049
        );

    \I__6329\ : Odrv4
    port map (
            O => \N__35230\,
            I => n2049
        );

    \I__6328\ : Odrv4
    port map (
            O => \N__35225\,
            I => n2049
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__35218\,
            I => n2049
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__35215\,
            I => n2049
        );

    \I__6325\ : Odrv4
    port map (
            O => \N__35210\,
            I => n2049
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__35203\,
            I => n2049
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__35200\,
            I => n2049
        );

    \I__6322\ : InMux
    port map (
            O => \N__35181\,
            I => n12964
        );

    \I__6321\ : InMux
    port map (
            O => \N__35178\,
            I => \N__35173\
        );

    \I__6320\ : InMux
    port map (
            O => \N__35177\,
            I => \N__35170\
        );

    \I__6319\ : InMux
    port map (
            O => \N__35176\,
            I => \N__35167\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__35173\,
            I => \N__35164\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__35170\,
            I => \N__35161\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__35167\,
            I => \N__35158\
        );

    \I__6315\ : Span4Mux_v
    port map (
            O => \N__35164\,
            I => \N__35153\
        );

    \I__6314\ : Span4Mux_v
    port map (
            O => \N__35161\,
            I => \N__35153\
        );

    \I__6313\ : Span4Mux_v
    port map (
            O => \N__35158\,
            I => \N__35148\
        );

    \I__6312\ : Span4Mux_h
    port map (
            O => \N__35153\,
            I => \N__35148\
        );

    \I__6311\ : Odrv4
    port map (
            O => \N__35148\,
            I => n315
        );

    \I__6310\ : InMux
    port map (
            O => \N__35145\,
            I => \N__35142\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__35142\,
            I => \N__35138\
        );

    \I__6308\ : InMux
    port map (
            O => \N__35141\,
            I => \N__35134\
        );

    \I__6307\ : Span4Mux_h
    port map (
            O => \N__35138\,
            I => \N__35131\
        );

    \I__6306\ : InMux
    port map (
            O => \N__35137\,
            I => \N__35128\
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__35134\,
            I => \N__35125\
        );

    \I__6304\ : Odrv4
    port map (
            O => \N__35131\,
            I => n311
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__35128\,
            I => n311
        );

    \I__6302\ : Odrv4
    port map (
            O => \N__35125\,
            I => n311
        );

    \I__6301\ : InMux
    port map (
            O => \N__35118\,
            I => \bfn_7_25_0_\
        );

    \I__6300\ : InMux
    port map (
            O => \N__35115\,
            I => \N__35112\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__35112\,
            I => \N__35109\
        );

    \I__6298\ : Span4Mux_h
    port map (
            O => \N__35109\,
            I => \N__35106\
        );

    \I__6297\ : Odrv4
    port map (
            O => \N__35106\,
            I => n15485
        );

    \I__6296\ : InMux
    port map (
            O => \N__35103\,
            I => \N__35100\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__35100\,
            I => \N__35096\
        );

    \I__6294\ : InMux
    port map (
            O => \N__35099\,
            I => \N__35084\
        );

    \I__6293\ : Span4Mux_v
    port map (
            O => \N__35096\,
            I => \N__35081\
        );

    \I__6292\ : CascadeMux
    port map (
            O => \N__35095\,
            I => \N__35073\
        );

    \I__6291\ : CascadeMux
    port map (
            O => \N__35094\,
            I => \N__35069\
        );

    \I__6290\ : CascadeMux
    port map (
            O => \N__35093\,
            I => \N__35063\
        );

    \I__6289\ : InMux
    port map (
            O => \N__35092\,
            I => \N__35058\
        );

    \I__6288\ : InMux
    port map (
            O => \N__35091\,
            I => \N__35058\
        );

    \I__6287\ : CascadeMux
    port map (
            O => \N__35090\,
            I => \N__35054\
        );

    \I__6286\ : CascadeMux
    port map (
            O => \N__35089\,
            I => \N__35051\
        );

    \I__6285\ : CascadeMux
    port map (
            O => \N__35088\,
            I => \N__35046\
        );

    \I__6284\ : CascadeMux
    port map (
            O => \N__35087\,
            I => \N__35042\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__35084\,
            I => \N__35032\
        );

    \I__6282\ : Span4Mux_v
    port map (
            O => \N__35081\,
            I => \N__35029\
        );

    \I__6281\ : InMux
    port map (
            O => \N__35080\,
            I => \N__35016\
        );

    \I__6280\ : InMux
    port map (
            O => \N__35079\,
            I => \N__35016\
        );

    \I__6279\ : InMux
    port map (
            O => \N__35078\,
            I => \N__35016\
        );

    \I__6278\ : InMux
    port map (
            O => \N__35077\,
            I => \N__35016\
        );

    \I__6277\ : InMux
    port map (
            O => \N__35076\,
            I => \N__35016\
        );

    \I__6276\ : InMux
    port map (
            O => \N__35073\,
            I => \N__35016\
        );

    \I__6275\ : InMux
    port map (
            O => \N__35072\,
            I => \N__35003\
        );

    \I__6274\ : InMux
    port map (
            O => \N__35069\,
            I => \N__35003\
        );

    \I__6273\ : InMux
    port map (
            O => \N__35068\,
            I => \N__35003\
        );

    \I__6272\ : InMux
    port map (
            O => \N__35067\,
            I => \N__35003\
        );

    \I__6271\ : InMux
    port map (
            O => \N__35066\,
            I => \N__35003\
        );

    \I__6270\ : InMux
    port map (
            O => \N__35063\,
            I => \N__35003\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__35058\,
            I => \N__35000\
        );

    \I__6268\ : InMux
    port map (
            O => \N__35057\,
            I => \N__34987\
        );

    \I__6267\ : InMux
    port map (
            O => \N__35054\,
            I => \N__34987\
        );

    \I__6266\ : InMux
    port map (
            O => \N__35051\,
            I => \N__34987\
        );

    \I__6265\ : InMux
    port map (
            O => \N__35050\,
            I => \N__34987\
        );

    \I__6264\ : InMux
    port map (
            O => \N__35049\,
            I => \N__34987\
        );

    \I__6263\ : InMux
    port map (
            O => \N__35046\,
            I => \N__34987\
        );

    \I__6262\ : InMux
    port map (
            O => \N__35045\,
            I => \N__34980\
        );

    \I__6261\ : InMux
    port map (
            O => \N__35042\,
            I => \N__34980\
        );

    \I__6260\ : InMux
    port map (
            O => \N__35041\,
            I => \N__34980\
        );

    \I__6259\ : InMux
    port map (
            O => \N__35040\,
            I => \N__34967\
        );

    \I__6258\ : InMux
    port map (
            O => \N__35039\,
            I => \N__34967\
        );

    \I__6257\ : InMux
    port map (
            O => \N__35038\,
            I => \N__34967\
        );

    \I__6256\ : InMux
    port map (
            O => \N__35037\,
            I => \N__34967\
        );

    \I__6255\ : InMux
    port map (
            O => \N__35036\,
            I => \N__34967\
        );

    \I__6254\ : InMux
    port map (
            O => \N__35035\,
            I => \N__34967\
        );

    \I__6253\ : Odrv4
    port map (
            O => \N__35032\,
            I => n3237
        );

    \I__6252\ : Odrv4
    port map (
            O => \N__35029\,
            I => n3237
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__35016\,
            I => n3237
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__35003\,
            I => n3237
        );

    \I__6249\ : Odrv4
    port map (
            O => \N__35000\,
            I => n3237
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__34987\,
            I => n3237
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__34980\,
            I => n3237
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__34967\,
            I => n3237
        );

    \I__6245\ : InMux
    port map (
            O => \N__34950\,
            I => n12952
        );

    \I__6244\ : InMux
    port map (
            O => \N__34947\,
            I => \N__34944\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__34944\,
            I => \N__34941\
        );

    \I__6242\ : Span4Mux_v
    port map (
            O => \N__34941\,
            I => \N__34937\
        );

    \I__6241\ : CascadeMux
    port map (
            O => \N__34940\,
            I => \N__34934\
        );

    \I__6240\ : Span4Mux_h
    port map (
            O => \N__34937\,
            I => \N__34931\
        );

    \I__6239\ : InMux
    port map (
            O => \N__34934\,
            I => \N__34928\
        );

    \I__6238\ : Odrv4
    port map (
            O => \N__34931\,
            I => n15451
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__34928\,
            I => n15451
        );

    \I__6236\ : CascadeMux
    port map (
            O => \N__34923\,
            I => \N__34919\
        );

    \I__6235\ : InMux
    port map (
            O => \N__34922\,
            I => \N__34912\
        );

    \I__6234\ : InMux
    port map (
            O => \N__34919\,
            I => \N__34901\
        );

    \I__6233\ : InMux
    port map (
            O => \N__34918\,
            I => \N__34901\
        );

    \I__6232\ : InMux
    port map (
            O => \N__34917\,
            I => \N__34898\
        );

    \I__6231\ : CascadeMux
    port map (
            O => \N__34916\,
            I => \N__34895\
        );

    \I__6230\ : CascadeMux
    port map (
            O => \N__34915\,
            I => \N__34892\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__34912\,
            I => \N__34885\
        );

    \I__6228\ : InMux
    port map (
            O => \N__34911\,
            I => \N__34882\
        );

    \I__6227\ : CascadeMux
    port map (
            O => \N__34910\,
            I => \N__34877\
        );

    \I__6226\ : CascadeMux
    port map (
            O => \N__34909\,
            I => \N__34871\
        );

    \I__6225\ : CascadeMux
    port map (
            O => \N__34908\,
            I => \N__34867\
        );

    \I__6224\ : CascadeMux
    port map (
            O => \N__34907\,
            I => \N__34863\
        );

    \I__6223\ : CascadeMux
    port map (
            O => \N__34906\,
            I => \N__34859\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__34901\,
            I => \N__34855\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__34898\,
            I => \N__34852\
        );

    \I__6220\ : InMux
    port map (
            O => \N__34895\,
            I => \N__34843\
        );

    \I__6219\ : InMux
    port map (
            O => \N__34892\,
            I => \N__34843\
        );

    \I__6218\ : InMux
    port map (
            O => \N__34891\,
            I => \N__34843\
        );

    \I__6217\ : InMux
    port map (
            O => \N__34890\,
            I => \N__34843\
        );

    \I__6216\ : InMux
    port map (
            O => \N__34889\,
            I => \N__34840\
        );

    \I__6215\ : CascadeMux
    port map (
            O => \N__34888\,
            I => \N__34836\
        );

    \I__6214\ : Span4Mux_h
    port map (
            O => \N__34885\,
            I => \N__34832\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__34882\,
            I => \N__34829\
        );

    \I__6212\ : CascadeMux
    port map (
            O => \N__34881\,
            I => \N__34826\
        );

    \I__6211\ : InMux
    port map (
            O => \N__34880\,
            I => \N__34814\
        );

    \I__6210\ : InMux
    port map (
            O => \N__34877\,
            I => \N__34814\
        );

    \I__6209\ : InMux
    port map (
            O => \N__34876\,
            I => \N__34814\
        );

    \I__6208\ : InMux
    port map (
            O => \N__34875\,
            I => \N__34814\
        );

    \I__6207\ : InMux
    port map (
            O => \N__34874\,
            I => \N__34807\
        );

    \I__6206\ : InMux
    port map (
            O => \N__34871\,
            I => \N__34807\
        );

    \I__6205\ : InMux
    port map (
            O => \N__34870\,
            I => \N__34807\
        );

    \I__6204\ : InMux
    port map (
            O => \N__34867\,
            I => \N__34802\
        );

    \I__6203\ : InMux
    port map (
            O => \N__34866\,
            I => \N__34802\
        );

    \I__6202\ : InMux
    port map (
            O => \N__34863\,
            I => \N__34793\
        );

    \I__6201\ : InMux
    port map (
            O => \N__34862\,
            I => \N__34793\
        );

    \I__6200\ : InMux
    port map (
            O => \N__34859\,
            I => \N__34793\
        );

    \I__6199\ : InMux
    port map (
            O => \N__34858\,
            I => \N__34793\
        );

    \I__6198\ : Span4Mux_v
    port map (
            O => \N__34855\,
            I => \N__34790\
        );

    \I__6197\ : Span4Mux_h
    port map (
            O => \N__34852\,
            I => \N__34783\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__34843\,
            I => \N__34783\
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__34840\,
            I => \N__34783\
        );

    \I__6194\ : InMux
    port map (
            O => \N__34839\,
            I => \N__34776\
        );

    \I__6193\ : InMux
    port map (
            O => \N__34836\,
            I => \N__34776\
        );

    \I__6192\ : InMux
    port map (
            O => \N__34835\,
            I => \N__34776\
        );

    \I__6191\ : Span4Mux_v
    port map (
            O => \N__34832\,
            I => \N__34771\
        );

    \I__6190\ : Span4Mux_s3_h
    port map (
            O => \N__34829\,
            I => \N__34771\
        );

    \I__6189\ : InMux
    port map (
            O => \N__34826\,
            I => \N__34762\
        );

    \I__6188\ : InMux
    port map (
            O => \N__34825\,
            I => \N__34762\
        );

    \I__6187\ : InMux
    port map (
            O => \N__34824\,
            I => \N__34762\
        );

    \I__6186\ : InMux
    port map (
            O => \N__34823\,
            I => \N__34762\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__34814\,
            I => n3138
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__34807\,
            I => n3138
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__34802\,
            I => n3138
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__34793\,
            I => n3138
        );

    \I__6181\ : Odrv4
    port map (
            O => \N__34790\,
            I => n3138
        );

    \I__6180\ : Odrv4
    port map (
            O => \N__34783\,
            I => n3138
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__34776\,
            I => n3138
        );

    \I__6178\ : Odrv4
    port map (
            O => \N__34771\,
            I => n3138
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__34762\,
            I => n3138
        );

    \I__6176\ : InMux
    port map (
            O => \N__34743\,
            I => n12953
        );

    \I__6175\ : InMux
    port map (
            O => \N__34740\,
            I => \N__34736\
        );

    \I__6174\ : InMux
    port map (
            O => \N__34739\,
            I => \N__34733\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__34736\,
            I => \N__34730\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__34733\,
            I => \N__34727\
        );

    \I__6171\ : Span4Mux_h
    port map (
            O => \N__34730\,
            I => \N__34724\
        );

    \I__6170\ : Span12Mux_s4_h
    port map (
            O => \N__34727\,
            I => \N__34721\
        );

    \I__6169\ : Odrv4
    port map (
            O => \N__34724\,
            I => n15418
        );

    \I__6168\ : Odrv12
    port map (
            O => \N__34721\,
            I => n15418
        );

    \I__6167\ : CascadeMux
    port map (
            O => \N__34716\,
            I => \N__34711\
        );

    \I__6166\ : InMux
    port map (
            O => \N__34715\,
            I => \N__34705\
        );

    \I__6165\ : CascadeMux
    port map (
            O => \N__34714\,
            I => \N__34700\
        );

    \I__6164\ : InMux
    port map (
            O => \N__34711\,
            I => \N__34690\
        );

    \I__6163\ : InMux
    port map (
            O => \N__34710\,
            I => \N__34690\
        );

    \I__6162\ : CascadeMux
    port map (
            O => \N__34709\,
            I => \N__34687\
        );

    \I__6161\ : CascadeMux
    port map (
            O => \N__34708\,
            I => \N__34683\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__34705\,
            I => \N__34678\
        );

    \I__6159\ : InMux
    port map (
            O => \N__34704\,
            I => \N__34673\
        );

    \I__6158\ : InMux
    port map (
            O => \N__34703\,
            I => \N__34673\
        );

    \I__6157\ : InMux
    port map (
            O => \N__34700\,
            I => \N__34666\
        );

    \I__6156\ : InMux
    port map (
            O => \N__34699\,
            I => \N__34666\
        );

    \I__6155\ : InMux
    port map (
            O => \N__34698\,
            I => \N__34666\
        );

    \I__6154\ : CascadeMux
    port map (
            O => \N__34697\,
            I => \N__34661\
        );

    \I__6153\ : CascadeMux
    port map (
            O => \N__34696\,
            I => \N__34654\
        );

    \I__6152\ : CascadeMux
    port map (
            O => \N__34695\,
            I => \N__34650\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__34690\,
            I => \N__34646\
        );

    \I__6150\ : InMux
    port map (
            O => \N__34687\,
            I => \N__34635\
        );

    \I__6149\ : InMux
    port map (
            O => \N__34686\,
            I => \N__34635\
        );

    \I__6148\ : InMux
    port map (
            O => \N__34683\,
            I => \N__34635\
        );

    \I__6147\ : InMux
    port map (
            O => \N__34682\,
            I => \N__34635\
        );

    \I__6146\ : InMux
    port map (
            O => \N__34681\,
            I => \N__34635\
        );

    \I__6145\ : Span4Mux_v
    port map (
            O => \N__34678\,
            I => \N__34632\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__34673\,
            I => \N__34627\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__34666\,
            I => \N__34627\
        );

    \I__6142\ : InMux
    port map (
            O => \N__34665\,
            I => \N__34620\
        );

    \I__6141\ : InMux
    port map (
            O => \N__34664\,
            I => \N__34620\
        );

    \I__6140\ : InMux
    port map (
            O => \N__34661\,
            I => \N__34620\
        );

    \I__6139\ : InMux
    port map (
            O => \N__34660\,
            I => \N__34617\
        );

    \I__6138\ : InMux
    port map (
            O => \N__34659\,
            I => \N__34614\
        );

    \I__6137\ : CascadeMux
    port map (
            O => \N__34658\,
            I => \N__34608\
        );

    \I__6136\ : CascadeMux
    port map (
            O => \N__34657\,
            I => \N__34605\
        );

    \I__6135\ : InMux
    port map (
            O => \N__34654\,
            I => \N__34594\
        );

    \I__6134\ : InMux
    port map (
            O => \N__34653\,
            I => \N__34594\
        );

    \I__6133\ : InMux
    port map (
            O => \N__34650\,
            I => \N__34594\
        );

    \I__6132\ : InMux
    port map (
            O => \N__34649\,
            I => \N__34594\
        );

    \I__6131\ : Span4Mux_s1_h
    port map (
            O => \N__34646\,
            I => \N__34589\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__34635\,
            I => \N__34589\
        );

    \I__6129\ : Span4Mux_h
    port map (
            O => \N__34632\,
            I => \N__34582\
        );

    \I__6128\ : Span4Mux_s1_v
    port map (
            O => \N__34627\,
            I => \N__34582\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__34620\,
            I => \N__34582\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__34617\,
            I => \N__34579\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__34614\,
            I => \N__34576\
        );

    \I__6124\ : InMux
    port map (
            O => \N__34613\,
            I => \N__34563\
        );

    \I__6123\ : InMux
    port map (
            O => \N__34612\,
            I => \N__34563\
        );

    \I__6122\ : InMux
    port map (
            O => \N__34611\,
            I => \N__34563\
        );

    \I__6121\ : InMux
    port map (
            O => \N__34608\,
            I => \N__34563\
        );

    \I__6120\ : InMux
    port map (
            O => \N__34605\,
            I => \N__34563\
        );

    \I__6119\ : InMux
    port map (
            O => \N__34604\,
            I => \N__34563\
        );

    \I__6118\ : InMux
    port map (
            O => \N__34603\,
            I => \N__34560\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__34594\,
            I => \N__34555\
        );

    \I__6116\ : Span4Mux_v
    port map (
            O => \N__34589\,
            I => \N__34555\
        );

    \I__6115\ : Odrv4
    port map (
            O => \N__34582\,
            I => n3039
        );

    \I__6114\ : Odrv4
    port map (
            O => \N__34579\,
            I => n3039
        );

    \I__6113\ : Odrv4
    port map (
            O => \N__34576\,
            I => n3039
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__34563\,
            I => n3039
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__34560\,
            I => n3039
        );

    \I__6110\ : Odrv4
    port map (
            O => \N__34555\,
            I => n3039
        );

    \I__6109\ : InMux
    port map (
            O => \N__34542\,
            I => n12954
        );

    \I__6108\ : InMux
    port map (
            O => \N__34539\,
            I => \N__34536\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__34536\,
            I => \N__34533\
        );

    \I__6106\ : Span4Mux_h
    port map (
            O => \N__34533\,
            I => \N__34529\
        );

    \I__6105\ : CascadeMux
    port map (
            O => \N__34532\,
            I => \N__34526\
        );

    \I__6104\ : Span4Mux_h
    port map (
            O => \N__34529\,
            I => \N__34523\
        );

    \I__6103\ : InMux
    port map (
            O => \N__34526\,
            I => \N__34520\
        );

    \I__6102\ : Odrv4
    port map (
            O => \N__34523\,
            I => n15384
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__34520\,
            I => n15384
        );

    \I__6100\ : InMux
    port map (
            O => \N__34515\,
            I => \N__34506\
        );

    \I__6099\ : InMux
    port map (
            O => \N__34514\,
            I => \N__34499\
        );

    \I__6098\ : InMux
    port map (
            O => \N__34513\,
            I => \N__34494\
        );

    \I__6097\ : InMux
    port map (
            O => \N__34512\,
            I => \N__34494\
        );

    \I__6096\ : CascadeMux
    port map (
            O => \N__34511\,
            I => \N__34490\
        );

    \I__6095\ : CascadeMux
    port map (
            O => \N__34510\,
            I => \N__34487\
        );

    \I__6094\ : CascadeMux
    port map (
            O => \N__34509\,
            I => \N__34484\
        );

    \I__6093\ : LocalMux
    port map (
            O => \N__34506\,
            I => \N__34480\
        );

    \I__6092\ : InMux
    port map (
            O => \N__34505\,
            I => \N__34476\
        );

    \I__6091\ : CascadeMux
    port map (
            O => \N__34504\,
            I => \N__34469\
        );

    \I__6090\ : CascadeMux
    port map (
            O => \N__34503\,
            I => \N__34463\
        );

    \I__6089\ : CascadeMux
    port map (
            O => \N__34502\,
            I => \N__34455\
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__34499\,
            I => \N__34450\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__34494\,
            I => \N__34447\
        );

    \I__6086\ : InMux
    port map (
            O => \N__34493\,
            I => \N__34436\
        );

    \I__6085\ : InMux
    port map (
            O => \N__34490\,
            I => \N__34436\
        );

    \I__6084\ : InMux
    port map (
            O => \N__34487\,
            I => \N__34436\
        );

    \I__6083\ : InMux
    port map (
            O => \N__34484\,
            I => \N__34436\
        );

    \I__6082\ : InMux
    port map (
            O => \N__34483\,
            I => \N__34436\
        );

    \I__6081\ : Span4Mux_h
    port map (
            O => \N__34480\,
            I => \N__34433\
        );

    \I__6080\ : InMux
    port map (
            O => \N__34479\,
            I => \N__34430\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__34476\,
            I => \N__34427\
        );

    \I__6078\ : InMux
    port map (
            O => \N__34475\,
            I => \N__34420\
        );

    \I__6077\ : InMux
    port map (
            O => \N__34474\,
            I => \N__34420\
        );

    \I__6076\ : InMux
    port map (
            O => \N__34473\,
            I => \N__34420\
        );

    \I__6075\ : InMux
    port map (
            O => \N__34472\,
            I => \N__34413\
        );

    \I__6074\ : InMux
    port map (
            O => \N__34469\,
            I => \N__34413\
        );

    \I__6073\ : InMux
    port map (
            O => \N__34468\,
            I => \N__34413\
        );

    \I__6072\ : InMux
    port map (
            O => \N__34467\,
            I => \N__34406\
        );

    \I__6071\ : InMux
    port map (
            O => \N__34466\,
            I => \N__34406\
        );

    \I__6070\ : InMux
    port map (
            O => \N__34463\,
            I => \N__34406\
        );

    \I__6069\ : InMux
    port map (
            O => \N__34462\,
            I => \N__34403\
        );

    \I__6068\ : InMux
    port map (
            O => \N__34461\,
            I => \N__34398\
        );

    \I__6067\ : InMux
    port map (
            O => \N__34460\,
            I => \N__34398\
        );

    \I__6066\ : InMux
    port map (
            O => \N__34459\,
            I => \N__34387\
        );

    \I__6065\ : InMux
    port map (
            O => \N__34458\,
            I => \N__34387\
        );

    \I__6064\ : InMux
    port map (
            O => \N__34455\,
            I => \N__34387\
        );

    \I__6063\ : InMux
    port map (
            O => \N__34454\,
            I => \N__34387\
        );

    \I__6062\ : InMux
    port map (
            O => \N__34453\,
            I => \N__34387\
        );

    \I__6061\ : Span4Mux_v
    port map (
            O => \N__34450\,
            I => \N__34380\
        );

    \I__6060\ : Span4Mux_v
    port map (
            O => \N__34447\,
            I => \N__34380\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__34436\,
            I => \N__34380\
        );

    \I__6058\ : Odrv4
    port map (
            O => \N__34433\,
            I => n2940
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__34430\,
            I => n2940
        );

    \I__6056\ : Odrv4
    port map (
            O => \N__34427\,
            I => n2940
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__34420\,
            I => n2940
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__34413\,
            I => n2940
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__34406\,
            I => n2940
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__34403\,
            I => n2940
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__34398\,
            I => n2940
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__34387\,
            I => n2940
        );

    \I__6049\ : Odrv4
    port map (
            O => \N__34380\,
            I => n2940
        );

    \I__6048\ : InMux
    port map (
            O => \N__34359\,
            I => n12955
        );

    \I__6047\ : InMux
    port map (
            O => \N__34356\,
            I => \N__34353\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__34353\,
            I => \N__34349\
        );

    \I__6045\ : InMux
    port map (
            O => \N__34352\,
            I => \N__34346\
        );

    \I__6044\ : Span4Mux_h
    port map (
            O => \N__34349\,
            I => \N__34341\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__34346\,
            I => \N__34341\
        );

    \I__6042\ : Span4Mux_s3_h
    port map (
            O => \N__34341\,
            I => \N__34338\
        );

    \I__6041\ : Odrv4
    port map (
            O => \N__34338\,
            I => n15352
        );

    \I__6040\ : CascadeMux
    port map (
            O => \N__34335\,
            I => \N__34329\
        );

    \I__6039\ : InMux
    port map (
            O => \N__34334\,
            I => \N__34325\
        );

    \I__6038\ : CascadeMux
    port map (
            O => \N__34333\,
            I => \N__34317\
        );

    \I__6037\ : InMux
    port map (
            O => \N__34332\,
            I => \N__34311\
        );

    \I__6036\ : InMux
    port map (
            O => \N__34329\,
            I => \N__34306\
        );

    \I__6035\ : InMux
    port map (
            O => \N__34328\,
            I => \N__34306\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__34325\,
            I => \N__34303\
        );

    \I__6033\ : CascadeMux
    port map (
            O => \N__34324\,
            I => \N__34298\
        );

    \I__6032\ : CascadeMux
    port map (
            O => \N__34323\,
            I => \N__34294\
        );

    \I__6031\ : InMux
    port map (
            O => \N__34322\,
            I => \N__34286\
        );

    \I__6030\ : CascadeMux
    port map (
            O => \N__34321\,
            I => \N__34283\
        );

    \I__6029\ : CascadeMux
    port map (
            O => \N__34320\,
            I => \N__34279\
        );

    \I__6028\ : InMux
    port map (
            O => \N__34317\,
            I => \N__34272\
        );

    \I__6027\ : InMux
    port map (
            O => \N__34316\,
            I => \N__34272\
        );

    \I__6026\ : CascadeMux
    port map (
            O => \N__34315\,
            I => \N__34268\
        );

    \I__6025\ : CascadeMux
    port map (
            O => \N__34314\,
            I => \N__34264\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__34311\,
            I => \N__34260\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__34306\,
            I => \N__34257\
        );

    \I__6022\ : Span4Mux_h
    port map (
            O => \N__34303\,
            I => \N__34254\
        );

    \I__6021\ : InMux
    port map (
            O => \N__34302\,
            I => \N__34249\
        );

    \I__6020\ : InMux
    port map (
            O => \N__34301\,
            I => \N__34249\
        );

    \I__6019\ : InMux
    port map (
            O => \N__34298\,
            I => \N__34244\
        );

    \I__6018\ : InMux
    port map (
            O => \N__34297\,
            I => \N__34244\
        );

    \I__6017\ : InMux
    port map (
            O => \N__34294\,
            I => \N__34239\
        );

    \I__6016\ : InMux
    port map (
            O => \N__34293\,
            I => \N__34239\
        );

    \I__6015\ : InMux
    port map (
            O => \N__34292\,
            I => \N__34230\
        );

    \I__6014\ : InMux
    port map (
            O => \N__34291\,
            I => \N__34230\
        );

    \I__6013\ : InMux
    port map (
            O => \N__34290\,
            I => \N__34230\
        );

    \I__6012\ : InMux
    port map (
            O => \N__34289\,
            I => \N__34230\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__34286\,
            I => \N__34227\
        );

    \I__6010\ : InMux
    port map (
            O => \N__34283\,
            I => \N__34222\
        );

    \I__6009\ : InMux
    port map (
            O => \N__34282\,
            I => \N__34222\
        );

    \I__6008\ : InMux
    port map (
            O => \N__34279\,
            I => \N__34215\
        );

    \I__6007\ : InMux
    port map (
            O => \N__34278\,
            I => \N__34215\
        );

    \I__6006\ : InMux
    port map (
            O => \N__34277\,
            I => \N__34215\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__34272\,
            I => \N__34212\
        );

    \I__6004\ : InMux
    port map (
            O => \N__34271\,
            I => \N__34201\
        );

    \I__6003\ : InMux
    port map (
            O => \N__34268\,
            I => \N__34201\
        );

    \I__6002\ : InMux
    port map (
            O => \N__34267\,
            I => \N__34201\
        );

    \I__6001\ : InMux
    port map (
            O => \N__34264\,
            I => \N__34201\
        );

    \I__6000\ : InMux
    port map (
            O => \N__34263\,
            I => \N__34201\
        );

    \I__5999\ : Span4Mux_v
    port map (
            O => \N__34260\,
            I => \N__34196\
        );

    \I__5998\ : Span4Mux_s3_h
    port map (
            O => \N__34257\,
            I => \N__34196\
        );

    \I__5997\ : Odrv4
    port map (
            O => \N__34254\,
            I => n2841
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__34249\,
            I => n2841
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__34244\,
            I => n2841
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__34239\,
            I => n2841
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__34230\,
            I => n2841
        );

    \I__5992\ : Odrv4
    port map (
            O => \N__34227\,
            I => n2841
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__34222\,
            I => n2841
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__34215\,
            I => n2841
        );

    \I__5989\ : Odrv4
    port map (
            O => \N__34212\,
            I => n2841
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__34201\,
            I => n2841
        );

    \I__5987\ : Odrv4
    port map (
            O => \N__34196\,
            I => n2841
        );

    \I__5986\ : InMux
    port map (
            O => \N__34173\,
            I => n12956
        );

    \I__5985\ : InMux
    port map (
            O => \N__34170\,
            I => \N__34167\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__34167\,
            I => \N__34162\
        );

    \I__5983\ : InMux
    port map (
            O => \N__34166\,
            I => \N__34159\
        );

    \I__5982\ : InMux
    port map (
            O => \N__34165\,
            I => \N__34156\
        );

    \I__5981\ : Span4Mux_s3_h
    port map (
            O => \N__34162\,
            I => \N__34151\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__34159\,
            I => \N__34151\
        );

    \I__5979\ : LocalMux
    port map (
            O => \N__34156\,
            I => \N__34148\
        );

    \I__5978\ : Span4Mux_h
    port map (
            O => \N__34151\,
            I => \N__34145\
        );

    \I__5977\ : Sp12to4
    port map (
            O => \N__34148\,
            I => \N__34142\
        );

    \I__5976\ : Span4Mux_v
    port map (
            O => \N__34145\,
            I => \N__34139\
        );

    \I__5975\ : Odrv12
    port map (
            O => \N__34142\,
            I => n317
        );

    \I__5974\ : Odrv4
    port map (
            O => \N__34139\,
            I => n317
        );

    \I__5973\ : InMux
    port map (
            O => \N__34134\,
            I => \N__34131\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__34131\,
            I => \N__34128\
        );

    \I__5971\ : Odrv4
    port map (
            O => \N__34128\,
            I => n14184
        );

    \I__5970\ : InMux
    port map (
            O => \N__34125\,
            I => \N__34122\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__34122\,
            I => n2490
        );

    \I__5968\ : CascadeMux
    port map (
            O => \N__34119\,
            I => \N__34115\
        );

    \I__5967\ : InMux
    port map (
            O => \N__34118\,
            I => \N__34112\
        );

    \I__5966\ : InMux
    port map (
            O => \N__34115\,
            I => \N__34109\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__34112\,
            I => \N__34106\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__34109\,
            I => \N__34103\
        );

    \I__5963\ : Span4Mux_v
    port map (
            O => \N__34106\,
            I => \N__34099\
        );

    \I__5962\ : Span4Mux_h
    port map (
            O => \N__34103\,
            I => \N__34096\
        );

    \I__5961\ : InMux
    port map (
            O => \N__34102\,
            I => \N__34093\
        );

    \I__5960\ : Odrv4
    port map (
            O => \N__34099\,
            I => n2423
        );

    \I__5959\ : Odrv4
    port map (
            O => \N__34096\,
            I => n2423
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__34093\,
            I => n2423
        );

    \I__5957\ : InMux
    port map (
            O => \N__34086\,
            I => \N__34083\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__34083\,
            I => \N__34079\
        );

    \I__5955\ : CascadeMux
    port map (
            O => \N__34082\,
            I => \N__34076\
        );

    \I__5954\ : Span4Mux_v
    port map (
            O => \N__34079\,
            I => \N__34072\
        );

    \I__5953\ : InMux
    port map (
            O => \N__34076\,
            I => \N__34069\
        );

    \I__5952\ : CascadeMux
    port map (
            O => \N__34075\,
            I => \N__34066\
        );

    \I__5951\ : Span4Mux_h
    port map (
            O => \N__34072\,
            I => \N__34061\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__34069\,
            I => \N__34061\
        );

    \I__5949\ : InMux
    port map (
            O => \N__34066\,
            I => \N__34058\
        );

    \I__5948\ : Odrv4
    port map (
            O => \N__34061\,
            I => n2522
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__34058\,
            I => n2522
        );

    \I__5946\ : InMux
    port map (
            O => \N__34053\,
            I => \N__34050\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__34050\,
            I => n2489
        );

    \I__5944\ : CascadeMux
    port map (
            O => \N__34047\,
            I => \N__34044\
        );

    \I__5943\ : InMux
    port map (
            O => \N__34044\,
            I => \N__34040\
        );

    \I__5942\ : CascadeMux
    port map (
            O => \N__34043\,
            I => \N__34037\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__34040\,
            I => \N__34034\
        );

    \I__5940\ : InMux
    port map (
            O => \N__34037\,
            I => \N__34031\
        );

    \I__5939\ : Span4Mux_v
    port map (
            O => \N__34034\,
            I => \N__34027\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__34031\,
            I => \N__34024\
        );

    \I__5937\ : InMux
    port map (
            O => \N__34030\,
            I => \N__34021\
        );

    \I__5936\ : Odrv4
    port map (
            O => \N__34027\,
            I => n2422
        );

    \I__5935\ : Odrv4
    port map (
            O => \N__34024\,
            I => n2422
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__34021\,
            I => n2422
        );

    \I__5933\ : CascadeMux
    port map (
            O => \N__34014\,
            I => \N__34011\
        );

    \I__5932\ : InMux
    port map (
            O => \N__34011\,
            I => \N__34007\
        );

    \I__5931\ : CascadeMux
    port map (
            O => \N__34010\,
            I => \N__34004\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__34007\,
            I => \N__34001\
        );

    \I__5929\ : InMux
    port map (
            O => \N__34004\,
            I => \N__33998\
        );

    \I__5928\ : Span4Mux_h
    port map (
            O => \N__34001\,
            I => \N__33992\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__33998\,
            I => \N__33992\
        );

    \I__5926\ : InMux
    port map (
            O => \N__33997\,
            I => \N__33989\
        );

    \I__5925\ : Odrv4
    port map (
            O => \N__33992\,
            I => n2521
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__33989\,
            I => n2521
        );

    \I__5923\ : CascadeMux
    port map (
            O => \N__33984\,
            I => \N__33980\
        );

    \I__5922\ : InMux
    port map (
            O => \N__33983\,
            I => \N__33977\
        );

    \I__5921\ : InMux
    port map (
            O => \N__33980\,
            I => \N__33974\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__33977\,
            I => \N__33969\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__33974\,
            I => \N__33969\
        );

    \I__5918\ : Span4Mux_v
    port map (
            O => \N__33969\,
            I => \N__33965\
        );

    \I__5917\ : InMux
    port map (
            O => \N__33968\,
            I => \N__33962\
        );

    \I__5916\ : Odrv4
    port map (
            O => \N__33965\,
            I => n2426
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__33962\,
            I => n2426
        );

    \I__5914\ : InMux
    port map (
            O => \N__33957\,
            I => \N__33954\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__33954\,
            I => n2493
        );

    \I__5912\ : CascadeMux
    port map (
            O => \N__33951\,
            I => \N__33948\
        );

    \I__5911\ : InMux
    port map (
            O => \N__33948\,
            I => \N__33945\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__33945\,
            I => \N__33941\
        );

    \I__5909\ : InMux
    port map (
            O => \N__33944\,
            I => \N__33938\
        );

    \I__5908\ : Odrv4
    port map (
            O => \N__33941\,
            I => n2525
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__33938\,
            I => n2525
        );

    \I__5906\ : InMux
    port map (
            O => \N__33933\,
            I => \N__33930\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__33930\,
            I => \N__33927\
        );

    \I__5904\ : Odrv4
    port map (
            O => \N__33927\,
            I => n2592
        );

    \I__5903\ : CascadeMux
    port map (
            O => \N__33924\,
            I => \n2525_cascade_\
        );

    \I__5902\ : CascadeMux
    port map (
            O => \N__33921\,
            I => \N__33918\
        );

    \I__5901\ : InMux
    port map (
            O => \N__33918\,
            I => \N__33914\
        );

    \I__5900\ : InMux
    port map (
            O => \N__33917\,
            I => \N__33911\
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__33914\,
            I => \N__33908\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__33911\,
            I => \N__33904\
        );

    \I__5897\ : Span4Mux_v
    port map (
            O => \N__33908\,
            I => \N__33901\
        );

    \I__5896\ : InMux
    port map (
            O => \N__33907\,
            I => \N__33898\
        );

    \I__5895\ : Span4Mux_v
    port map (
            O => \N__33904\,
            I => \N__33891\
        );

    \I__5894\ : Span4Mux_v
    port map (
            O => \N__33901\,
            I => \N__33891\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__33898\,
            I => \N__33891\
        );

    \I__5892\ : Span4Mux_h
    port map (
            O => \N__33891\,
            I => \N__33888\
        );

    \I__5891\ : Odrv4
    port map (
            O => \N__33888\,
            I => n2624
        );

    \I__5890\ : InMux
    port map (
            O => \N__33885\,
            I => \N__33882\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__33882\,
            I => n2486
        );

    \I__5888\ : CascadeMux
    port map (
            O => \N__33879\,
            I => \N__33875\
        );

    \I__5887\ : CascadeMux
    port map (
            O => \N__33878\,
            I => \N__33872\
        );

    \I__5886\ : InMux
    port map (
            O => \N__33875\,
            I => \N__33868\
        );

    \I__5885\ : InMux
    port map (
            O => \N__33872\,
            I => \N__33865\
        );

    \I__5884\ : CascadeMux
    port map (
            O => \N__33871\,
            I => \N__33862\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__33868\,
            I => \N__33859\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__33865\,
            I => \N__33856\
        );

    \I__5881\ : InMux
    port map (
            O => \N__33862\,
            I => \N__33853\
        );

    \I__5880\ : Span4Mux_v
    port map (
            O => \N__33859\,
            I => \N__33850\
        );

    \I__5879\ : Span4Mux_h
    port map (
            O => \N__33856\,
            I => \N__33845\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__33853\,
            I => \N__33845\
        );

    \I__5877\ : Odrv4
    port map (
            O => \N__33850\,
            I => n2419
        );

    \I__5876\ : Odrv4
    port map (
            O => \N__33845\,
            I => n2419
        );

    \I__5875\ : InMux
    port map (
            O => \N__33840\,
            I => \N__33836\
        );

    \I__5874\ : InMux
    port map (
            O => \N__33839\,
            I => \N__33833\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__33836\,
            I => \N__33829\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__33833\,
            I => \N__33826\
        );

    \I__5871\ : InMux
    port map (
            O => \N__33832\,
            I => \N__33823\
        );

    \I__5870\ : Odrv4
    port map (
            O => \N__33829\,
            I => n2518
        );

    \I__5869\ : Odrv4
    port map (
            O => \N__33826\,
            I => n2518
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__33823\,
            I => n2518
        );

    \I__5867\ : InMux
    port map (
            O => \N__33816\,
            I => \N__33813\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__33813\,
            I => n11981
        );

    \I__5865\ : InMux
    port map (
            O => \N__33810\,
            I => \N__33807\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__33807\,
            I => \N__33802\
        );

    \I__5863\ : CascadeMux
    port map (
            O => \N__33806\,
            I => \N__33799\
        );

    \I__5862\ : InMux
    port map (
            O => \N__33805\,
            I => \N__33796\
        );

    \I__5861\ : Span4Mux_h
    port map (
            O => \N__33802\,
            I => \N__33793\
        );

    \I__5860\ : InMux
    port map (
            O => \N__33799\,
            I => \N__33790\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__33796\,
            I => \N__33787\
        );

    \I__5858\ : Odrv4
    port map (
            O => \N__33793\,
            I => n2029
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__33790\,
            I => n2029
        );

    \I__5856\ : Odrv4
    port map (
            O => \N__33787\,
            I => n2029
        );

    \I__5855\ : CascadeMux
    port map (
            O => \N__33780\,
            I => \n14550_cascade_\
        );

    \I__5854\ : InMux
    port map (
            O => \N__33777\,
            I => \N__33772\
        );

    \I__5853\ : CascadeMux
    port map (
            O => \N__33776\,
            I => \N__33769\
        );

    \I__5852\ : InMux
    port map (
            O => \N__33775\,
            I => \N__33766\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__33772\,
            I => \N__33763\
        );

    \I__5850\ : InMux
    port map (
            O => \N__33769\,
            I => \N__33760\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__33766\,
            I => \N__33757\
        );

    \I__5848\ : Odrv4
    port map (
            O => \N__33763\,
            I => n2030
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__33760\,
            I => n2030
        );

    \I__5846\ : Odrv12
    port map (
            O => \N__33757\,
            I => n2030
        );

    \I__5845\ : InMux
    port map (
            O => \N__33750\,
            I => \N__33747\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__33747\,
            I => n14552
        );

    \I__5843\ : InMux
    port map (
            O => \N__33744\,
            I => \N__33741\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__33741\,
            I => \N__33738\
        );

    \I__5841\ : Span4Mux_v
    port map (
            O => \N__33738\,
            I => \N__33735\
        );

    \I__5840\ : Odrv4
    port map (
            O => \N__33735\,
            I => n2100
        );

    \I__5839\ : CascadeMux
    port map (
            O => \N__33732\,
            I => \N__33728\
        );

    \I__5838\ : CascadeMux
    port map (
            O => \N__33731\,
            I => \N__33725\
        );

    \I__5837\ : InMux
    port map (
            O => \N__33728\,
            I => \N__33722\
        );

    \I__5836\ : InMux
    port map (
            O => \N__33725\,
            I => \N__33718\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__33722\,
            I => \N__33715\
        );

    \I__5834\ : InMux
    port map (
            O => \N__33721\,
            I => \N__33712\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__33718\,
            I => n2033
        );

    \I__5832\ : Odrv4
    port map (
            O => \N__33715\,
            I => n2033
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__33712\,
            I => n2033
        );

    \I__5830\ : InMux
    port map (
            O => \N__33705\,
            I => \N__33701\
        );

    \I__5829\ : CascadeMux
    port map (
            O => \N__33704\,
            I => \N__33698\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__33701\,
            I => \N__33695\
        );

    \I__5827\ : InMux
    port map (
            O => \N__33698\,
            I => \N__33692\
        );

    \I__5826\ : Span4Mux_v
    port map (
            O => \N__33695\,
            I => \N__33687\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__33692\,
            I => \N__33687\
        );

    \I__5824\ : Span4Mux_v
    port map (
            O => \N__33687\,
            I => \N__33684\
        );

    \I__5823\ : Odrv4
    port map (
            O => \N__33684\,
            I => n2132
        );

    \I__5822\ : CascadeMux
    port map (
            O => \N__33681\,
            I => \n2132_cascade_\
        );

    \I__5821\ : CascadeMux
    port map (
            O => \N__33678\,
            I => \N__33674\
        );

    \I__5820\ : InMux
    port map (
            O => \N__33677\,
            I => \N__33671\
        );

    \I__5819\ : InMux
    port map (
            O => \N__33674\,
            I => \N__33668\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__33671\,
            I => \N__33665\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__33668\,
            I => \N__33662\
        );

    \I__5816\ : Span12Mux_v
    port map (
            O => \N__33665\,
            I => \N__33658\
        );

    \I__5815\ : Span4Mux_h
    port map (
            O => \N__33662\,
            I => \N__33655\
        );

    \I__5814\ : InMux
    port map (
            O => \N__33661\,
            I => \N__33652\
        );

    \I__5813\ : Odrv12
    port map (
            O => \N__33658\,
            I => n2133
        );

    \I__5812\ : Odrv4
    port map (
            O => \N__33655\,
            I => n2133
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__33652\,
            I => n2133
        );

    \I__5810\ : InMux
    port map (
            O => \N__33645\,
            I => \N__33642\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__33642\,
            I => \N__33639\
        );

    \I__5808\ : Span4Mux_h
    port map (
            O => \N__33639\,
            I => \N__33636\
        );

    \I__5807\ : Odrv4
    port map (
            O => \N__33636\,
            I => n11909
        );

    \I__5806\ : InMux
    port map (
            O => \N__33633\,
            I => \N__33629\
        );

    \I__5805\ : InMux
    port map (
            O => \N__33632\,
            I => \N__33626\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__33629\,
            I => \N__33621\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__33626\,
            I => \N__33621\
        );

    \I__5802\ : Span4Mux_h
    port map (
            O => \N__33621\,
            I => \N__33617\
        );

    \I__5801\ : InMux
    port map (
            O => \N__33620\,
            I => \N__33614\
        );

    \I__5800\ : Odrv4
    port map (
            O => \N__33617\,
            I => n307
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__33614\,
            I => n307
        );

    \I__5798\ : InMux
    port map (
            O => \N__33609\,
            I => \N__33606\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__33606\,
            I => \N__33602\
        );

    \I__5796\ : InMux
    port map (
            O => \N__33605\,
            I => \N__33598\
        );

    \I__5795\ : Span4Mux_h
    port map (
            O => \N__33602\,
            I => \N__33595\
        );

    \I__5794\ : InMux
    port map (
            O => \N__33601\,
            I => \N__33592\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__33598\,
            I => \N__33589\
        );

    \I__5792\ : Odrv4
    port map (
            O => \N__33595\,
            I => n310
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__33592\,
            I => n310
        );

    \I__5790\ : Odrv12
    port map (
            O => \N__33589\,
            I => n310
        );

    \I__5789\ : InMux
    port map (
            O => \N__33582\,
            I => \N__33578\
        );

    \I__5788\ : InMux
    port map (
            O => \N__33581\,
            I => \N__33574\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__33578\,
            I => \N__33571\
        );

    \I__5786\ : InMux
    port map (
            O => \N__33577\,
            I => \N__33568\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__33574\,
            I => \N__33565\
        );

    \I__5784\ : Span4Mux_s2_h
    port map (
            O => \N__33571\,
            I => \N__33562\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__33568\,
            I => \N__33559\
        );

    \I__5782\ : Span4Mux_v
    port map (
            O => \N__33565\,
            I => \N__33556\
        );

    \I__5781\ : Span4Mux_v
    port map (
            O => \N__33562\,
            I => \N__33553\
        );

    \I__5780\ : Span4Mux_v
    port map (
            O => \N__33559\,
            I => \N__33548\
        );

    \I__5779\ : Span4Mux_s3_h
    port map (
            O => \N__33556\,
            I => \N__33548\
        );

    \I__5778\ : Span4Mux_h
    port map (
            O => \N__33553\,
            I => \N__33545\
        );

    \I__5777\ : Odrv4
    port map (
            O => \N__33548\,
            I => n312
        );

    \I__5776\ : Odrv4
    port map (
            O => \N__33545\,
            I => n312
        );

    \I__5775\ : InMux
    port map (
            O => \N__33540\,
            I => \N__33536\
        );

    \I__5774\ : InMux
    port map (
            O => \N__33539\,
            I => \N__33533\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__33536\,
            I => \N__33530\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__33533\,
            I => \N__33527\
        );

    \I__5771\ : Span4Mux_v
    port map (
            O => \N__33530\,
            I => \N__33524\
        );

    \I__5770\ : Span4Mux_v
    port map (
            O => \N__33527\,
            I => \N__33520\
        );

    \I__5769\ : Span4Mux_h
    port map (
            O => \N__33524\,
            I => \N__33517\
        );

    \I__5768\ : InMux
    port map (
            O => \N__33523\,
            I => \N__33514\
        );

    \I__5767\ : Span4Mux_h
    port map (
            O => \N__33520\,
            I => \N__33509\
        );

    \I__5766\ : Span4Mux_v
    port map (
            O => \N__33517\,
            I => \N__33509\
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__33514\,
            I => \N__33506\
        );

    \I__5764\ : Odrv4
    port map (
            O => \N__33509\,
            I => n313
        );

    \I__5763\ : Odrv12
    port map (
            O => \N__33506\,
            I => n313
        );

    \I__5762\ : InMux
    port map (
            O => \N__33501\,
            I => \N__33497\
        );

    \I__5761\ : InMux
    port map (
            O => \N__33500\,
            I => \N__33493\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__33497\,
            I => \N__33490\
        );

    \I__5759\ : InMux
    port map (
            O => \N__33496\,
            I => \N__33487\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__33493\,
            I => \N__33484\
        );

    \I__5757\ : Span4Mux_s1_h
    port map (
            O => \N__33490\,
            I => \N__33481\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__33487\,
            I => \N__33478\
        );

    \I__5755\ : Span4Mux_v
    port map (
            O => \N__33484\,
            I => \N__33473\
        );

    \I__5754\ : Span4Mux_h
    port map (
            O => \N__33481\,
            I => \N__33473\
        );

    \I__5753\ : Span4Mux_h
    port map (
            O => \N__33478\,
            I => \N__33470\
        );

    \I__5752\ : Odrv4
    port map (
            O => \N__33473\,
            I => n314
        );

    \I__5751\ : Odrv4
    port map (
            O => \N__33470\,
            I => n314
        );

    \I__5750\ : InMux
    port map (
            O => \N__33465\,
            I => \N__33461\
        );

    \I__5749\ : CascadeMux
    port map (
            O => \N__33464\,
            I => \N__33458\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__33461\,
            I => \N__33455\
        );

    \I__5747\ : InMux
    port map (
            O => \N__33458\,
            I => \N__33452\
        );

    \I__5746\ : Odrv4
    port map (
            O => \N__33455\,
            I => n2025
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__33452\,
            I => n2025
        );

    \I__5744\ : InMux
    port map (
            O => \N__33447\,
            I => \N__33444\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__33444\,
            I => \N__33440\
        );

    \I__5742\ : CascadeMux
    port map (
            O => \N__33443\,
            I => \N__33437\
        );

    \I__5741\ : Span4Mux_v
    port map (
            O => \N__33440\,
            I => \N__33433\
        );

    \I__5740\ : InMux
    port map (
            O => \N__33437\,
            I => \N__33430\
        );

    \I__5739\ : InMux
    port map (
            O => \N__33436\,
            I => \N__33427\
        );

    \I__5738\ : Odrv4
    port map (
            O => \N__33433\,
            I => n2028
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__33430\,
            I => n2028
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__33427\,
            I => n2028
        );

    \I__5735\ : InMux
    port map (
            O => \N__33420\,
            I => \N__33416\
        );

    \I__5734\ : CascadeMux
    port map (
            O => \N__33419\,
            I => \N__33413\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__33416\,
            I => \N__33409\
        );

    \I__5732\ : InMux
    port map (
            O => \N__33413\,
            I => \N__33406\
        );

    \I__5731\ : InMux
    port map (
            O => \N__33412\,
            I => \N__33403\
        );

    \I__5730\ : Odrv4
    port map (
            O => \N__33409\,
            I => n2026
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__33406\,
            I => n2026
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__33403\,
            I => n2026
        );

    \I__5727\ : CascadeMux
    port map (
            O => \N__33396\,
            I => \n2025_cascade_\
        );

    \I__5726\ : InMux
    port map (
            O => \N__33393\,
            I => \N__33389\
        );

    \I__5725\ : CascadeMux
    port map (
            O => \N__33392\,
            I => \N__33386\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__33389\,
            I => \N__33382\
        );

    \I__5723\ : InMux
    port map (
            O => \N__33386\,
            I => \N__33379\
        );

    \I__5722\ : InMux
    port map (
            O => \N__33385\,
            I => \N__33376\
        );

    \I__5721\ : Odrv4
    port map (
            O => \N__33382\,
            I => n2027
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__33379\,
            I => n2027
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__33376\,
            I => n2027
        );

    \I__5718\ : InMux
    port map (
            O => \N__33369\,
            I => \N__33365\
        );

    \I__5717\ : CascadeMux
    port map (
            O => \N__33368\,
            I => \N__33362\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__33365\,
            I => \N__33359\
        );

    \I__5715\ : InMux
    port map (
            O => \N__33362\,
            I => \N__33356\
        );

    \I__5714\ : Span4Mux_h
    port map (
            O => \N__33359\,
            I => \N__33353\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__33356\,
            I => \N__33350\
        );

    \I__5712\ : Odrv4
    port map (
            O => \N__33353\,
            I => n2032
        );

    \I__5711\ : Odrv4
    port map (
            O => \N__33350\,
            I => n2032
        );

    \I__5710\ : InMux
    port map (
            O => \N__33345\,
            I => \N__33342\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__33342\,
            I => \N__33338\
        );

    \I__5708\ : CascadeMux
    port map (
            O => \N__33341\,
            I => \N__33335\
        );

    \I__5707\ : Span4Mux_h
    port map (
            O => \N__33338\,
            I => \N__33331\
        );

    \I__5706\ : InMux
    port map (
            O => \N__33335\,
            I => \N__33328\
        );

    \I__5705\ : InMux
    port map (
            O => \N__33334\,
            I => \N__33325\
        );

    \I__5704\ : Odrv4
    port map (
            O => \N__33331\,
            I => n2031
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__33328\,
            I => n2031
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__33325\,
            I => n2031
        );

    \I__5701\ : CascadeMux
    port map (
            O => \N__33318\,
            I => \n2032_cascade_\
        );

    \I__5700\ : CascadeMux
    port map (
            O => \N__33315\,
            I => \N__33311\
        );

    \I__5699\ : CascadeMux
    port map (
            O => \N__33314\,
            I => \N__33308\
        );

    \I__5698\ : InMux
    port map (
            O => \N__33311\,
            I => \N__33304\
        );

    \I__5697\ : InMux
    port map (
            O => \N__33308\,
            I => \N__33301\
        );

    \I__5696\ : InMux
    port map (
            O => \N__33307\,
            I => \N__33298\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__33304\,
            I => n2022
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__33301\,
            I => n2022
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__33298\,
            I => n2022
        );

    \I__5692\ : CascadeMux
    port map (
            O => \N__33291\,
            I => \N__33288\
        );

    \I__5691\ : InMux
    port map (
            O => \N__33288\,
            I => \N__33283\
        );

    \I__5690\ : InMux
    port map (
            O => \N__33287\,
            I => \N__33280\
        );

    \I__5689\ : InMux
    port map (
            O => \N__33286\,
            I => \N__33277\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__33283\,
            I => n2024
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__33280\,
            I => n2024
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__33277\,
            I => n2024
        );

    \I__5685\ : CascadeMux
    port map (
            O => \N__33270\,
            I => \N__33265\
        );

    \I__5684\ : CascadeMux
    port map (
            O => \N__33269\,
            I => \N__33262\
        );

    \I__5683\ : CascadeMux
    port map (
            O => \N__33268\,
            I => \N__33259\
        );

    \I__5682\ : InMux
    port map (
            O => \N__33265\,
            I => \N__33256\
        );

    \I__5681\ : InMux
    port map (
            O => \N__33262\,
            I => \N__33253\
        );

    \I__5680\ : InMux
    port map (
            O => \N__33259\,
            I => \N__33250\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__33256\,
            I => n2023
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__33253\,
            I => n2023
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__33250\,
            I => n2023
        );

    \I__5676\ : InMux
    port map (
            O => \N__33243\,
            I => \N__33240\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__33240\,
            I => n14544
        );

    \I__5674\ : InMux
    port map (
            O => \N__33237\,
            I => \N__33234\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__33234\,
            I => n2087
        );

    \I__5672\ : CascadeMux
    port map (
            O => \N__33231\,
            I => \n2020_cascade_\
        );

    \I__5671\ : InMux
    port map (
            O => \N__33228\,
            I => \N__33224\
        );

    \I__5670\ : InMux
    port map (
            O => \N__33227\,
            I => \N__33221\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__33224\,
            I => \N__33217\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__33221\,
            I => \N__33214\
        );

    \I__5667\ : InMux
    port map (
            O => \N__33220\,
            I => \N__33211\
        );

    \I__5666\ : Span4Mux_h
    port map (
            O => \N__33217\,
            I => \N__33208\
        );

    \I__5665\ : Span4Mux_h
    port map (
            O => \N__33214\,
            I => \N__33205\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__33211\,
            I => \N__33202\
        );

    \I__5663\ : Odrv4
    port map (
            O => \N__33208\,
            I => n2119
        );

    \I__5662\ : Odrv4
    port map (
            O => \N__33205\,
            I => n2119
        );

    \I__5661\ : Odrv4
    port map (
            O => \N__33202\,
            I => n2119
        );

    \I__5660\ : CascadeMux
    port map (
            O => \N__33195\,
            I => \n14446_cascade_\
        );

    \I__5659\ : InMux
    port map (
            O => \N__33192\,
            I => \N__33189\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__33189\,
            I => n11985
        );

    \I__5657\ : CascadeMux
    port map (
            O => \N__33186\,
            I => \n14450_cascade_\
        );

    \I__5656\ : CascadeMux
    port map (
            O => \N__33183\,
            I => \n1950_cascade_\
        );

    \I__5655\ : InMux
    port map (
            O => \N__33180\,
            I => \N__33177\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__33177\,
            I => \N__33172\
        );

    \I__5653\ : InMux
    port map (
            O => \N__33176\,
            I => \N__33167\
        );

    \I__5652\ : InMux
    port map (
            O => \N__33175\,
            I => \N__33167\
        );

    \I__5651\ : Odrv12
    port map (
            O => \N__33172\,
            I => n2017
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__33167\,
            I => n2017
        );

    \I__5649\ : InMux
    port map (
            O => \N__33162\,
            I => \N__33159\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__33159\,
            I => n45_adj_720
        );

    \I__5647\ : InMux
    port map (
            O => \N__33156\,
            I => \N__33153\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__33153\,
            I => \N__33150\
        );

    \I__5645\ : IoSpan4Mux
    port map (
            O => \N__33150\,
            I => \N__33147\
        );

    \I__5644\ : Odrv4
    port map (
            O => \N__33147\,
            I => \ENCODER0_A_N\
        );

    \I__5643\ : CascadeMux
    port map (
            O => \N__33144\,
            I => \n1922_cascade_\
        );

    \I__5642\ : CascadeMux
    port map (
            O => \N__33141\,
            I => \N__33137\
        );

    \I__5641\ : InMux
    port map (
            O => \N__33140\,
            I => \N__33134\
        );

    \I__5640\ : InMux
    port map (
            O => \N__33137\,
            I => \N__33131\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__33134\,
            I => \N__33128\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__33131\,
            I => n2021
        );

    \I__5637\ : Odrv4
    port map (
            O => \N__33128\,
            I => n2021
        );

    \I__5636\ : InMux
    port map (
            O => \N__33123\,
            I => \N__33120\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__33120\,
            I => n2088
        );

    \I__5634\ : CascadeMux
    port map (
            O => \N__33117\,
            I => \n2021_cascade_\
        );

    \I__5633\ : CascadeMux
    port map (
            O => \N__33114\,
            I => \N__33111\
        );

    \I__5632\ : InMux
    port map (
            O => \N__33111\,
            I => \N__33107\
        );

    \I__5631\ : InMux
    port map (
            O => \N__33110\,
            I => \N__33104\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__33107\,
            I => \N__33098\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__33104\,
            I => \N__33098\
        );

    \I__5628\ : InMux
    port map (
            O => \N__33103\,
            I => \N__33095\
        );

    \I__5627\ : Span4Mux_h
    port map (
            O => \N__33098\,
            I => \N__33092\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__33095\,
            I => \N__33089\
        );

    \I__5625\ : Odrv4
    port map (
            O => \N__33092\,
            I => n2120
        );

    \I__5624\ : Odrv12
    port map (
            O => \N__33089\,
            I => n2120
        );

    \I__5623\ : CascadeMux
    port map (
            O => \N__33084\,
            I => \N__33080\
        );

    \I__5622\ : InMux
    port map (
            O => \N__33083\,
            I => \N__33077\
        );

    \I__5621\ : InMux
    port map (
            O => \N__33080\,
            I => \N__33074\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__33077\,
            I => \N__33071\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__33074\,
            I => n2020
        );

    \I__5618\ : Odrv4
    port map (
            O => \N__33071\,
            I => n2020
        );

    \I__5617\ : CascadeMux
    port map (
            O => \N__33066\,
            I => \n14304_cascade_\
        );

    \I__5616\ : CascadeMux
    port map (
            O => \N__33063\,
            I => \n14306_cascade_\
        );

    \I__5615\ : InMux
    port map (
            O => \N__33060\,
            I => \N__33057\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__33057\,
            I => n14308
        );

    \I__5613\ : InMux
    port map (
            O => \N__33054\,
            I => \N__33051\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__33051\,
            I => n5_adj_704
        );

    \I__5611\ : CascadeMux
    port map (
            O => \N__33048\,
            I => \N__33045\
        );

    \I__5610\ : InMux
    port map (
            O => \N__33045\,
            I => \N__33042\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__33042\,
            I => \N__33039\
        );

    \I__5608\ : Odrv4
    port map (
            O => \N__33039\,
            I => n12039
        );

    \I__5607\ : CascadeMux
    port map (
            O => \N__33036\,
            I => \n14292_cascade_\
        );

    \I__5606\ : InMux
    port map (
            O => \N__33033\,
            I => \N__33030\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__33030\,
            I => n14284
        );

    \I__5604\ : CascadeMux
    port map (
            O => \N__33027\,
            I => \n14286_cascade_\
        );

    \I__5603\ : InMux
    port map (
            O => \N__33024\,
            I => \N__33021\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__33021\,
            I => n14288
        );

    \I__5601\ : InMux
    port map (
            O => \N__33018\,
            I => \N__33015\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__33015\,
            I => n14294
        );

    \I__5599\ : CascadeMux
    port map (
            O => \N__33012\,
            I => \n14296_cascade_\
        );

    \I__5598\ : InMux
    port map (
            O => \N__33009\,
            I => \N__33006\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__33006\,
            I => n14298
        );

    \I__5596\ : CascadeMux
    port map (
            O => \N__33003\,
            I => \n29_adj_717_cascade_\
        );

    \I__5595\ : InMux
    port map (
            O => \N__33000\,
            I => \N__32997\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__32997\,
            I => \N__32994\
        );

    \I__5593\ : Span4Mux_h
    port map (
            O => \N__32994\,
            I => \N__32991\
        );

    \I__5592\ : Odrv4
    port map (
            O => \N__32991\,
            I => n14270
        );

    \I__5591\ : CascadeMux
    port map (
            O => \N__32988\,
            I => \n11941_cascade_\
        );

    \I__5590\ : InMux
    port map (
            O => \N__32985\,
            I => \N__32982\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__32982\,
            I => n11878
        );

    \I__5588\ : InMux
    port map (
            O => \N__32979\,
            I => \N__32976\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__32976\,
            I => n14782
        );

    \I__5586\ : InMux
    port map (
            O => \N__32973\,
            I => \N__32970\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__32970\,
            I => n14788
        );

    \I__5584\ : CascadeMux
    port map (
            O => \N__32967\,
            I => \n14300_cascade_\
        );

    \I__5583\ : CascadeMux
    port map (
            O => \N__32964\,
            I => \n14302_cascade_\
        );

    \I__5582\ : InMux
    port map (
            O => \N__32961\,
            I => \N__32958\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__32958\,
            I => \N__32954\
        );

    \I__5580\ : InMux
    port map (
            O => \N__32957\,
            I => \N__32951\
        );

    \I__5579\ : Span4Mux_v
    port map (
            O => \N__32954\,
            I => \N__32946\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__32951\,
            I => \N__32946\
        );

    \I__5577\ : Odrv4
    port map (
            O => \N__32946\,
            I => n3130
        );

    \I__5576\ : CascadeMux
    port map (
            O => \N__32943\,
            I => \N__32940\
        );

    \I__5575\ : InMux
    port map (
            O => \N__32940\,
            I => \N__32937\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__32937\,
            I => \N__32934\
        );

    \I__5573\ : Span4Mux_h
    port map (
            O => \N__32934\,
            I => \N__32931\
        );

    \I__5572\ : Odrv4
    port map (
            O => \N__32931\,
            I => n3197
        );

    \I__5571\ : InMux
    port map (
            O => \N__32928\,
            I => \N__32925\
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__32925\,
            I => \N__32922\
        );

    \I__5569\ : Span4Mux_h
    port map (
            O => \N__32922\,
            I => \N__32919\
        );

    \I__5568\ : Odrv4
    port map (
            O => \N__32919\,
            I => n3193
        );

    \I__5567\ : CascadeMux
    port map (
            O => \N__32916\,
            I => \N__32912\
        );

    \I__5566\ : InMux
    port map (
            O => \N__32915\,
            I => \N__32909\
        );

    \I__5565\ : InMux
    port map (
            O => \N__32912\,
            I => \N__32906\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__32909\,
            I => \N__32902\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__32906\,
            I => \N__32899\
        );

    \I__5562\ : InMux
    port map (
            O => \N__32905\,
            I => \N__32896\
        );

    \I__5561\ : Odrv12
    port map (
            O => \N__32902\,
            I => n3126
        );

    \I__5560\ : Odrv4
    port map (
            O => \N__32899\,
            I => n3126
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__32896\,
            I => n3126
        );

    \I__5558\ : InMux
    port map (
            O => \N__32889\,
            I => \N__32886\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__32886\,
            I => \N__32883\
        );

    \I__5556\ : Span4Mux_v
    port map (
            O => \N__32883\,
            I => \N__32880\
        );

    \I__5555\ : Span4Mux_h
    port map (
            O => \N__32880\,
            I => \N__32877\
        );

    \I__5554\ : Odrv4
    port map (
            O => \N__32877\,
            I => n3201
        );

    \I__5553\ : CascadeMux
    port map (
            O => \N__32874\,
            I => \n3233_cascade_\
        );

    \I__5552\ : CascadeMux
    port map (
            O => \N__32871\,
            I => \n11943_cascade_\
        );

    \I__5551\ : InMux
    port map (
            O => \N__32868\,
            I => \N__32865\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__32865\,
            I => n13875
        );

    \I__5549\ : CascadeMux
    port map (
            O => \N__32862\,
            I => \N__32859\
        );

    \I__5548\ : InMux
    port map (
            O => \N__32859\,
            I => \N__32855\
        );

    \I__5547\ : InMux
    port map (
            O => \N__32858\,
            I => \N__32852\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__32855\,
            I => \N__32849\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__32852\,
            I => n2515
        );

    \I__5544\ : Odrv4
    port map (
            O => \N__32849\,
            I => n2515
        );

    \I__5543\ : InMux
    port map (
            O => \N__32844\,
            I => \N__32841\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__32841\,
            I => \N__32838\
        );

    \I__5541\ : Span4Mux_h
    port map (
            O => \N__32838\,
            I => \N__32835\
        );

    \I__5540\ : Odrv4
    port map (
            O => \N__32835\,
            I => n2582
        );

    \I__5539\ : InMux
    port map (
            O => \N__32832\,
            I => n12757
        );

    \I__5538\ : CascadeMux
    port map (
            O => \N__32829\,
            I => \N__32826\
        );

    \I__5537\ : InMux
    port map (
            O => \N__32826\,
            I => \N__32823\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__32823\,
            I => \N__32819\
        );

    \I__5535\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32815\
        );

    \I__5534\ : Span4Mux_v
    port map (
            O => \N__32819\,
            I => \N__32812\
        );

    \I__5533\ : InMux
    port map (
            O => \N__32818\,
            I => \N__32809\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__32815\,
            I => n2514
        );

    \I__5531\ : Odrv4
    port map (
            O => \N__32812\,
            I => n2514
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__32809\,
            I => n2514
        );

    \I__5529\ : CascadeMux
    port map (
            O => \N__32802\,
            I => \N__32799\
        );

    \I__5528\ : InMux
    port map (
            O => \N__32799\,
            I => \N__32796\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__32796\,
            I => \N__32793\
        );

    \I__5526\ : Span4Mux_v
    port map (
            O => \N__32793\,
            I => \N__32790\
        );

    \I__5525\ : Odrv4
    port map (
            O => \N__32790\,
            I => n2581
        );

    \I__5524\ : InMux
    port map (
            O => \N__32787\,
            I => n12758
        );

    \I__5523\ : CascadeMux
    port map (
            O => \N__32784\,
            I => \N__32781\
        );

    \I__5522\ : InMux
    port map (
            O => \N__32781\,
            I => \N__32777\
        );

    \I__5521\ : InMux
    port map (
            O => \N__32780\,
            I => \N__32774\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__32777\,
            I => n2513
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__32774\,
            I => n2513
        );

    \I__5518\ : InMux
    port map (
            O => \N__32769\,
            I => \N__32766\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__32766\,
            I => n2580
        );

    \I__5516\ : InMux
    port map (
            O => \N__32763\,
            I => n12759
        );

    \I__5515\ : InMux
    port map (
            O => \N__32760\,
            I => n12760
        );

    \I__5514\ : CascadeMux
    port map (
            O => \N__32757\,
            I => \N__32754\
        );

    \I__5513\ : InMux
    port map (
            O => \N__32754\,
            I => \N__32751\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__32751\,
            I => \N__32747\
        );

    \I__5511\ : InMux
    port map (
            O => \N__32750\,
            I => \N__32744\
        );

    \I__5510\ : Odrv12
    port map (
            O => \N__32747\,
            I => n2511
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__32744\,
            I => n2511
        );

    \I__5508\ : InMux
    port map (
            O => \N__32739\,
            I => n12761
        );

    \I__5507\ : CascadeMux
    port map (
            O => \N__32736\,
            I => \N__32733\
        );

    \I__5506\ : InMux
    port map (
            O => \N__32733\,
            I => \N__32729\
        );

    \I__5505\ : InMux
    port map (
            O => \N__32732\,
            I => \N__32726\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__32729\,
            I => \N__32723\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__32726\,
            I => \N__32717\
        );

    \I__5502\ : Span4Mux_v
    port map (
            O => \N__32723\,
            I => \N__32717\
        );

    \I__5501\ : InMux
    port map (
            O => \N__32722\,
            I => \N__32714\
        );

    \I__5500\ : Span4Mux_v
    port map (
            O => \N__32717\,
            I => \N__32709\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__32714\,
            I => \N__32709\
        );

    \I__5498\ : Span4Mux_h
    port map (
            O => \N__32709\,
            I => \N__32706\
        );

    \I__5497\ : Odrv4
    port map (
            O => \N__32706\,
            I => n2610
        );

    \I__5496\ : InMux
    port map (
            O => \N__32703\,
            I => \N__32699\
        );

    \I__5495\ : CascadeMux
    port map (
            O => \N__32702\,
            I => \N__32696\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__32699\,
            I => \N__32692\
        );

    \I__5493\ : InMux
    port map (
            O => \N__32696\,
            I => \N__32689\
        );

    \I__5492\ : InMux
    port map (
            O => \N__32695\,
            I => \N__32686\
        );

    \I__5491\ : Span4Mux_v
    port map (
            O => \N__32692\,
            I => \N__32679\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__32689\,
            I => \N__32679\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__32686\,
            I => \N__32679\
        );

    \I__5488\ : Span4Mux_v
    port map (
            O => \N__32679\,
            I => \N__32676\
        );

    \I__5487\ : Odrv4
    port map (
            O => \N__32676\,
            I => n2418
        );

    \I__5486\ : CascadeMux
    port map (
            O => \N__32673\,
            I => \N__32670\
        );

    \I__5485\ : InMux
    port map (
            O => \N__32670\,
            I => \N__32667\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__32667\,
            I => \N__32664\
        );

    \I__5483\ : Odrv12
    port map (
            O => \N__32664\,
            I => n2485
        );

    \I__5482\ : InMux
    port map (
            O => \N__32661\,
            I => \N__32658\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__32658\,
            I => \N__32654\
        );

    \I__5480\ : CascadeMux
    port map (
            O => \N__32657\,
            I => \N__32651\
        );

    \I__5479\ : Span4Mux_v
    port map (
            O => \N__32654\,
            I => \N__32648\
        );

    \I__5478\ : InMux
    port map (
            O => \N__32651\,
            I => \N__32645\
        );

    \I__5477\ : Span4Mux_v
    port map (
            O => \N__32648\,
            I => \N__32642\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__32645\,
            I => n2517
        );

    \I__5475\ : Odrv4
    port map (
            O => \N__32642\,
            I => n2517
        );

    \I__5474\ : InMux
    port map (
            O => \N__32637\,
            I => \N__32634\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__32634\,
            I => n2584
        );

    \I__5472\ : CascadeMux
    port map (
            O => \N__32631\,
            I => \n2517_cascade_\
        );

    \I__5471\ : InMux
    port map (
            O => \N__32628\,
            I => \N__32625\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__32625\,
            I => \N__32621\
        );

    \I__5469\ : InMux
    port map (
            O => \N__32624\,
            I => \N__32618\
        );

    \I__5468\ : Span4Mux_h
    port map (
            O => \N__32621\,
            I => \N__32614\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__32618\,
            I => \N__32611\
        );

    \I__5466\ : InMux
    port map (
            O => \N__32617\,
            I => \N__32608\
        );

    \I__5465\ : Span4Mux_v
    port map (
            O => \N__32614\,
            I => \N__32605\
        );

    \I__5464\ : Span4Mux_v
    port map (
            O => \N__32611\,
            I => \N__32600\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__32608\,
            I => \N__32600\
        );

    \I__5462\ : Span4Mux_v
    port map (
            O => \N__32605\,
            I => \N__32595\
        );

    \I__5461\ : Span4Mux_h
    port map (
            O => \N__32600\,
            I => \N__32595\
        );

    \I__5460\ : Odrv4
    port map (
            O => \N__32595\,
            I => n2616
        );

    \I__5459\ : InMux
    port map (
            O => \N__32592\,
            I => \N__32588\
        );

    \I__5458\ : InMux
    port map (
            O => \N__32591\,
            I => \N__32585\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__32588\,
            I => \N__32580\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__32585\,
            I => \N__32580\
        );

    \I__5455\ : Span4Mux_v
    port map (
            O => \N__32580\,
            I => \N__32576\
        );

    \I__5454\ : InMux
    port map (
            O => \N__32579\,
            I => \N__32573\
        );

    \I__5453\ : Odrv4
    port map (
            O => \N__32576\,
            I => n2512
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__32573\,
            I => n2512
        );

    \I__5451\ : CascadeMux
    port map (
            O => \N__32568\,
            I => \N__32565\
        );

    \I__5450\ : InMux
    port map (
            O => \N__32565\,
            I => \N__32562\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__32562\,
            I => n2579
        );

    \I__5448\ : InMux
    port map (
            O => \N__32559\,
            I => \N__32556\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__32556\,
            I => \N__32552\
        );

    \I__5446\ : InMux
    port map (
            O => \N__32555\,
            I => \N__32549\
        );

    \I__5445\ : Span4Mux_h
    port map (
            O => \N__32552\,
            I => \N__32545\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__32549\,
            I => \N__32542\
        );

    \I__5443\ : InMux
    port map (
            O => \N__32548\,
            I => \N__32539\
        );

    \I__5442\ : Span4Mux_v
    port map (
            O => \N__32545\,
            I => \N__32536\
        );

    \I__5441\ : Span4Mux_v
    port map (
            O => \N__32542\,
            I => \N__32531\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__32539\,
            I => \N__32531\
        );

    \I__5439\ : Span4Mux_v
    port map (
            O => \N__32536\,
            I => \N__32526\
        );

    \I__5438\ : Span4Mux_h
    port map (
            O => \N__32531\,
            I => \N__32526\
        );

    \I__5437\ : Odrv4
    port map (
            O => \N__32526\,
            I => n2611
        );

    \I__5436\ : InMux
    port map (
            O => \N__32523\,
            I => n12748
        );

    \I__5435\ : CascadeMux
    port map (
            O => \N__32520\,
            I => \N__32517\
        );

    \I__5434\ : InMux
    port map (
            O => \N__32517\,
            I => \N__32514\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__32514\,
            I => \N__32510\
        );

    \I__5432\ : InMux
    port map (
            O => \N__32513\,
            I => \N__32507\
        );

    \I__5431\ : Span4Mux_h
    port map (
            O => \N__32510\,
            I => \N__32504\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__32507\,
            I => n2523
        );

    \I__5429\ : Odrv4
    port map (
            O => \N__32504\,
            I => n2523
        );

    \I__5428\ : InMux
    port map (
            O => \N__32499\,
            I => \N__32496\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__32496\,
            I => \N__32493\
        );

    \I__5426\ : Span4Mux_h
    port map (
            O => \N__32493\,
            I => \N__32490\
        );

    \I__5425\ : Odrv4
    port map (
            O => \N__32490\,
            I => n2590
        );

    \I__5424\ : InMux
    port map (
            O => \N__32487\,
            I => n12749
        );

    \I__5423\ : CascadeMux
    port map (
            O => \N__32484\,
            I => \N__32481\
        );

    \I__5422\ : InMux
    port map (
            O => \N__32481\,
            I => \N__32478\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__32478\,
            I => \N__32475\
        );

    \I__5420\ : Span4Mux_h
    port map (
            O => \N__32475\,
            I => \N__32472\
        );

    \I__5419\ : Odrv4
    port map (
            O => \N__32472\,
            I => n2589
        );

    \I__5418\ : InMux
    port map (
            O => \N__32469\,
            I => n12750
        );

    \I__5417\ : InMux
    port map (
            O => \N__32466\,
            I => \N__32463\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__32463\,
            I => \N__32460\
        );

    \I__5415\ : Odrv4
    port map (
            O => \N__32460\,
            I => n2588
        );

    \I__5414\ : InMux
    port map (
            O => \N__32457\,
            I => n12751
        );

    \I__5413\ : CascadeMux
    port map (
            O => \N__32454\,
            I => \N__32451\
        );

    \I__5412\ : InMux
    port map (
            O => \N__32451\,
            I => \N__32447\
        );

    \I__5411\ : InMux
    port map (
            O => \N__32450\,
            I => \N__32443\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__32447\,
            I => \N__32440\
        );

    \I__5409\ : InMux
    port map (
            O => \N__32446\,
            I => \N__32437\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__32443\,
            I => n2520
        );

    \I__5407\ : Odrv4
    port map (
            O => \N__32440\,
            I => n2520
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__32437\,
            I => n2520
        );

    \I__5405\ : InMux
    port map (
            O => \N__32430\,
            I => \N__32427\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__32427\,
            I => \N__32424\
        );

    \I__5403\ : Span4Mux_h
    port map (
            O => \N__32424\,
            I => \N__32421\
        );

    \I__5402\ : Odrv4
    port map (
            O => \N__32421\,
            I => n2587
        );

    \I__5401\ : InMux
    port map (
            O => \N__32418\,
            I => n12752
        );

    \I__5400\ : CascadeMux
    port map (
            O => \N__32415\,
            I => \N__32412\
        );

    \I__5399\ : InMux
    port map (
            O => \N__32412\,
            I => \N__32409\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__32409\,
            I => \N__32405\
        );

    \I__5397\ : InMux
    port map (
            O => \N__32408\,
            I => \N__32401\
        );

    \I__5396\ : Span4Mux_v
    port map (
            O => \N__32405\,
            I => \N__32398\
        );

    \I__5395\ : InMux
    port map (
            O => \N__32404\,
            I => \N__32395\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__32401\,
            I => n2519
        );

    \I__5393\ : Odrv4
    port map (
            O => \N__32398\,
            I => n2519
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__32395\,
            I => n2519
        );

    \I__5391\ : CascadeMux
    port map (
            O => \N__32388\,
            I => \N__32385\
        );

    \I__5390\ : InMux
    port map (
            O => \N__32385\,
            I => \N__32382\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__32382\,
            I => \N__32379\
        );

    \I__5388\ : Span4Mux_v
    port map (
            O => \N__32379\,
            I => \N__32376\
        );

    \I__5387\ : Odrv4
    port map (
            O => \N__32376\,
            I => n2586
        );

    \I__5386\ : InMux
    port map (
            O => \N__32373\,
            I => n12753
        );

    \I__5385\ : CascadeMux
    port map (
            O => \N__32370\,
            I => \N__32367\
        );

    \I__5384\ : InMux
    port map (
            O => \N__32367\,
            I => \N__32364\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__32364\,
            I => \N__32361\
        );

    \I__5382\ : Span4Mux_h
    port map (
            O => \N__32361\,
            I => \N__32358\
        );

    \I__5381\ : Odrv4
    port map (
            O => \N__32358\,
            I => n2585
        );

    \I__5380\ : InMux
    port map (
            O => \N__32355\,
            I => \bfn_6_26_0_\
        );

    \I__5379\ : InMux
    port map (
            O => \N__32352\,
            I => n12755
        );

    \I__5378\ : InMux
    port map (
            O => \N__32349\,
            I => \N__32345\
        );

    \I__5377\ : CascadeMux
    port map (
            O => \N__32348\,
            I => \N__32342\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__32345\,
            I => \N__32339\
        );

    \I__5375\ : InMux
    port map (
            O => \N__32342\,
            I => \N__32336\
        );

    \I__5374\ : Span4Mux_v
    port map (
            O => \N__32339\,
            I => \N__32331\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__32336\,
            I => \N__32331\
        );

    \I__5372\ : Span4Mux_v
    port map (
            O => \N__32331\,
            I => \N__32327\
        );

    \I__5371\ : InMux
    port map (
            O => \N__32330\,
            I => \N__32324\
        );

    \I__5370\ : Odrv4
    port map (
            O => \N__32327\,
            I => n2516
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__32324\,
            I => n2516
        );

    \I__5368\ : InMux
    port map (
            O => \N__32319\,
            I => \N__32316\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__32316\,
            I => n2583
        );

    \I__5366\ : InMux
    port map (
            O => \N__32313\,
            I => n12756
        );

    \I__5365\ : CascadeMux
    port map (
            O => \N__32310\,
            I => \N__32307\
        );

    \I__5364\ : InMux
    port map (
            O => \N__32307\,
            I => \N__32302\
        );

    \I__5363\ : InMux
    port map (
            O => \N__32306\,
            I => \N__32299\
        );

    \I__5362\ : InMux
    port map (
            O => \N__32305\,
            I => \N__32296\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__32302\,
            I => \N__32293\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__32299\,
            I => \N__32288\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__32296\,
            I => \N__32288\
        );

    \I__5358\ : Odrv4
    port map (
            O => \N__32293\,
            I => n2531
        );

    \I__5357\ : Odrv4
    port map (
            O => \N__32288\,
            I => n2531
        );

    \I__5356\ : InMux
    port map (
            O => \N__32283\,
            I => \N__32280\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__32280\,
            I => n2598
        );

    \I__5354\ : InMux
    port map (
            O => \N__32277\,
            I => n12741
        );

    \I__5353\ : CascadeMux
    port map (
            O => \N__32274\,
            I => \N__32271\
        );

    \I__5352\ : InMux
    port map (
            O => \N__32271\,
            I => \N__32267\
        );

    \I__5351\ : CascadeMux
    port map (
            O => \N__32270\,
            I => \N__32264\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__32267\,
            I => \N__32261\
        );

    \I__5349\ : InMux
    port map (
            O => \N__32264\,
            I => \N__32258\
        );

    \I__5348\ : Odrv4
    port map (
            O => \N__32261\,
            I => n2530
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__32258\,
            I => n2530
        );

    \I__5346\ : InMux
    port map (
            O => \N__32253\,
            I => \N__32250\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__32250\,
            I => n2597
        );

    \I__5344\ : InMux
    port map (
            O => \N__32247\,
            I => n12742
        );

    \I__5343\ : InMux
    port map (
            O => \N__32244\,
            I => \N__32241\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__32241\,
            I => \N__32237\
        );

    \I__5341\ : CascadeMux
    port map (
            O => \N__32240\,
            I => \N__32234\
        );

    \I__5340\ : Span4Mux_h
    port map (
            O => \N__32237\,
            I => \N__32230\
        );

    \I__5339\ : InMux
    port map (
            O => \N__32234\,
            I => \N__32227\
        );

    \I__5338\ : InMux
    port map (
            O => \N__32233\,
            I => \N__32224\
        );

    \I__5337\ : Odrv4
    port map (
            O => \N__32230\,
            I => n2529
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__32227\,
            I => n2529
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__32224\,
            I => n2529
        );

    \I__5334\ : CascadeMux
    port map (
            O => \N__32217\,
            I => \N__32214\
        );

    \I__5333\ : InMux
    port map (
            O => \N__32214\,
            I => \N__32211\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__32211\,
            I => \N__32208\
        );

    \I__5331\ : Span4Mux_v
    port map (
            O => \N__32208\,
            I => \N__32205\
        );

    \I__5330\ : Odrv4
    port map (
            O => \N__32205\,
            I => n2596
        );

    \I__5329\ : InMux
    port map (
            O => \N__32202\,
            I => n12743
        );

    \I__5328\ : CascadeMux
    port map (
            O => \N__32199\,
            I => \N__32196\
        );

    \I__5327\ : InMux
    port map (
            O => \N__32196\,
            I => \N__32193\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__32193\,
            I => \N__32190\
        );

    \I__5325\ : Span4Mux_h
    port map (
            O => \N__32190\,
            I => \N__32186\
        );

    \I__5324\ : InMux
    port map (
            O => \N__32189\,
            I => \N__32183\
        );

    \I__5323\ : Odrv4
    port map (
            O => \N__32186\,
            I => n2528
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__32183\,
            I => n2528
        );

    \I__5321\ : InMux
    port map (
            O => \N__32178\,
            I => \N__32175\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__32175\,
            I => \N__32172\
        );

    \I__5319\ : Odrv4
    port map (
            O => \N__32172\,
            I => n2595
        );

    \I__5318\ : InMux
    port map (
            O => \N__32169\,
            I => n12744
        );

    \I__5317\ : CascadeMux
    port map (
            O => \N__32166\,
            I => \N__32163\
        );

    \I__5316\ : InMux
    port map (
            O => \N__32163\,
            I => \N__32160\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__32160\,
            I => \N__32157\
        );

    \I__5314\ : Span4Mux_h
    port map (
            O => \N__32157\,
            I => \N__32153\
        );

    \I__5313\ : InMux
    port map (
            O => \N__32156\,
            I => \N__32150\
        );

    \I__5312\ : Odrv4
    port map (
            O => \N__32153\,
            I => n2527
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__32150\,
            I => n2527
        );

    \I__5310\ : InMux
    port map (
            O => \N__32145\,
            I => \N__32142\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__32142\,
            I => \N__32139\
        );

    \I__5308\ : Span4Mux_h
    port map (
            O => \N__32139\,
            I => \N__32136\
        );

    \I__5307\ : Odrv4
    port map (
            O => \N__32136\,
            I => n2594
        );

    \I__5306\ : InMux
    port map (
            O => \N__32133\,
            I => n12745
        );

    \I__5305\ : CascadeMux
    port map (
            O => \N__32130\,
            I => \N__32127\
        );

    \I__5304\ : InMux
    port map (
            O => \N__32127\,
            I => \N__32124\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__32124\,
            I => \N__32121\
        );

    \I__5302\ : Span4Mux_v
    port map (
            O => \N__32121\,
            I => \N__32117\
        );

    \I__5301\ : InMux
    port map (
            O => \N__32120\,
            I => \N__32114\
        );

    \I__5300\ : Odrv4
    port map (
            O => \N__32117\,
            I => n2526
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__32114\,
            I => n2526
        );

    \I__5298\ : InMux
    port map (
            O => \N__32109\,
            I => \N__32106\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__32106\,
            I => \N__32103\
        );

    \I__5296\ : Span4Mux_h
    port map (
            O => \N__32103\,
            I => \N__32100\
        );

    \I__5295\ : Odrv4
    port map (
            O => \N__32100\,
            I => n2593
        );

    \I__5294\ : InMux
    port map (
            O => \N__32097\,
            I => \bfn_6_25_0_\
        );

    \I__5293\ : InMux
    port map (
            O => \N__32094\,
            I => n12747
        );

    \I__5292\ : InMux
    port map (
            O => \N__32091\,
            I => \N__32087\
        );

    \I__5291\ : CascadeMux
    port map (
            O => \N__32090\,
            I => \N__32084\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__32087\,
            I => \N__32081\
        );

    \I__5289\ : InMux
    port map (
            O => \N__32084\,
            I => \N__32078\
        );

    \I__5288\ : Span4Mux_v
    port map (
            O => \N__32081\,
            I => \N__32075\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__32078\,
            I => n2524
        );

    \I__5286\ : Odrv4
    port map (
            O => \N__32075\,
            I => n2524
        );

    \I__5285\ : InMux
    port map (
            O => \N__32070\,
            I => \N__32067\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__32067\,
            I => \N__32064\
        );

    \I__5283\ : Span4Mux_h
    port map (
            O => \N__32064\,
            I => \N__32061\
        );

    \I__5282\ : Odrv4
    port map (
            O => \N__32061\,
            I => n2591
        );

    \I__5281\ : InMux
    port map (
            O => \N__32058\,
            I => n12734
        );

    \I__5280\ : CascadeMux
    port map (
            O => \N__32055\,
            I => \N__32050\
        );

    \I__5279\ : InMux
    port map (
            O => \N__32054\,
            I => \N__32047\
        );

    \I__5278\ : InMux
    port map (
            O => \N__32053\,
            I => \N__32042\
        );

    \I__5277\ : InMux
    port map (
            O => \N__32050\,
            I => \N__32042\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__32047\,
            I => \N__32037\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__32042\,
            I => \N__32037\
        );

    \I__5274\ : Span4Mux_h
    port map (
            O => \N__32037\,
            I => \N__32034\
        );

    \I__5273\ : Odrv4
    port map (
            O => \N__32034\,
            I => n2415
        );

    \I__5272\ : InMux
    port map (
            O => \N__32031\,
            I => \N__32028\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__32028\,
            I => n2482
        );

    \I__5270\ : InMux
    port map (
            O => \N__32025\,
            I => n12735
        );

    \I__5269\ : CascadeMux
    port map (
            O => \N__32022\,
            I => \N__32019\
        );

    \I__5268\ : InMux
    port map (
            O => \N__32019\,
            I => \N__32016\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__32016\,
            I => \N__32012\
        );

    \I__5266\ : InMux
    port map (
            O => \N__32015\,
            I => \N__32009\
        );

    \I__5265\ : Span4Mux_v
    port map (
            O => \N__32012\,
            I => \N__32003\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__32009\,
            I => \N__32003\
        );

    \I__5263\ : InMux
    port map (
            O => \N__32008\,
            I => \N__32000\
        );

    \I__5262\ : Span4Mux_h
    port map (
            O => \N__32003\,
            I => \N__31995\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__32000\,
            I => \N__31995\
        );

    \I__5260\ : Odrv4
    port map (
            O => \N__31995\,
            I => n2414
        );

    \I__5259\ : InMux
    port map (
            O => \N__31992\,
            I => \N__31989\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__31989\,
            I => \N__31986\
        );

    \I__5257\ : Odrv4
    port map (
            O => \N__31986\,
            I => n2481
        );

    \I__5256\ : InMux
    port map (
            O => \N__31983\,
            I => n12736
        );

    \I__5255\ : InMux
    port map (
            O => \N__31980\,
            I => \N__31976\
        );

    \I__5254\ : InMux
    port map (
            O => \N__31979\,
            I => \N__31973\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__31976\,
            I => \N__31969\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__31973\,
            I => \N__31966\
        );

    \I__5251\ : InMux
    port map (
            O => \N__31972\,
            I => \N__31963\
        );

    \I__5250\ : Span4Mux_v
    port map (
            O => \N__31969\,
            I => \N__31956\
        );

    \I__5249\ : Span4Mux_h
    port map (
            O => \N__31966\,
            I => \N__31956\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__31963\,
            I => \N__31956\
        );

    \I__5247\ : Odrv4
    port map (
            O => \N__31956\,
            I => n2413
        );

    \I__5246\ : InMux
    port map (
            O => \N__31953\,
            I => \N__31950\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__31950\,
            I => n2480
        );

    \I__5244\ : InMux
    port map (
            O => \N__31947\,
            I => n12737
        );

    \I__5243\ : InMux
    port map (
            O => \N__31944\,
            I => \N__31941\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__31941\,
            I => \N__31937\
        );

    \I__5241\ : InMux
    port map (
            O => \N__31940\,
            I => \N__31934\
        );

    \I__5240\ : Span4Mux_h
    port map (
            O => \N__31937\,
            I => \N__31929\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__31934\,
            I => \N__31929\
        );

    \I__5238\ : Span4Mux_h
    port map (
            O => \N__31929\,
            I => \N__31926\
        );

    \I__5237\ : Odrv4
    port map (
            O => \N__31926\,
            I => n2412
        );

    \I__5236\ : InMux
    port map (
            O => \N__31923\,
            I => n12738
        );

    \I__5235\ : InMux
    port map (
            O => \N__31920\,
            I => \N__31917\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__31917\,
            I => \N__31913\
        );

    \I__5233\ : CascadeMux
    port map (
            O => \N__31916\,
            I => \N__31910\
        );

    \I__5232\ : Span4Mux_v
    port map (
            O => \N__31913\,
            I => \N__31906\
        );

    \I__5231\ : InMux
    port map (
            O => \N__31910\,
            I => \N__31903\
        );

    \I__5230\ : InMux
    port map (
            O => \N__31909\,
            I => \N__31900\
        );

    \I__5229\ : Odrv4
    port map (
            O => \N__31906\,
            I => n2433
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__31903\,
            I => n2433
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__31900\,
            I => n2433
        );

    \I__5226\ : CascadeMux
    port map (
            O => \N__31893\,
            I => \N__31890\
        );

    \I__5225\ : InMux
    port map (
            O => \N__31890\,
            I => \N__31887\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__31887\,
            I => \N__31884\
        );

    \I__5223\ : Odrv4
    port map (
            O => \N__31884\,
            I => n2500
        );

    \I__5222\ : InMux
    port map (
            O => \N__31881\,
            I => \N__31878\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__31878\,
            I => \N__31875\
        );

    \I__5220\ : Span4Mux_v
    port map (
            O => \N__31875\,
            I => \N__31872\
        );

    \I__5219\ : Odrv4
    port map (
            O => \N__31872\,
            I => n2601
        );

    \I__5218\ : InMux
    port map (
            O => \N__31869\,
            I => \bfn_6_24_0_\
        );

    \I__5217\ : CascadeMux
    port map (
            O => \N__31866\,
            I => \N__31862\
        );

    \I__5216\ : InMux
    port map (
            O => \N__31865\,
            I => \N__31859\
        );

    \I__5215\ : InMux
    port map (
            O => \N__31862\,
            I => \N__31856\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__31859\,
            I => n2533
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__31856\,
            I => n2533
        );

    \I__5212\ : CascadeMux
    port map (
            O => \N__31851\,
            I => \N__31848\
        );

    \I__5211\ : InMux
    port map (
            O => \N__31848\,
            I => \N__31845\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__31845\,
            I => n2600
        );

    \I__5209\ : InMux
    port map (
            O => \N__31842\,
            I => n12739
        );

    \I__5208\ : CascadeMux
    port map (
            O => \N__31839\,
            I => \N__31836\
        );

    \I__5207\ : InMux
    port map (
            O => \N__31836\,
            I => \N__31831\
        );

    \I__5206\ : InMux
    port map (
            O => \N__31835\,
            I => \N__31826\
        );

    \I__5205\ : InMux
    port map (
            O => \N__31834\,
            I => \N__31826\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__31831\,
            I => n2532
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__31826\,
            I => n2532
        );

    \I__5202\ : InMux
    port map (
            O => \N__31821\,
            I => \N__31818\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__31818\,
            I => n2599
        );

    \I__5200\ : InMux
    port map (
            O => \N__31815\,
            I => n12740
        );

    \I__5199\ : CascadeMux
    port map (
            O => \N__31812\,
            I => \N__31809\
        );

    \I__5198\ : InMux
    port map (
            O => \N__31809\,
            I => \N__31805\
        );

    \I__5197\ : InMux
    port map (
            O => \N__31808\,
            I => \N__31802\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__31805\,
            I => \N__31799\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__31802\,
            I => \N__31793\
        );

    \I__5194\ : Span4Mux_h
    port map (
            O => \N__31799\,
            I => \N__31793\
        );

    \I__5193\ : InMux
    port map (
            O => \N__31798\,
            I => \N__31790\
        );

    \I__5192\ : Odrv4
    port map (
            O => \N__31793\,
            I => n2424
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__31790\,
            I => n2424
        );

    \I__5190\ : CascadeMux
    port map (
            O => \N__31785\,
            I => \N__31782\
        );

    \I__5189\ : InMux
    port map (
            O => \N__31782\,
            I => \N__31779\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__31779\,
            I => \N__31776\
        );

    \I__5187\ : Odrv4
    port map (
            O => \N__31776\,
            I => n2491
        );

    \I__5186\ : InMux
    port map (
            O => \N__31773\,
            I => n12726
        );

    \I__5185\ : InMux
    port map (
            O => \N__31770\,
            I => n12727
        );

    \I__5184\ : InMux
    port map (
            O => \N__31767\,
            I => n12728
        );

    \I__5183\ : CascadeMux
    port map (
            O => \N__31764\,
            I => \N__31761\
        );

    \I__5182\ : InMux
    port map (
            O => \N__31761\,
            I => \N__31757\
        );

    \I__5181\ : InMux
    port map (
            O => \N__31760\,
            I => \N__31754\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__31757\,
            I => \N__31750\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__31754\,
            I => \N__31747\
        );

    \I__5178\ : InMux
    port map (
            O => \N__31753\,
            I => \N__31744\
        );

    \I__5177\ : Odrv12
    port map (
            O => \N__31750\,
            I => n2421
        );

    \I__5176\ : Odrv4
    port map (
            O => \N__31747\,
            I => n2421
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__31744\,
            I => n2421
        );

    \I__5174\ : InMux
    port map (
            O => \N__31737\,
            I => \N__31734\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__31734\,
            I => n2488
        );

    \I__5172\ : InMux
    port map (
            O => \N__31731\,
            I => n12729
        );

    \I__5171\ : CascadeMux
    port map (
            O => \N__31728\,
            I => \N__31724\
        );

    \I__5170\ : CascadeMux
    port map (
            O => \N__31727\,
            I => \N__31721\
        );

    \I__5169\ : InMux
    port map (
            O => \N__31724\,
            I => \N__31718\
        );

    \I__5168\ : InMux
    port map (
            O => \N__31721\,
            I => \N__31715\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__31718\,
            I => n2420
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__31715\,
            I => n2420
        );

    \I__5165\ : InMux
    port map (
            O => \N__31710\,
            I => \N__31707\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__31707\,
            I => \N__31704\
        );

    \I__5163\ : Odrv4
    port map (
            O => \N__31704\,
            I => n2487
        );

    \I__5162\ : InMux
    port map (
            O => \N__31701\,
            I => n12730
        );

    \I__5161\ : InMux
    port map (
            O => \N__31698\,
            I => n12731
        );

    \I__5160\ : InMux
    port map (
            O => \N__31695\,
            I => \bfn_6_23_0_\
        );

    \I__5159\ : InMux
    port map (
            O => \N__31692\,
            I => \N__31688\
        );

    \I__5158\ : InMux
    port map (
            O => \N__31691\,
            I => \N__31685\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__31688\,
            I => n2417
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__31685\,
            I => n2417
        );

    \I__5155\ : InMux
    port map (
            O => \N__31680\,
            I => \N__31677\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__31677\,
            I => n2484
        );

    \I__5153\ : InMux
    port map (
            O => \N__31674\,
            I => n12733
        );

    \I__5152\ : InMux
    port map (
            O => \N__31671\,
            I => \N__31668\
        );

    \I__5151\ : LocalMux
    port map (
            O => \N__31668\,
            I => \N__31663\
        );

    \I__5150\ : InMux
    port map (
            O => \N__31667\,
            I => \N__31660\
        );

    \I__5149\ : InMux
    port map (
            O => \N__31666\,
            I => \N__31657\
        );

    \I__5148\ : Odrv4
    port map (
            O => \N__31663\,
            I => n2416
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__31660\,
            I => n2416
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__31657\,
            I => n2416
        );

    \I__5145\ : CascadeMux
    port map (
            O => \N__31650\,
            I => \N__31647\
        );

    \I__5144\ : InMux
    port map (
            O => \N__31647\,
            I => \N__31644\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__31644\,
            I => n2483
        );

    \I__5142\ : CascadeMux
    port map (
            O => \N__31641\,
            I => \N__31637\
        );

    \I__5141\ : CascadeMux
    port map (
            O => \N__31640\,
            I => \N__31634\
        );

    \I__5140\ : InMux
    port map (
            O => \N__31637\,
            I => \N__31631\
        );

    \I__5139\ : InMux
    port map (
            O => \N__31634\,
            I => \N__31628\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__31631\,
            I => n2432
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__31628\,
            I => n2432
        );

    \I__5136\ : InMux
    port map (
            O => \N__31623\,
            I => \N__31620\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__31620\,
            I => \N__31617\
        );

    \I__5134\ : Odrv4
    port map (
            O => \N__31617\,
            I => n2499
        );

    \I__5133\ : InMux
    port map (
            O => \N__31614\,
            I => n12718
        );

    \I__5132\ : InMux
    port map (
            O => \N__31611\,
            I => \N__31607\
        );

    \I__5131\ : CascadeMux
    port map (
            O => \N__31610\,
            I => \N__31603\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__31607\,
            I => \N__31600\
        );

    \I__5129\ : InMux
    port map (
            O => \N__31606\,
            I => \N__31597\
        );

    \I__5128\ : InMux
    port map (
            O => \N__31603\,
            I => \N__31594\
        );

    \I__5127\ : Odrv4
    port map (
            O => \N__31600\,
            I => n2431
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__31597\,
            I => n2431
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__31594\,
            I => n2431
        );

    \I__5124\ : CascadeMux
    port map (
            O => \N__31587\,
            I => \N__31584\
        );

    \I__5123\ : InMux
    port map (
            O => \N__31584\,
            I => \N__31581\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__31581\,
            I => \N__31578\
        );

    \I__5121\ : Odrv4
    port map (
            O => \N__31578\,
            I => n2498
        );

    \I__5120\ : InMux
    port map (
            O => \N__31575\,
            I => n12719
        );

    \I__5119\ : InMux
    port map (
            O => \N__31572\,
            I => \N__31568\
        );

    \I__5118\ : CascadeMux
    port map (
            O => \N__31571\,
            I => \N__31565\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__31568\,
            I => \N__31562\
        );

    \I__5116\ : InMux
    port map (
            O => \N__31565\,
            I => \N__31559\
        );

    \I__5115\ : Odrv12
    port map (
            O => \N__31562\,
            I => n2430
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__31559\,
            I => n2430
        );

    \I__5113\ : InMux
    port map (
            O => \N__31554\,
            I => \N__31551\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__31551\,
            I => \N__31548\
        );

    \I__5111\ : Odrv4
    port map (
            O => \N__31548\,
            I => n2497
        );

    \I__5110\ : InMux
    port map (
            O => \N__31545\,
            I => n12720
        );

    \I__5109\ : CascadeMux
    port map (
            O => \N__31542\,
            I => \N__31539\
        );

    \I__5108\ : InMux
    port map (
            O => \N__31539\,
            I => \N__31535\
        );

    \I__5107\ : CascadeMux
    port map (
            O => \N__31538\,
            I => \N__31532\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__31535\,
            I => \N__31528\
        );

    \I__5105\ : InMux
    port map (
            O => \N__31532\,
            I => \N__31525\
        );

    \I__5104\ : InMux
    port map (
            O => \N__31531\,
            I => \N__31522\
        );

    \I__5103\ : Odrv4
    port map (
            O => \N__31528\,
            I => n2429
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__31525\,
            I => n2429
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__31522\,
            I => n2429
        );

    \I__5100\ : InMux
    port map (
            O => \N__31515\,
            I => \N__31512\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__31512\,
            I => n2496
        );

    \I__5098\ : InMux
    port map (
            O => \N__31509\,
            I => n12721
        );

    \I__5097\ : CascadeMux
    port map (
            O => \N__31506\,
            I => \N__31503\
        );

    \I__5096\ : InMux
    port map (
            O => \N__31503\,
            I => \N__31499\
        );

    \I__5095\ : InMux
    port map (
            O => \N__31502\,
            I => \N__31495\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__31499\,
            I => \N__31492\
        );

    \I__5093\ : InMux
    port map (
            O => \N__31498\,
            I => \N__31489\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__31495\,
            I => n2428
        );

    \I__5091\ : Odrv4
    port map (
            O => \N__31492\,
            I => n2428
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__31489\,
            I => n2428
        );

    \I__5089\ : CascadeMux
    port map (
            O => \N__31482\,
            I => \N__31479\
        );

    \I__5088\ : InMux
    port map (
            O => \N__31479\,
            I => \N__31476\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__31476\,
            I => \N__31473\
        );

    \I__5086\ : Span4Mux_h
    port map (
            O => \N__31473\,
            I => \N__31470\
        );

    \I__5085\ : Odrv4
    port map (
            O => \N__31470\,
            I => n2495
        );

    \I__5084\ : InMux
    port map (
            O => \N__31467\,
            I => n12722
        );

    \I__5083\ : InMux
    port map (
            O => \N__31464\,
            I => \N__31460\
        );

    \I__5082\ : InMux
    port map (
            O => \N__31463\,
            I => \N__31457\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__31460\,
            I => \N__31452\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__31457\,
            I => \N__31452\
        );

    \I__5079\ : Odrv4
    port map (
            O => \N__31452\,
            I => n2427
        );

    \I__5078\ : CascadeMux
    port map (
            O => \N__31449\,
            I => \N__31446\
        );

    \I__5077\ : InMux
    port map (
            O => \N__31446\,
            I => \N__31443\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__31443\,
            I => \N__31440\
        );

    \I__5075\ : Odrv4
    port map (
            O => \N__31440\,
            I => n2494
        );

    \I__5074\ : InMux
    port map (
            O => \N__31437\,
            I => n12723
        );

    \I__5073\ : InMux
    port map (
            O => \N__31434\,
            I => \bfn_6_22_0_\
        );

    \I__5072\ : CascadeMux
    port map (
            O => \N__31431\,
            I => \N__31427\
        );

    \I__5071\ : InMux
    port map (
            O => \N__31430\,
            I => \N__31424\
        );

    \I__5070\ : InMux
    port map (
            O => \N__31427\,
            I => \N__31421\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__31424\,
            I => \N__31417\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__31421\,
            I => \N__31414\
        );

    \I__5067\ : InMux
    port map (
            O => \N__31420\,
            I => \N__31411\
        );

    \I__5066\ : Odrv4
    port map (
            O => \N__31417\,
            I => n2425
        );

    \I__5065\ : Odrv4
    port map (
            O => \N__31414\,
            I => n2425
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__31411\,
            I => n2425
        );

    \I__5063\ : InMux
    port map (
            O => \N__31404\,
            I => \N__31401\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__31401\,
            I => \N__31398\
        );

    \I__5061\ : Odrv4
    port map (
            O => \N__31398\,
            I => n2492
        );

    \I__5060\ : InMux
    port map (
            O => \N__31395\,
            I => n12725
        );

    \I__5059\ : CascadeMux
    port map (
            O => \N__31392\,
            I => \n14558_cascade_\
        );

    \I__5058\ : InMux
    port map (
            O => \N__31389\,
            I => \N__31386\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__31386\,
            I => \N__31383\
        );

    \I__5056\ : Odrv4
    port map (
            O => \N__31383\,
            I => n2101
        );

    \I__5055\ : CascadeMux
    port map (
            O => \N__31380\,
            I => \n2049_cascade_\
        );

    \I__5054\ : InMux
    port map (
            O => \N__31377\,
            I => \N__31371\
        );

    \I__5053\ : InMux
    port map (
            O => \N__31376\,
            I => \N__31371\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__31371\,
            I => \N__31368\
        );

    \I__5051\ : Odrv4
    port map (
            O => \N__31368\,
            I => n2018
        );

    \I__5050\ : InMux
    port map (
            O => \N__31365\,
            I => \N__31362\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__31362\,
            I => n2085
        );

    \I__5048\ : CascadeMux
    port map (
            O => \N__31359\,
            I => \n2018_cascade_\
        );

    \I__5047\ : InMux
    port map (
            O => \N__31356\,
            I => \N__31352\
        );

    \I__5046\ : InMux
    port map (
            O => \N__31355\,
            I => \N__31349\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__31352\,
            I => \N__31346\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__31349\,
            I => \N__31342\
        );

    \I__5043\ : Span4Mux_v
    port map (
            O => \N__31346\,
            I => \N__31339\
        );

    \I__5042\ : InMux
    port map (
            O => \N__31345\,
            I => \N__31336\
        );

    \I__5041\ : Span4Mux_h
    port map (
            O => \N__31342\,
            I => \N__31333\
        );

    \I__5040\ : Span4Mux_h
    port map (
            O => \N__31339\,
            I => \N__31330\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__31336\,
            I => n2117
        );

    \I__5038\ : Odrv4
    port map (
            O => \N__31333\,
            I => n2117
        );

    \I__5037\ : Odrv4
    port map (
            O => \N__31330\,
            I => n2117
        );

    \I__5036\ : InMux
    port map (
            O => \N__31323\,
            I => \N__31320\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__31320\,
            I => \N__31317\
        );

    \I__5034\ : Odrv4
    port map (
            O => \N__31317\,
            I => n2089
        );

    \I__5033\ : InMux
    port map (
            O => \N__31314\,
            I => \N__31309\
        );

    \I__5032\ : InMux
    port map (
            O => \N__31313\,
            I => \N__31306\
        );

    \I__5031\ : CascadeMux
    port map (
            O => \N__31312\,
            I => \N__31303\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__31309\,
            I => \N__31300\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__31306\,
            I => \N__31297\
        );

    \I__5028\ : InMux
    port map (
            O => \N__31303\,
            I => \N__31294\
        );

    \I__5027\ : Span4Mux_h
    port map (
            O => \N__31300\,
            I => \N__31291\
        );

    \I__5026\ : Span4Mux_h
    port map (
            O => \N__31297\,
            I => \N__31288\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__31294\,
            I => \N__31285\
        );

    \I__5024\ : Odrv4
    port map (
            O => \N__31291\,
            I => n2121
        );

    \I__5023\ : Odrv4
    port map (
            O => \N__31288\,
            I => n2121
        );

    \I__5022\ : Odrv4
    port map (
            O => \N__31285\,
            I => n2121
        );

    \I__5021\ : InMux
    port map (
            O => \N__31278\,
            I => \N__31275\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__31275\,
            I => \N__31272\
        );

    \I__5019\ : Span4Mux_v
    port map (
            O => \N__31272\,
            I => \N__31269\
        );

    \I__5018\ : Odrv4
    port map (
            O => \N__31269\,
            I => n2501
        );

    \I__5017\ : InMux
    port map (
            O => \N__31266\,
            I => \bfn_6_21_0_\
        );

    \I__5016\ : InMux
    port map (
            O => \N__31263\,
            I => n12717
        );

    \I__5015\ : InMux
    port map (
            O => \N__31260\,
            I => n12651
        );

    \I__5014\ : InMux
    port map (
            O => \N__31257\,
            I => n12652
        );

    \I__5013\ : InMux
    port map (
            O => \N__31254\,
            I => \N__31251\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__31251\,
            I => \N__31248\
        );

    \I__5011\ : Odrv4
    port map (
            O => \N__31248\,
            I => n2086
        );

    \I__5010\ : InMux
    port map (
            O => \N__31245\,
            I => n12653
        );

    \I__5009\ : InMux
    port map (
            O => \N__31242\,
            I => \bfn_6_19_0_\
        );

    \I__5008\ : CascadeMux
    port map (
            O => \N__31239\,
            I => \N__31236\
        );

    \I__5007\ : InMux
    port map (
            O => \N__31236\,
            I => \N__31233\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__31233\,
            I => n2084
        );

    \I__5005\ : InMux
    port map (
            O => \N__31230\,
            I => n12655
        );

    \I__5004\ : InMux
    port map (
            O => \N__31227\,
            I => n12656
        );

    \I__5003\ : CascadeMux
    port map (
            O => \N__31224\,
            I => \N__31221\
        );

    \I__5002\ : InMux
    port map (
            O => \N__31221\,
            I => \N__31218\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__31218\,
            I => \N__31214\
        );

    \I__5000\ : InMux
    port map (
            O => \N__31217\,
            I => \N__31211\
        );

    \I__4999\ : Odrv4
    port map (
            O => \N__31214\,
            I => n2115
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__31211\,
            I => n2115
        );

    \I__4997\ : InMux
    port map (
            O => \N__31206\,
            I => \N__31203\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__31203\,
            I => n2091
        );

    \I__4995\ : CascadeMux
    port map (
            O => \N__31200\,
            I => \N__31196\
        );

    \I__4994\ : CascadeMux
    port map (
            O => \N__31199\,
            I => \N__31193\
        );

    \I__4993\ : InMux
    port map (
            O => \N__31196\,
            I => \N__31190\
        );

    \I__4992\ : InMux
    port map (
            O => \N__31193\,
            I => \N__31187\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__31190\,
            I => \N__31182\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__31187\,
            I => \N__31182\
        );

    \I__4989\ : Span4Mux_h
    port map (
            O => \N__31182\,
            I => \N__31178\
        );

    \I__4988\ : InMux
    port map (
            O => \N__31181\,
            I => \N__31175\
        );

    \I__4987\ : Odrv4
    port map (
            O => \N__31178\,
            I => n2123
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__31175\,
            I => n2123
        );

    \I__4985\ : CascadeMux
    port map (
            O => \N__31170\,
            I => \N__31167\
        );

    \I__4984\ : InMux
    port map (
            O => \N__31167\,
            I => \N__31164\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__31164\,
            I => \N__31161\
        );

    \I__4982\ : Span4Mux_h
    port map (
            O => \N__31161\,
            I => \N__31158\
        );

    \I__4981\ : Odrv4
    port map (
            O => \N__31158\,
            I => n2097
        );

    \I__4980\ : InMux
    port map (
            O => \N__31155\,
            I => n12642
        );

    \I__4979\ : InMux
    port map (
            O => \N__31152\,
            I => \N__31149\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__31149\,
            I => n2096
        );

    \I__4977\ : InMux
    port map (
            O => \N__31146\,
            I => n12643
        );

    \I__4976\ : InMux
    port map (
            O => \N__31143\,
            I => \N__31140\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__31140\,
            I => n2095
        );

    \I__4974\ : InMux
    port map (
            O => \N__31137\,
            I => n12644
        );

    \I__4973\ : CascadeMux
    port map (
            O => \N__31134\,
            I => \N__31131\
        );

    \I__4972\ : InMux
    port map (
            O => \N__31131\,
            I => \N__31128\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__31128\,
            I => n2094
        );

    \I__4970\ : InMux
    port map (
            O => \N__31125\,
            I => n12645
        );

    \I__4969\ : InMux
    port map (
            O => \N__31122\,
            I => \N__31119\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__31119\,
            I => n2093
        );

    \I__4967\ : InMux
    port map (
            O => \N__31116\,
            I => \bfn_6_18_0_\
        );

    \I__4966\ : InMux
    port map (
            O => \N__31113\,
            I => \N__31110\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__31110\,
            I => n2092
        );

    \I__4964\ : InMux
    port map (
            O => \N__31107\,
            I => n12647
        );

    \I__4963\ : InMux
    port map (
            O => \N__31104\,
            I => n12648
        );

    \I__4962\ : InMux
    port map (
            O => \N__31101\,
            I => \N__31098\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__31098\,
            I => n2090
        );

    \I__4960\ : InMux
    port map (
            O => \N__31095\,
            I => n12649
        );

    \I__4959\ : InMux
    port map (
            O => \N__31092\,
            I => n12650
        );

    \I__4958\ : InMux
    port map (
            O => \N__31089\,
            I => \N__31086\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__31086\,
            I => n14272
        );

    \I__4956\ : InMux
    port map (
            O => \N__31083\,
            I => \N__31080\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__31080\,
            I => n14268
        );

    \I__4954\ : CascadeMux
    port map (
            O => \N__31077\,
            I => \n14262_cascade_\
        );

    \I__4953\ : InMux
    port map (
            O => \N__31074\,
            I => \N__31071\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__31071\,
            I => n14282
        );

    \I__4951\ : InMux
    port map (
            O => \N__31068\,
            I => \N__31065\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__31065\,
            I => \N__31060\
        );

    \I__4949\ : InMux
    port map (
            O => \N__31064\,
            I => \N__31057\
        );

    \I__4948\ : InMux
    port map (
            O => \N__31063\,
            I => \N__31054\
        );

    \I__4947\ : Odrv4
    port map (
            O => \N__31060\,
            I => n3111
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__31057\,
            I => n3111
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__31054\,
            I => n3111
        );

    \I__4944\ : CascadeMux
    port map (
            O => \N__31047\,
            I => \N__31044\
        );

    \I__4943\ : InMux
    port map (
            O => \N__31044\,
            I => \N__31041\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__31041\,
            I => \N__31038\
        );

    \I__4941\ : Span4Mux_s1_v
    port map (
            O => \N__31038\,
            I => \N__31035\
        );

    \I__4940\ : Odrv4
    port map (
            O => \N__31035\,
            I => n3178
        );

    \I__4939\ : InMux
    port map (
            O => \N__31032\,
            I => \N__31029\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__31029\,
            I => \N__31024\
        );

    \I__4937\ : InMux
    port map (
            O => \N__31028\,
            I => \N__31021\
        );

    \I__4936\ : InMux
    port map (
            O => \N__31027\,
            I => \N__31018\
        );

    \I__4935\ : Odrv4
    port map (
            O => \N__31024\,
            I => n3110
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__31021\,
            I => n3110
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__31018\,
            I => n3110
        );

    \I__4932\ : InMux
    port map (
            O => \N__31011\,
            I => \N__31008\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__31008\,
            I => \N__31005\
        );

    \I__4930\ : Odrv4
    port map (
            O => \N__31005\,
            I => n3177
        );

    \I__4929\ : InMux
    port map (
            O => \N__31002\,
            I => \N__30999\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__30999\,
            I => \N__30996\
        );

    \I__4927\ : Odrv4
    port map (
            O => \N__30996\,
            I => n2283
        );

    \I__4926\ : CascadeMux
    port map (
            O => \N__30993\,
            I => \N__30989\
        );

    \I__4925\ : InMux
    port map (
            O => \N__30992\,
            I => \N__30986\
        );

    \I__4924\ : InMux
    port map (
            O => \N__30989\,
            I => \N__30982\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__30986\,
            I => \N__30979\
        );

    \I__4922\ : InMux
    port map (
            O => \N__30985\,
            I => \N__30976\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__30982\,
            I => \N__30973\
        );

    \I__4920\ : Span4Mux_v
    port map (
            O => \N__30979\,
            I => \N__30968\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__30976\,
            I => \N__30968\
        );

    \I__4918\ : Odrv4
    port map (
            O => \N__30973\,
            I => n2216
        );

    \I__4917\ : Odrv4
    port map (
            O => \N__30968\,
            I => n2216
        );

    \I__4916\ : InMux
    port map (
            O => \N__30963\,
            I => \N__30959\
        );

    \I__4915\ : InMux
    port map (
            O => \N__30962\,
            I => \N__30956\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__30959\,
            I => \N__30953\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__30956\,
            I => \N__30949\
        );

    \I__4912\ : Span4Mux_v
    port map (
            O => \N__30953\,
            I => \N__30946\
        );

    \I__4911\ : InMux
    port map (
            O => \N__30952\,
            I => \N__30943\
        );

    \I__4910\ : Span4Mux_v
    port map (
            O => \N__30949\,
            I => \N__30936\
        );

    \I__4909\ : Span4Mux_h
    port map (
            O => \N__30946\,
            I => \N__30936\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__30943\,
            I => \N__30936\
        );

    \I__4907\ : Span4Mux_v
    port map (
            O => \N__30936\,
            I => \N__30933\
        );

    \I__4906\ : Odrv4
    port map (
            O => \N__30933\,
            I => n2315
        );

    \I__4905\ : InMux
    port map (
            O => \N__30930\,
            I => \bfn_6_17_0_\
        );

    \I__4904\ : InMux
    port map (
            O => \N__30927\,
            I => n12639
        );

    \I__4903\ : CascadeMux
    port map (
            O => \N__30924\,
            I => \N__30921\
        );

    \I__4902\ : InMux
    port map (
            O => \N__30921\,
            I => \N__30918\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__30918\,
            I => n2099
        );

    \I__4900\ : InMux
    port map (
            O => \N__30915\,
            I => n12640
        );

    \I__4899\ : InMux
    port map (
            O => \N__30912\,
            I => \N__30909\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__30909\,
            I => n2098
        );

    \I__4897\ : InMux
    port map (
            O => \N__30906\,
            I => n12641
        );

    \I__4896\ : InMux
    port map (
            O => \N__30903\,
            I => \N__30900\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__30900\,
            I => \N__30897\
        );

    \I__4894\ : Odrv12
    port map (
            O => \N__30897\,
            I => n3185
        );

    \I__4893\ : InMux
    port map (
            O => \N__30894\,
            I => \N__30891\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__30891\,
            I => \N__30887\
        );

    \I__4891\ : InMux
    port map (
            O => \N__30890\,
            I => \N__30884\
        );

    \I__4890\ : Span4Mux_h
    port map (
            O => \N__30887\,
            I => \N__30878\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__30884\,
            I => \N__30878\
        );

    \I__4888\ : InMux
    port map (
            O => \N__30883\,
            I => \N__30875\
        );

    \I__4887\ : Odrv4
    port map (
            O => \N__30878\,
            I => n3118
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__30875\,
            I => n3118
        );

    \I__4885\ : CascadeMux
    port map (
            O => \N__30870\,
            I => \n27_adj_716_cascade_\
        );

    \I__4884\ : InMux
    port map (
            O => \N__30867\,
            I => \N__30864\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__30864\,
            I => n14266
        );

    \I__4882\ : InMux
    port map (
            O => \N__30861\,
            I => \N__30858\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__30858\,
            I => n35_adj_719
        );

    \I__4880\ : CascadeMux
    port map (
            O => \N__30855\,
            I => \n17_adj_714_cascade_\
        );

    \I__4879\ : InMux
    port map (
            O => \N__30852\,
            I => \N__30848\
        );

    \I__4878\ : InMux
    port map (
            O => \N__30851\,
            I => \N__30844\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__30848\,
            I => \N__30841\
        );

    \I__4876\ : InMux
    port map (
            O => \N__30847\,
            I => \N__30838\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__30844\,
            I => n3109
        );

    \I__4874\ : Odrv4
    port map (
            O => \N__30841\,
            I => n3109
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__30838\,
            I => n3109
        );

    \I__4872\ : CascadeMux
    port map (
            O => \N__30831\,
            I => \N__30828\
        );

    \I__4871\ : InMux
    port map (
            O => \N__30828\,
            I => \N__30825\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__30825\,
            I => \N__30822\
        );

    \I__4869\ : Odrv4
    port map (
            O => \N__30822\,
            I => n3176
        );

    \I__4868\ : CascadeMux
    port map (
            O => \N__30819\,
            I => \n33_adj_718_cascade_\
        );

    \I__4867\ : InMux
    port map (
            O => \N__30816\,
            I => \N__30813\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__30813\,
            I => \N__30808\
        );

    \I__4865\ : CascadeMux
    port map (
            O => \N__30812\,
            I => \N__30805\
        );

    \I__4864\ : CascadeMux
    port map (
            O => \N__30811\,
            I => \N__30802\
        );

    \I__4863\ : Span4Mux_h
    port map (
            O => \N__30808\,
            I => \N__30799\
        );

    \I__4862\ : InMux
    port map (
            O => \N__30805\,
            I => \N__30796\
        );

    \I__4861\ : InMux
    port map (
            O => \N__30802\,
            I => \N__30793\
        );

    \I__4860\ : Odrv4
    port map (
            O => \N__30799\,
            I => n3124
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__30796\,
            I => n3124
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__30793\,
            I => n3124
        );

    \I__4857\ : CascadeMux
    port map (
            O => \N__30786\,
            I => \N__30783\
        );

    \I__4856\ : InMux
    port map (
            O => \N__30783\,
            I => \N__30780\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__30780\,
            I => \N__30777\
        );

    \I__4854\ : Odrv4
    port map (
            O => \N__30777\,
            I => n3191
        );

    \I__4853\ : InMux
    port map (
            O => \N__30774\,
            I => \N__30771\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__30771\,
            I => n14804
        );

    \I__4851\ : CascadeMux
    port map (
            O => \N__30768\,
            I => \N__30765\
        );

    \I__4850\ : InMux
    port map (
            O => \N__30765\,
            I => \N__30762\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__30762\,
            I => n14025
        );

    \I__4848\ : CascadeMux
    port map (
            O => \N__30759\,
            I => \n3237_cascade_\
        );

    \I__4847\ : InMux
    port map (
            O => \N__30756\,
            I => \N__30753\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__30753\,
            I => n13_adj_713
        );

    \I__4845\ : InMux
    port map (
            O => \N__30750\,
            I => \N__30747\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__30747\,
            I => \N__30744\
        );

    \I__4843\ : Span4Mux_h
    port map (
            O => \N__30744\,
            I => \N__30741\
        );

    \I__4842\ : Odrv4
    port map (
            O => \N__30741\,
            I => n3179
        );

    \I__4841\ : InMux
    port map (
            O => \N__30738\,
            I => \N__30734\
        );

    \I__4840\ : InMux
    port map (
            O => \N__30737\,
            I => \N__30731\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__30734\,
            I => \N__30727\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__30731\,
            I => \N__30724\
        );

    \I__4837\ : InMux
    port map (
            O => \N__30730\,
            I => \N__30721\
        );

    \I__4836\ : Span4Mux_s3_h
    port map (
            O => \N__30727\,
            I => \N__30716\
        );

    \I__4835\ : Span4Mux_s1_v
    port map (
            O => \N__30724\,
            I => \N__30716\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__30721\,
            I => n3112
        );

    \I__4833\ : Odrv4
    port map (
            O => \N__30716\,
            I => n3112
        );

    \I__4832\ : InMux
    port map (
            O => \N__30711\,
            I => \N__30708\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__30708\,
            I => n14770
        );

    \I__4830\ : CascadeMux
    port map (
            O => \N__30705\,
            I => \n14776_cascade_\
        );

    \I__4829\ : InMux
    port map (
            O => \N__30702\,
            I => \N__30699\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__30699\,
            I => \N__30696\
        );

    \I__4827\ : Span4Mux_s3_v
    port map (
            O => \N__30696\,
            I => \N__30693\
        );

    \I__4826\ : Span4Mux_h
    port map (
            O => \N__30693\,
            I => \N__30689\
        );

    \I__4825\ : InMux
    port map (
            O => \N__30692\,
            I => \N__30686\
        );

    \I__4824\ : Odrv4
    port map (
            O => \N__30689\,
            I => n3122
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__30686\,
            I => n3122
        );

    \I__4822\ : CascadeMux
    port map (
            O => \N__30681\,
            I => \N__30678\
        );

    \I__4821\ : InMux
    port map (
            O => \N__30678\,
            I => \N__30675\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__30675\,
            I => \N__30672\
        );

    \I__4819\ : Odrv4
    port map (
            O => \N__30672\,
            I => n3189
        );

    \I__4818\ : InMux
    port map (
            O => \N__30669\,
            I => \N__30666\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__30666\,
            I => \N__30662\
        );

    \I__4816\ : InMux
    port map (
            O => \N__30665\,
            I => \N__30659\
        );

    \I__4815\ : Span4Mux_h
    port map (
            O => \N__30662\,
            I => \N__30653\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__30659\,
            I => \N__30653\
        );

    \I__4813\ : InMux
    port map (
            O => \N__30658\,
            I => \N__30650\
        );

    \I__4812\ : Odrv4
    port map (
            O => \N__30653\,
            I => n3116
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__30650\,
            I => n3116
        );

    \I__4810\ : CascadeMux
    port map (
            O => \N__30645\,
            I => \N__30642\
        );

    \I__4809\ : InMux
    port map (
            O => \N__30642\,
            I => \N__30639\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__30639\,
            I => \N__30636\
        );

    \I__4807\ : Odrv4
    port map (
            O => \N__30636\,
            I => n3183
        );

    \I__4806\ : CascadeMux
    port map (
            O => \N__30633\,
            I => \n3030_cascade_\
        );

    \I__4805\ : InMux
    port map (
            O => \N__30630\,
            I => \N__30627\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__30627\,
            I => n11947
        );

    \I__4803\ : CascadeMux
    port map (
            O => \N__30624\,
            I => \N__30620\
        );

    \I__4802\ : InMux
    port map (
            O => \N__30623\,
            I => \N__30617\
        );

    \I__4801\ : InMux
    port map (
            O => \N__30620\,
            I => \N__30614\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__30617\,
            I => \N__30609\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__30614\,
            I => \N__30609\
        );

    \I__4798\ : Span4Mux_h
    port map (
            O => \N__30609\,
            I => \N__30605\
        );

    \I__4797\ : InMux
    port map (
            O => \N__30608\,
            I => \N__30602\
        );

    \I__4796\ : Odrv4
    port map (
            O => \N__30605\,
            I => n3019
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__30602\,
            I => n3019
        );

    \I__4794\ : CascadeMux
    port map (
            O => \N__30597\,
            I => \N__30594\
        );

    \I__4793\ : InMux
    port map (
            O => \N__30594\,
            I => \N__30591\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__30591\,
            I => \N__30588\
        );

    \I__4791\ : Span4Mux_v
    port map (
            O => \N__30588\,
            I => \N__30584\
        );

    \I__4790\ : CascadeMux
    port map (
            O => \N__30587\,
            I => \N__30581\
        );

    \I__4789\ : Span4Mux_s0_h
    port map (
            O => \N__30584\,
            I => \N__30577\
        );

    \I__4788\ : InMux
    port map (
            O => \N__30581\,
            I => \N__30574\
        );

    \I__4787\ : InMux
    port map (
            O => \N__30580\,
            I => \N__30571\
        );

    \I__4786\ : Odrv4
    port map (
            O => \N__30577\,
            I => n3027
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__30574\,
            I => n3027
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__30571\,
            I => n3027
        );

    \I__4783\ : CascadeMux
    port map (
            O => \N__30564\,
            I => \n13871_cascade_\
        );

    \I__4782\ : CascadeMux
    port map (
            O => \N__30561\,
            I => \N__30557\
        );

    \I__4781\ : InMux
    port map (
            O => \N__30560\,
            I => \N__30554\
        );

    \I__4780\ : InMux
    port map (
            O => \N__30557\,
            I => \N__30551\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__30554\,
            I => \N__30548\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__30551\,
            I => \N__30545\
        );

    \I__4777\ : Span4Mux_v
    port map (
            O => \N__30548\,
            I => \N__30541\
        );

    \I__4776\ : Span4Mux_v
    port map (
            O => \N__30545\,
            I => \N__30538\
        );

    \I__4775\ : InMux
    port map (
            O => \N__30544\,
            I => \N__30535\
        );

    \I__4774\ : Odrv4
    port map (
            O => \N__30541\,
            I => n3023
        );

    \I__4773\ : Odrv4
    port map (
            O => \N__30538\,
            I => n3023
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__30535\,
            I => n3023
        );

    \I__4771\ : CascadeMux
    port map (
            O => \N__30528\,
            I => \N__30525\
        );

    \I__4770\ : InMux
    port map (
            O => \N__30525\,
            I => \N__30522\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__30522\,
            I => n14078
        );

    \I__4768\ : InMux
    port map (
            O => \N__30519\,
            I => \N__30516\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__30516\,
            I => \N__30513\
        );

    \I__4766\ : Odrv4
    port map (
            O => \N__30513\,
            I => n3199
        );

    \I__4765\ : CascadeMux
    port map (
            O => \N__30510\,
            I => \N__30507\
        );

    \I__4764\ : InMux
    port map (
            O => \N__30507\,
            I => \N__30503\
        );

    \I__4763\ : InMux
    port map (
            O => \N__30506\,
            I => \N__30500\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__30503\,
            I => \N__30497\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__30500\,
            I => n3132
        );

    \I__4760\ : Odrv4
    port map (
            O => \N__30497\,
            I => n3132
        );

    \I__4759\ : CascadeMux
    port map (
            O => \N__30492\,
            I => \N__30489\
        );

    \I__4758\ : InMux
    port map (
            O => \N__30489\,
            I => \N__30485\
        );

    \I__4757\ : InMux
    port map (
            O => \N__30488\,
            I => \N__30481\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__30485\,
            I => \N__30478\
        );

    \I__4755\ : InMux
    port map (
            O => \N__30484\,
            I => \N__30475\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__30481\,
            I => n3129
        );

    \I__4753\ : Odrv4
    port map (
            O => \N__30478\,
            I => n3129
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__30475\,
            I => n3129
        );

    \I__4751\ : CascadeMux
    port map (
            O => \N__30468\,
            I => \N__30465\
        );

    \I__4750\ : InMux
    port map (
            O => \N__30465\,
            I => \N__30462\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__30462\,
            I => \N__30459\
        );

    \I__4748\ : Span4Mux_h
    port map (
            O => \N__30459\,
            I => \N__30456\
        );

    \I__4747\ : Odrv4
    port map (
            O => \N__30456\,
            I => n3196
        );

    \I__4746\ : CascadeMux
    port map (
            O => \N__30453\,
            I => \n3228_cascade_\
        );

    \I__4745\ : InMux
    port map (
            O => \N__30450\,
            I => \N__30447\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__30447\,
            I => n14768
        );

    \I__4743\ : InMux
    port map (
            O => \N__30444\,
            I => \N__30441\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__30441\,
            I => \N__30438\
        );

    \I__4741\ : Span4Mux_h
    port map (
            O => \N__30438\,
            I => \N__30435\
        );

    \I__4740\ : Odrv4
    port map (
            O => \N__30435\,
            I => n3200
        );

    \I__4739\ : CascadeMux
    port map (
            O => \N__30432\,
            I => \N__30428\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__30431\,
            I => \N__30425\
        );

    \I__4737\ : InMux
    port map (
            O => \N__30428\,
            I => \N__30422\
        );

    \I__4736\ : InMux
    port map (
            O => \N__30425\,
            I => \N__30418\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__30422\,
            I => \N__30415\
        );

    \I__4734\ : InMux
    port map (
            O => \N__30421\,
            I => \N__30412\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__30418\,
            I => n3133
        );

    \I__4732\ : Odrv4
    port map (
            O => \N__30415\,
            I => n3133
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__30412\,
            I => n3133
        );

    \I__4730\ : InMux
    port map (
            O => \N__30405\,
            I => \N__30402\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__30402\,
            I => \N__30399\
        );

    \I__4728\ : Odrv4
    port map (
            O => \N__30399\,
            I => n3198
        );

    \I__4727\ : CascadeMux
    port map (
            O => \N__30396\,
            I => \N__30393\
        );

    \I__4726\ : InMux
    port map (
            O => \N__30393\,
            I => \N__30390\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__30390\,
            I => \N__30386\
        );

    \I__4724\ : InMux
    port map (
            O => \N__30389\,
            I => \N__30382\
        );

    \I__4723\ : Span4Mux_v
    port map (
            O => \N__30386\,
            I => \N__30379\
        );

    \I__4722\ : InMux
    port map (
            O => \N__30385\,
            I => \N__30376\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__30382\,
            I => n3131
        );

    \I__4720\ : Odrv4
    port map (
            O => \N__30379\,
            I => n3131
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__30376\,
            I => n3131
        );

    \I__4718\ : InMux
    port map (
            O => \N__30369\,
            I => \N__30365\
        );

    \I__4717\ : InMux
    port map (
            O => \N__30368\,
            I => \N__30362\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__30365\,
            I => \N__30359\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__30362\,
            I => \N__30356\
        );

    \I__4714\ : Span4Mux_v
    port map (
            O => \N__30359\,
            I => \N__30352\
        );

    \I__4713\ : Span4Mux_s3_h
    port map (
            O => \N__30356\,
            I => \N__30349\
        );

    \I__4712\ : InMux
    port map (
            O => \N__30355\,
            I => \N__30346\
        );

    \I__4711\ : Odrv4
    port map (
            O => \N__30352\,
            I => n2917
        );

    \I__4710\ : Odrv4
    port map (
            O => \N__30349\,
            I => n2917
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__30346\,
            I => n2917
        );

    \I__4708\ : CascadeMux
    port map (
            O => \N__30339\,
            I => \N__30336\
        );

    \I__4707\ : InMux
    port map (
            O => \N__30336\,
            I => \N__30333\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__30333\,
            I => \N__30330\
        );

    \I__4705\ : Span4Mux_v
    port map (
            O => \N__30330\,
            I => \N__30327\
        );

    \I__4704\ : Odrv4
    port map (
            O => \N__30327\,
            I => n2984
        );

    \I__4703\ : InMux
    port map (
            O => \N__30324\,
            I => \N__30320\
        );

    \I__4702\ : InMux
    port map (
            O => \N__30323\,
            I => \N__30317\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__30320\,
            I => \N__30314\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__30317\,
            I => \N__30311\
        );

    \I__4699\ : Span4Mux_s1_v
    port map (
            O => \N__30314\,
            I => \N__30307\
        );

    \I__4698\ : Span4Mux_s3_v
    port map (
            O => \N__30311\,
            I => \N__30304\
        );

    \I__4697\ : InMux
    port map (
            O => \N__30310\,
            I => \N__30301\
        );

    \I__4696\ : Odrv4
    port map (
            O => \N__30307\,
            I => n3016
        );

    \I__4695\ : Odrv4
    port map (
            O => \N__30304\,
            I => n3016
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__30301\,
            I => n3016
        );

    \I__4693\ : InMux
    port map (
            O => \N__30294\,
            I => \N__30291\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__30291\,
            I => \N__30287\
        );

    \I__4691\ : InMux
    port map (
            O => \N__30290\,
            I => \N__30283\
        );

    \I__4690\ : Span4Mux_h
    port map (
            O => \N__30287\,
            I => \N__30280\
        );

    \I__4689\ : InMux
    port map (
            O => \N__30286\,
            I => \N__30277\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__30283\,
            I => n2913
        );

    \I__4687\ : Odrv4
    port map (
            O => \N__30280\,
            I => n2913
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__30277\,
            I => n2913
        );

    \I__4685\ : CascadeMux
    port map (
            O => \N__30270\,
            I => \N__30267\
        );

    \I__4684\ : InMux
    port map (
            O => \N__30267\,
            I => \N__30264\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__30264\,
            I => \N__30261\
        );

    \I__4682\ : Odrv4
    port map (
            O => \N__30261\,
            I => n2980
        );

    \I__4681\ : CascadeMux
    port map (
            O => \N__30258\,
            I => \N__30255\
        );

    \I__4680\ : InMux
    port map (
            O => \N__30255\,
            I => \N__30252\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__30252\,
            I => \N__30248\
        );

    \I__4678\ : InMux
    port map (
            O => \N__30251\,
            I => \N__30245\
        );

    \I__4677\ : Span4Mux_s1_v
    port map (
            O => \N__30248\,
            I => \N__30242\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__30245\,
            I => \N__30239\
        );

    \I__4675\ : Span4Mux_v
    port map (
            O => \N__30242\,
            I => \N__30235\
        );

    \I__4674\ : Span4Mux_h
    port map (
            O => \N__30239\,
            I => \N__30232\
        );

    \I__4673\ : InMux
    port map (
            O => \N__30238\,
            I => \N__30229\
        );

    \I__4672\ : Odrv4
    port map (
            O => \N__30235\,
            I => n3012
        );

    \I__4671\ : Odrv4
    port map (
            O => \N__30232\,
            I => n3012
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__30229\,
            I => n3012
        );

    \I__4669\ : InMux
    port map (
            O => \N__30222\,
            I => \N__30217\
        );

    \I__4668\ : InMux
    port map (
            O => \N__30221\,
            I => \N__30214\
        );

    \I__4667\ : InMux
    port map (
            O => \N__30220\,
            I => \N__30211\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__30217\,
            I => \N__30208\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__30214\,
            I => \N__30203\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__30211\,
            I => \N__30203\
        );

    \I__4663\ : Odrv4
    port map (
            O => \N__30208\,
            I => n2933
        );

    \I__4662\ : Odrv4
    port map (
            O => \N__30203\,
            I => n2933
        );

    \I__4661\ : InMux
    port map (
            O => \N__30198\,
            I => \N__30195\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__30195\,
            I => n12053
        );

    \I__4659\ : InMux
    port map (
            O => \N__30192\,
            I => \N__30189\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__30189\,
            I => \N__30186\
        );

    \I__4657\ : Span4Mux_h
    port map (
            O => \N__30186\,
            I => \N__30183\
        );

    \I__4656\ : Odrv4
    port map (
            O => \N__30183\,
            I => n2987
        );

    \I__4655\ : CascadeMux
    port map (
            O => \N__30180\,
            I => \N__30176\
        );

    \I__4654\ : InMux
    port map (
            O => \N__30179\,
            I => \N__30173\
        );

    \I__4653\ : InMux
    port map (
            O => \N__30176\,
            I => \N__30169\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__30173\,
            I => \N__30166\
        );

    \I__4651\ : InMux
    port map (
            O => \N__30172\,
            I => \N__30163\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__30169\,
            I => n2920
        );

    \I__4649\ : Odrv4
    port map (
            O => \N__30166\,
            I => n2920
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__30163\,
            I => n2920
        );

    \I__4647\ : InMux
    port map (
            O => \N__30156\,
            I => \N__30153\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__30153\,
            I => \N__30150\
        );

    \I__4645\ : Span4Mux_h
    port map (
            O => \N__30150\,
            I => \N__30147\
        );

    \I__4644\ : Odrv4
    port map (
            O => \N__30147\,
            I => n2999
        );

    \I__4643\ : CascadeMux
    port map (
            O => \N__30144\,
            I => \N__30141\
        );

    \I__4642\ : InMux
    port map (
            O => \N__30141\,
            I => \N__30137\
        );

    \I__4641\ : InMux
    port map (
            O => \N__30140\,
            I => \N__30134\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__30137\,
            I => \N__30131\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__30134\,
            I => \N__30127\
        );

    \I__4638\ : Span4Mux_h
    port map (
            O => \N__30131\,
            I => \N__30124\
        );

    \I__4637\ : InMux
    port map (
            O => \N__30130\,
            I => \N__30121\
        );

    \I__4636\ : Span4Mux_h
    port map (
            O => \N__30127\,
            I => \N__30118\
        );

    \I__4635\ : Odrv4
    port map (
            O => \N__30124\,
            I => n2932
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__30121\,
            I => n2932
        );

    \I__4633\ : Odrv4
    port map (
            O => \N__30118\,
            I => n2932
        );

    \I__4632\ : InMux
    port map (
            O => \N__30111\,
            I => \N__30108\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__30108\,
            I => \N__30105\
        );

    \I__4630\ : Span4Mux_v
    port map (
            O => \N__30105\,
            I => \N__30102\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__30102\,
            I => n3001
        );

    \I__4628\ : CascadeMux
    port map (
            O => \N__30099\,
            I => \N__30096\
        );

    \I__4627\ : InMux
    port map (
            O => \N__30096\,
            I => \N__30092\
        );

    \I__4626\ : InMux
    port map (
            O => \N__30095\,
            I => \N__30089\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__30092\,
            I => \N__30086\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__30089\,
            I => n3033
        );

    \I__4623\ : Odrv4
    port map (
            O => \N__30086\,
            I => n3033
        );

    \I__4622\ : CascadeMux
    port map (
            O => \N__30081\,
            I => \n3033_cascade_\
        );

    \I__4621\ : CascadeMux
    port map (
            O => \N__30078\,
            I => \N__30074\
        );

    \I__4620\ : InMux
    port map (
            O => \N__30077\,
            I => \N__30070\
        );

    \I__4619\ : InMux
    port map (
            O => \N__30074\,
            I => \N__30067\
        );

    \I__4618\ : InMux
    port map (
            O => \N__30073\,
            I => \N__30064\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__30070\,
            I => n3032
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__30067\,
            I => n3032
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__30064\,
            I => n3032
        );

    \I__4614\ : InMux
    port map (
            O => \N__30057\,
            I => \N__30054\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__30054\,
            I => \N__30051\
        );

    \I__4612\ : Span4Mux_h
    port map (
            O => \N__30051\,
            I => \N__30048\
        );

    \I__4611\ : Odrv4
    port map (
            O => \N__30048\,
            I => n3182
        );

    \I__4610\ : CascadeMux
    port map (
            O => \N__30045\,
            I => \N__30042\
        );

    \I__4609\ : InMux
    port map (
            O => \N__30042\,
            I => \N__30039\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__30039\,
            I => \N__30035\
        );

    \I__4607\ : InMux
    port map (
            O => \N__30038\,
            I => \N__30032\
        );

    \I__4606\ : Span4Mux_h
    port map (
            O => \N__30035\,
            I => \N__30027\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__30032\,
            I => \N__30027\
        );

    \I__4604\ : Span4Mux_v
    port map (
            O => \N__30027\,
            I => \N__30024\
        );

    \I__4603\ : Odrv4
    port map (
            O => \N__30024\,
            I => n3115
        );

    \I__4602\ : InMux
    port map (
            O => \N__30021\,
            I => \N__30018\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__30018\,
            I => \N__30015\
        );

    \I__4600\ : Span4Mux_h
    port map (
            O => \N__30015\,
            I => \N__30012\
        );

    \I__4599\ : Odrv4
    port map (
            O => \N__30012\,
            I => n2998
        );

    \I__4598\ : CascadeMux
    port map (
            O => \N__30009\,
            I => \N__30004\
        );

    \I__4597\ : CascadeMux
    port map (
            O => \N__30008\,
            I => \N__30001\
        );

    \I__4596\ : InMux
    port map (
            O => \N__30007\,
            I => \N__29998\
        );

    \I__4595\ : InMux
    port map (
            O => \N__30004\,
            I => \N__29995\
        );

    \I__4594\ : InMux
    port map (
            O => \N__30001\,
            I => \N__29992\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__29998\,
            I => \N__29989\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__29995\,
            I => \N__29984\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__29992\,
            I => \N__29984\
        );

    \I__4590\ : Odrv4
    port map (
            O => \N__29989\,
            I => n2931
        );

    \I__4589\ : Odrv4
    port map (
            O => \N__29984\,
            I => n2931
        );

    \I__4588\ : CascadeMux
    port map (
            O => \N__29979\,
            I => \N__29975\
        );

    \I__4587\ : CascadeMux
    port map (
            O => \N__29978\,
            I => \N__29972\
        );

    \I__4586\ : InMux
    port map (
            O => \N__29975\,
            I => \N__29969\
        );

    \I__4585\ : InMux
    port map (
            O => \N__29972\,
            I => \N__29966\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__29969\,
            I => \N__29963\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__29966\,
            I => n3030
        );

    \I__4582\ : Odrv4
    port map (
            O => \N__29963\,
            I => n3030
        );

    \I__4581\ : InMux
    port map (
            O => \N__29958\,
            I => \N__29955\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__29955\,
            I => \N__29951\
        );

    \I__4579\ : CascadeMux
    port map (
            O => \N__29954\,
            I => \N__29948\
        );

    \I__4578\ : Span4Mux_v
    port map (
            O => \N__29951\,
            I => \N__29944\
        );

    \I__4577\ : InMux
    port map (
            O => \N__29948\,
            I => \N__29941\
        );

    \I__4576\ : InMux
    port map (
            O => \N__29947\,
            I => \N__29938\
        );

    \I__4575\ : Odrv4
    port map (
            O => \N__29944\,
            I => n3029
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__29941\,
            I => n3029
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__29938\,
            I => n3029
        );

    \I__4572\ : CascadeMux
    port map (
            O => \N__29931\,
            I => \N__29928\
        );

    \I__4571\ : InMux
    port map (
            O => \N__29928\,
            I => \N__29923\
        );

    \I__4570\ : InMux
    port map (
            O => \N__29927\,
            I => \N__29920\
        );

    \I__4569\ : InMux
    port map (
            O => \N__29926\,
            I => \N__29917\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__29923\,
            I => \N__29914\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__29920\,
            I => n3031
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__29917\,
            I => n3031
        );

    \I__4565\ : Odrv4
    port map (
            O => \N__29914\,
            I => n3031
        );

    \I__4564\ : InMux
    port map (
            O => \N__29907\,
            I => \N__29904\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__29904\,
            I => \N__29901\
        );

    \I__4562\ : Span4Mux_v
    port map (
            O => \N__29901\,
            I => \N__29898\
        );

    \I__4561\ : Odrv4
    port map (
            O => \N__29898\,
            I => n2896
        );

    \I__4560\ : CascadeMux
    port map (
            O => \N__29895\,
            I => \N__29892\
        );

    \I__4559\ : InMux
    port map (
            O => \N__29892\,
            I => \N__29889\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__29889\,
            I => \N__29885\
        );

    \I__4557\ : InMux
    port map (
            O => \N__29888\,
            I => \N__29881\
        );

    \I__4556\ : Span4Mux_v
    port map (
            O => \N__29885\,
            I => \N__29878\
        );

    \I__4555\ : CascadeMux
    port map (
            O => \N__29884\,
            I => \N__29875\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__29881\,
            I => \N__29872\
        );

    \I__4553\ : Span4Mux_h
    port map (
            O => \N__29878\,
            I => \N__29869\
        );

    \I__4552\ : InMux
    port map (
            O => \N__29875\,
            I => \N__29866\
        );

    \I__4551\ : Span4Mux_v
    port map (
            O => \N__29872\,
            I => \N__29863\
        );

    \I__4550\ : Odrv4
    port map (
            O => \N__29869\,
            I => n2829
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__29866\,
            I => n2829
        );

    \I__4548\ : Odrv4
    port map (
            O => \N__29863\,
            I => n2829
        );

    \I__4547\ : InMux
    port map (
            O => \N__29856\,
            I => \N__29853\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__29853\,
            I => \N__29849\
        );

    \I__4545\ : InMux
    port map (
            O => \N__29852\,
            I => \N__29845\
        );

    \I__4544\ : Span4Mux_h
    port map (
            O => \N__29849\,
            I => \N__29842\
        );

    \I__4543\ : InMux
    port map (
            O => \N__29848\,
            I => \N__29839\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__29845\,
            I => n2928
        );

    \I__4541\ : Odrv4
    port map (
            O => \N__29842\,
            I => n2928
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__29839\,
            I => n2928
        );

    \I__4539\ : InMux
    port map (
            O => \N__29832\,
            I => \N__29828\
        );

    \I__4538\ : CascadeMux
    port map (
            O => \N__29831\,
            I => \N__29824\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__29828\,
            I => \N__29821\
        );

    \I__4536\ : InMux
    port map (
            O => \N__29827\,
            I => \N__29818\
        );

    \I__4535\ : InMux
    port map (
            O => \N__29824\,
            I => \N__29815\
        );

    \I__4534\ : Span4Mux_h
    port map (
            O => \N__29821\,
            I => \N__29810\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__29818\,
            I => \N__29810\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__29815\,
            I => n2821
        );

    \I__4531\ : Odrv4
    port map (
            O => \N__29810\,
            I => n2821
        );

    \I__4530\ : InMux
    port map (
            O => \N__29805\,
            I => \N__29802\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__29802\,
            I => \N__29799\
        );

    \I__4528\ : Span4Mux_h
    port map (
            O => \N__29799\,
            I => \N__29796\
        );

    \I__4527\ : Odrv4
    port map (
            O => \N__29796\,
            I => n2888
        );

    \I__4526\ : InMux
    port map (
            O => \N__29793\,
            I => \N__29790\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__29790\,
            I => \N__29787\
        );

    \I__4524\ : Span4Mux_v
    port map (
            O => \N__29787\,
            I => \N__29784\
        );

    \I__4523\ : Odrv4
    port map (
            O => \N__29784\,
            I => n2881
        );

    \I__4522\ : CascadeMux
    port map (
            O => \N__29781\,
            I => \N__29778\
        );

    \I__4521\ : InMux
    port map (
            O => \N__29778\,
            I => \N__29775\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__29775\,
            I => \N__29771\
        );

    \I__4519\ : InMux
    port map (
            O => \N__29774\,
            I => \N__29768\
        );

    \I__4518\ : Span4Mux_v
    port map (
            O => \N__29771\,
            I => \N__29762\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__29768\,
            I => \N__29762\
        );

    \I__4516\ : InMux
    port map (
            O => \N__29767\,
            I => \N__29759\
        );

    \I__4515\ : Span4Mux_h
    port map (
            O => \N__29762\,
            I => \N__29756\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__29759\,
            I => n2814
        );

    \I__4513\ : Odrv4
    port map (
            O => \N__29756\,
            I => n2814
        );

    \I__4512\ : InMux
    port map (
            O => \N__29751\,
            I => \N__29748\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__29748\,
            I => \N__29745\
        );

    \I__4510\ : Span4Mux_v
    port map (
            O => \N__29745\,
            I => \N__29742\
        );

    \I__4509\ : Odrv4
    port map (
            O => \N__29742\,
            I => n2893
        );

    \I__4508\ : CascadeMux
    port map (
            O => \N__29739\,
            I => \N__29736\
        );

    \I__4507\ : InMux
    port map (
            O => \N__29736\,
            I => \N__29733\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__29733\,
            I => \N__29729\
        );

    \I__4505\ : CascadeMux
    port map (
            O => \N__29732\,
            I => \N__29726\
        );

    \I__4504\ : Span4Mux_v
    port map (
            O => \N__29729\,
            I => \N__29723\
        );

    \I__4503\ : InMux
    port map (
            O => \N__29726\,
            I => \N__29720\
        );

    \I__4502\ : Odrv4
    port map (
            O => \N__29723\,
            I => n2826
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__29720\,
            I => n2826
        );

    \I__4500\ : CascadeMux
    port map (
            O => \N__29715\,
            I => \N__29712\
        );

    \I__4499\ : InMux
    port map (
            O => \N__29712\,
            I => \N__29709\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__29709\,
            I => \N__29705\
        );

    \I__4497\ : InMux
    port map (
            O => \N__29708\,
            I => \N__29702\
        );

    \I__4496\ : Span4Mux_v
    port map (
            O => \N__29705\,
            I => \N__29696\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__29702\,
            I => \N__29696\
        );

    \I__4494\ : InMux
    port map (
            O => \N__29701\,
            I => \N__29693\
        );

    \I__4493\ : Odrv4
    port map (
            O => \N__29696\,
            I => n2925
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__29693\,
            I => n2925
        );

    \I__4491\ : CascadeMux
    port map (
            O => \N__29688\,
            I => \N__29685\
        );

    \I__4490\ : InMux
    port map (
            O => \N__29685\,
            I => \N__29680\
        );

    \I__4489\ : InMux
    port map (
            O => \N__29684\,
            I => \N__29677\
        );

    \I__4488\ : InMux
    port map (
            O => \N__29683\,
            I => \N__29674\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__29680\,
            I => \N__29671\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__29677\,
            I => \N__29668\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__29674\,
            I => \N__29665\
        );

    \I__4484\ : Span4Mux_h
    port map (
            O => \N__29671\,
            I => \N__29662\
        );

    \I__4483\ : Span12Mux_s4_h
    port map (
            O => \N__29668\,
            I => \N__29659\
        );

    \I__4482\ : Span4Mux_h
    port map (
            O => \N__29665\,
            I => \N__29656\
        );

    \I__4481\ : Odrv4
    port map (
            O => \N__29662\,
            I => n2615
        );

    \I__4480\ : Odrv12
    port map (
            O => \N__29659\,
            I => n2615
        );

    \I__4479\ : Odrv4
    port map (
            O => \N__29656\,
            I => n2615
        );

    \I__4478\ : CascadeMux
    port map (
            O => \N__29649\,
            I => \N__29645\
        );

    \I__4477\ : InMux
    port map (
            O => \N__29648\,
            I => \N__29642\
        );

    \I__4476\ : InMux
    port map (
            O => \N__29645\,
            I => \N__29639\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__29642\,
            I => \N__29636\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__29639\,
            I => \N__29632\
        );

    \I__4473\ : Span4Mux_v
    port map (
            O => \N__29636\,
            I => \N__29629\
        );

    \I__4472\ : InMux
    port map (
            O => \N__29635\,
            I => \N__29626\
        );

    \I__4471\ : Span4Mux_s2_h
    port map (
            O => \N__29632\,
            I => \N__29623\
        );

    \I__4470\ : Odrv4
    port map (
            O => \N__29629\,
            I => n2831
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__29626\,
            I => n2831
        );

    \I__4468\ : Odrv4
    port map (
            O => \N__29623\,
            I => n2831
        );

    \I__4467\ : CascadeMux
    port map (
            O => \N__29616\,
            I => \N__29613\
        );

    \I__4466\ : InMux
    port map (
            O => \N__29613\,
            I => \N__29610\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__29610\,
            I => \N__29607\
        );

    \I__4464\ : Span4Mux_v
    port map (
            O => \N__29607\,
            I => \N__29604\
        );

    \I__4463\ : Span4Mux_h
    port map (
            O => \N__29604\,
            I => \N__29601\
        );

    \I__4462\ : Odrv4
    port map (
            O => \N__29601\,
            I => n2898
        );

    \I__4461\ : CascadeMux
    port map (
            O => \N__29598\,
            I => \N__29595\
        );

    \I__4460\ : InMux
    port map (
            O => \N__29595\,
            I => \N__29592\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__29592\,
            I => \N__29587\
        );

    \I__4458\ : InMux
    port map (
            O => \N__29591\,
            I => \N__29582\
        );

    \I__4457\ : InMux
    port map (
            O => \N__29590\,
            I => \N__29582\
        );

    \I__4456\ : Span4Mux_v
    port map (
            O => \N__29587\,
            I => \N__29579\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__29582\,
            I => n2930
        );

    \I__4454\ : Odrv4
    port map (
            O => \N__29579\,
            I => n2930
        );

    \I__4453\ : InMux
    port map (
            O => \N__29574\,
            I => \N__29571\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__29571\,
            I => \N__29568\
        );

    \I__4451\ : Span4Mux_h
    port map (
            O => \N__29568\,
            I => \N__29565\
        );

    \I__4450\ : Odrv4
    port map (
            O => \N__29565\,
            I => n2991
        );

    \I__4449\ : InMux
    port map (
            O => \N__29562\,
            I => \N__29558\
        );

    \I__4448\ : InMux
    port map (
            O => \N__29561\,
            I => \N__29555\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__29558\,
            I => \N__29552\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__29555\,
            I => n2924
        );

    \I__4445\ : Odrv4
    port map (
            O => \N__29552\,
            I => n2924
        );

    \I__4444\ : CascadeMux
    port map (
            O => \N__29547\,
            I => \n2513_cascade_\
        );

    \I__4443\ : InMux
    port map (
            O => \N__29544\,
            I => \N__29541\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__29541\,
            I => \N__29537\
        );

    \I__4441\ : InMux
    port map (
            O => \N__29540\,
            I => \N__29534\
        );

    \I__4440\ : Span4Mux_h
    port map (
            O => \N__29537\,
            I => \N__29530\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__29534\,
            I => \N__29527\
        );

    \I__4438\ : InMux
    port map (
            O => \N__29533\,
            I => \N__29524\
        );

    \I__4437\ : Span4Mux_v
    port map (
            O => \N__29530\,
            I => \N__29521\
        );

    \I__4436\ : Span4Mux_v
    port map (
            O => \N__29527\,
            I => \N__29516\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__29524\,
            I => \N__29516\
        );

    \I__4434\ : Span4Mux_v
    port map (
            O => \N__29521\,
            I => \N__29511\
        );

    \I__4433\ : Span4Mux_h
    port map (
            O => \N__29516\,
            I => \N__29511\
        );

    \I__4432\ : Odrv4
    port map (
            O => \N__29511\,
            I => n2612
        );

    \I__4431\ : CascadeMux
    port map (
            O => \N__29508\,
            I => \N__29505\
        );

    \I__4430\ : InMux
    port map (
            O => \N__29505\,
            I => \N__29502\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__29502\,
            I => \N__29497\
        );

    \I__4428\ : InMux
    port map (
            O => \N__29501\,
            I => \N__29494\
        );

    \I__4427\ : InMux
    port map (
            O => \N__29500\,
            I => \N__29491\
        );

    \I__4426\ : Span4Mux_h
    port map (
            O => \N__29497\,
            I => \N__29488\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__29494\,
            I => \N__29483\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__29491\,
            I => \N__29483\
        );

    \I__4423\ : Span4Mux_v
    port map (
            O => \N__29488\,
            I => \N__29480\
        );

    \I__4422\ : Span4Mux_h
    port map (
            O => \N__29483\,
            I => \N__29475\
        );

    \I__4421\ : Span4Mux_v
    port map (
            O => \N__29480\,
            I => \N__29475\
        );

    \I__4420\ : Odrv4
    port map (
            O => \N__29475\,
            I => n2629
        );

    \I__4419\ : InMux
    port map (
            O => \N__29472\,
            I => \N__29469\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__29469\,
            I => \N__29466\
        );

    \I__4417\ : Span4Mux_v
    port map (
            O => \N__29466\,
            I => \N__29463\
        );

    \I__4416\ : Odrv4
    port map (
            O => \N__29463\,
            I => n2899
        );

    \I__4415\ : CascadeMux
    port map (
            O => \N__29460\,
            I => \N__29457\
        );

    \I__4414\ : InMux
    port map (
            O => \N__29457\,
            I => \N__29454\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__29454\,
            I => \N__29450\
        );

    \I__4412\ : InMux
    port map (
            O => \N__29453\,
            I => \N__29447\
        );

    \I__4411\ : Span4Mux_s3_h
    port map (
            O => \N__29450\,
            I => \N__29444\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__29447\,
            I => n2832
        );

    \I__4409\ : Odrv4
    port map (
            O => \N__29444\,
            I => n2832
        );

    \I__4408\ : CascadeMux
    port map (
            O => \N__29439\,
            I => \N__29435\
        );

    \I__4407\ : CascadeMux
    port map (
            O => \N__29438\,
            I => \N__29431\
        );

    \I__4406\ : InMux
    port map (
            O => \N__29435\,
            I => \N__29428\
        );

    \I__4405\ : InMux
    port map (
            O => \N__29434\,
            I => \N__29425\
        );

    \I__4404\ : InMux
    port map (
            O => \N__29431\,
            I => \N__29422\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__29428\,
            I => \N__29419\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__29425\,
            I => \N__29416\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__29422\,
            I => \N__29413\
        );

    \I__4400\ : Span12Mux_s3_h
    port map (
            O => \N__29419\,
            I => \N__29410\
        );

    \I__4399\ : Span4Mux_v
    port map (
            O => \N__29416\,
            I => \N__29407\
        );

    \I__4398\ : Span4Mux_h
    port map (
            O => \N__29413\,
            I => \N__29404\
        );

    \I__4397\ : Span12Mux_v
    port map (
            O => \N__29410\,
            I => \N__29401\
        );

    \I__4396\ : Odrv4
    port map (
            O => \N__29407\,
            I => n2630
        );

    \I__4395\ : Odrv4
    port map (
            O => \N__29404\,
            I => n2630
        );

    \I__4394\ : Odrv12
    port map (
            O => \N__29401\,
            I => n2630
        );

    \I__4393\ : CascadeMux
    port map (
            O => \N__29394\,
            I => \N__29391\
        );

    \I__4392\ : InMux
    port map (
            O => \N__29391\,
            I => \N__29388\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__29388\,
            I => \N__29384\
        );

    \I__4390\ : InMux
    port map (
            O => \N__29387\,
            I => \N__29380\
        );

    \I__4389\ : Span4Mux_h
    port map (
            O => \N__29384\,
            I => \N__29377\
        );

    \I__4388\ : InMux
    port map (
            O => \N__29383\,
            I => \N__29374\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__29380\,
            I => \N__29371\
        );

    \I__4386\ : Span4Mux_v
    port map (
            O => \N__29377\,
            I => \N__29368\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__29374\,
            I => \N__29365\
        );

    \I__4384\ : Span4Mux_h
    port map (
            O => \N__29371\,
            I => \N__29362\
        );

    \I__4383\ : Span4Mux_v
    port map (
            O => \N__29368\,
            I => \N__29357\
        );

    \I__4382\ : Span4Mux_h
    port map (
            O => \N__29365\,
            I => \N__29357\
        );

    \I__4381\ : Odrv4
    port map (
            O => \N__29362\,
            I => n2620
        );

    \I__4380\ : Odrv4
    port map (
            O => \N__29357\,
            I => n2620
        );

    \I__4379\ : InMux
    port map (
            O => \N__29352\,
            I => \N__29349\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__29349\,
            I => \N__29346\
        );

    \I__4377\ : Span4Mux_v
    port map (
            O => \N__29346\,
            I => \N__29343\
        );

    \I__4376\ : Odrv4
    port map (
            O => \N__29343\,
            I => n2901
        );

    \I__4375\ : InMux
    port map (
            O => \N__29340\,
            I => \N__29337\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__29337\,
            I => \N__29333\
        );

    \I__4373\ : CascadeMux
    port map (
            O => \N__29336\,
            I => \N__29330\
        );

    \I__4372\ : Span4Mux_h
    port map (
            O => \N__29333\,
            I => \N__29326\
        );

    \I__4371\ : InMux
    port map (
            O => \N__29330\,
            I => \N__29323\
        );

    \I__4370\ : InMux
    port map (
            O => \N__29329\,
            I => \N__29320\
        );

    \I__4369\ : Odrv4
    port map (
            O => \N__29326\,
            I => n2824
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__29323\,
            I => n2824
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__29320\,
            I => n2824
        );

    \I__4366\ : InMux
    port map (
            O => \N__29313\,
            I => \N__29310\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__29310\,
            I => \N__29307\
        );

    \I__4364\ : Span4Mux_h
    port map (
            O => \N__29307\,
            I => \N__29304\
        );

    \I__4363\ : Odrv4
    port map (
            O => \N__29304\,
            I => n2891
        );

    \I__4362\ : InMux
    port map (
            O => \N__29301\,
            I => \N__29297\
        );

    \I__4361\ : CascadeMux
    port map (
            O => \N__29300\,
            I => \N__29294\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__29297\,
            I => \N__29291\
        );

    \I__4359\ : InMux
    port map (
            O => \N__29294\,
            I => \N__29288\
        );

    \I__4358\ : Span12Mux_s6_v
    port map (
            O => \N__29291\,
            I => \N__29283\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__29288\,
            I => \N__29283\
        );

    \I__4356\ : Odrv12
    port map (
            O => \N__29283\,
            I => n2923
        );

    \I__4355\ : CascadeMux
    port map (
            O => \N__29280\,
            I => \n2923_cascade_\
        );

    \I__4354\ : InMux
    port map (
            O => \N__29277\,
            I => \N__29274\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__29274\,
            I => n14214
        );

    \I__4352\ : CascadeMux
    port map (
            O => \N__29271\,
            I => \n2533_cascade_\
        );

    \I__4351\ : CascadeMux
    port map (
            O => \N__29268\,
            I => \N__29265\
        );

    \I__4350\ : InMux
    port map (
            O => \N__29265\,
            I => \N__29262\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__29262\,
            I => n12063
        );

    \I__4348\ : CascadeMux
    port map (
            O => \N__29259\,
            I => \N__29256\
        );

    \I__4347\ : InMux
    port map (
            O => \N__29256\,
            I => \N__29253\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__29253\,
            I => \N__29249\
        );

    \I__4345\ : InMux
    port map (
            O => \N__29252\,
            I => \N__29246\
        );

    \I__4344\ : Span4Mux_h
    port map (
            O => \N__29249\,
            I => \N__29243\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__29246\,
            I => \N__29240\
        );

    \I__4342\ : Span4Mux_v
    port map (
            O => \N__29243\,
            I => \N__29236\
        );

    \I__4341\ : Span12Mux_s4_h
    port map (
            O => \N__29240\,
            I => \N__29233\
        );

    \I__4340\ : InMux
    port map (
            O => \N__29239\,
            I => \N__29230\
        );

    \I__4339\ : Span4Mux_v
    port map (
            O => \N__29236\,
            I => \N__29227\
        );

    \I__4338\ : Odrv12
    port map (
            O => \N__29233\,
            I => n2632
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__29230\,
            I => n2632
        );

    \I__4336\ : Odrv4
    port map (
            O => \N__29227\,
            I => n2632
        );

    \I__4335\ : InMux
    port map (
            O => \N__29220\,
            I => \N__29217\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__29217\,
            I => n14188
        );

    \I__4333\ : CascadeMux
    port map (
            O => \N__29214\,
            I => \n2515_cascade_\
        );

    \I__4332\ : InMux
    port map (
            O => \N__29211\,
            I => \N__29208\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__29208\,
            I => \N__29205\
        );

    \I__4330\ : Odrv4
    port map (
            O => \N__29205\,
            I => n14117
        );

    \I__4329\ : CascadeMux
    port map (
            O => \N__29202\,
            I => \n14194_cascade_\
        );

    \I__4328\ : CascadeMux
    port map (
            O => \N__29199\,
            I => \n2544_cascade_\
        );

    \I__4327\ : CascadeMux
    port map (
            O => \N__29196\,
            I => \N__29192\
        );

    \I__4326\ : InMux
    port map (
            O => \N__29195\,
            I => \N__29189\
        );

    \I__4325\ : InMux
    port map (
            O => \N__29192\,
            I => \N__29186\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__29189\,
            I => \N__29183\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__29186\,
            I => \N__29179\
        );

    \I__4322\ : Span4Mux_v
    port map (
            O => \N__29183\,
            I => \N__29176\
        );

    \I__4321\ : InMux
    port map (
            O => \N__29182\,
            I => \N__29173\
        );

    \I__4320\ : Span12Mux_v
    port map (
            O => \N__29179\,
            I => \N__29170\
        );

    \I__4319\ : Odrv4
    port map (
            O => \N__29176\,
            I => n2631
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__29173\,
            I => n2631
        );

    \I__4317\ : Odrv12
    port map (
            O => \N__29170\,
            I => n2631
        );

    \I__4316\ : CascadeMux
    port map (
            O => \N__29163\,
            I => \n2417_cascade_\
        );

    \I__4315\ : InMux
    port map (
            O => \N__29160\,
            I => \N__29157\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__29157\,
            I => n14634
        );

    \I__4313\ : CascadeMux
    port map (
            O => \N__29154\,
            I => \n14640_cascade_\
        );

    \I__4312\ : CascadeMux
    port map (
            O => \N__29151\,
            I => \n2445_cascade_\
        );

    \I__4311\ : CascadeMux
    port map (
            O => \N__29148\,
            I => \n2530_cascade_\
        );

    \I__4310\ : InMux
    port map (
            O => \N__29145\,
            I => \N__29142\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__29142\,
            I => n14646
        );

    \I__4308\ : CascadeMux
    port map (
            O => \N__29139\,
            I => \n2430_cascade_\
        );

    \I__4307\ : InMux
    port map (
            O => \N__29136\,
            I => \N__29133\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__29133\,
            I => \N__29130\
        );

    \I__4305\ : Span4Mux_v
    port map (
            O => \N__29130\,
            I => \N__29127\
        );

    \I__4304\ : Odrv4
    port map (
            O => \N__29127\,
            I => n2400
        );

    \I__4303\ : CascadeMux
    port map (
            O => \N__29124\,
            I => \N__29120\
        );

    \I__4302\ : CascadeMux
    port map (
            O => \N__29123\,
            I => \N__29117\
        );

    \I__4301\ : InMux
    port map (
            O => \N__29120\,
            I => \N__29114\
        );

    \I__4300\ : InMux
    port map (
            O => \N__29117\,
            I => \N__29111\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__29114\,
            I => \N__29108\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__29111\,
            I => \N__29105\
        );

    \I__4297\ : Span4Mux_v
    port map (
            O => \N__29108\,
            I => \N__29101\
        );

    \I__4296\ : Span4Mux_s2_h
    port map (
            O => \N__29105\,
            I => \N__29098\
        );

    \I__4295\ : InMux
    port map (
            O => \N__29104\,
            I => \N__29095\
        );

    \I__4294\ : Odrv4
    port map (
            O => \N__29101\,
            I => n2333
        );

    \I__4293\ : Odrv4
    port map (
            O => \N__29098\,
            I => n2333
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__29095\,
            I => n2333
        );

    \I__4291\ : CascadeMux
    port map (
            O => \N__29088\,
            I => \n2432_cascade_\
        );

    \I__4290\ : InMux
    port map (
            O => \N__29085\,
            I => \N__29082\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__29082\,
            I => n11967
        );

    \I__4288\ : CascadeMux
    port map (
            O => \N__29079\,
            I => \n2528_cascade_\
        );

    \I__4287\ : CascadeMux
    port map (
            O => \N__29076\,
            I => \N__29073\
        );

    \I__4286\ : InMux
    port map (
            O => \N__29073\,
            I => \N__29070\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__29070\,
            I => \N__29066\
        );

    \I__4284\ : InMux
    port map (
            O => \N__29069\,
            I => \N__29063\
        );

    \I__4283\ : Span4Mux_h
    port map (
            O => \N__29066\,
            I => \N__29060\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__29063\,
            I => \N__29056\
        );

    \I__4281\ : Span4Mux_v
    port map (
            O => \N__29060\,
            I => \N__29053\
        );

    \I__4280\ : InMux
    port map (
            O => \N__29059\,
            I => \N__29050\
        );

    \I__4279\ : Span4Mux_h
    port map (
            O => \N__29056\,
            I => \N__29045\
        );

    \I__4278\ : Span4Mux_v
    port map (
            O => \N__29053\,
            I => \N__29045\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__29050\,
            I => n2627
        );

    \I__4276\ : Odrv4
    port map (
            O => \N__29045\,
            I => n2627
        );

    \I__4275\ : InMux
    port map (
            O => \N__29040\,
            I => \N__29037\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__29037\,
            I => \N__29034\
        );

    \I__4273\ : Span4Mux_h
    port map (
            O => \N__29034\,
            I => \N__29031\
        );

    \I__4272\ : Odrv4
    port map (
            O => \N__29031\,
            I => n2384
        );

    \I__4271\ : CascadeMux
    port map (
            O => \N__29028\,
            I => \N__29025\
        );

    \I__4270\ : InMux
    port map (
            O => \N__29025\,
            I => \N__29021\
        );

    \I__4269\ : InMux
    port map (
            O => \N__29024\,
            I => \N__29018\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__29021\,
            I => \N__29014\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__29018\,
            I => \N__29011\
        );

    \I__4266\ : CascadeMux
    port map (
            O => \N__29017\,
            I => \N__29008\
        );

    \I__4265\ : Span4Mux_h
    port map (
            O => \N__29014\,
            I => \N__29005\
        );

    \I__4264\ : Span4Mux_s3_h
    port map (
            O => \N__29011\,
            I => \N__29002\
        );

    \I__4263\ : InMux
    port map (
            O => \N__29008\,
            I => \N__28999\
        );

    \I__4262\ : Odrv4
    port map (
            O => \N__29005\,
            I => n2317
        );

    \I__4261\ : Odrv4
    port map (
            O => \N__29002\,
            I => n2317
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__28999\,
            I => n2317
        );

    \I__4259\ : InMux
    port map (
            O => \N__28992\,
            I => \N__28989\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__28989\,
            I => n13828
        );

    \I__4257\ : InMux
    port map (
            O => \N__28986\,
            I => \N__28983\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__28983\,
            I => n14628
        );

    \I__4255\ : InMux
    port map (
            O => \N__28980\,
            I => \N__28976\
        );

    \I__4254\ : InMux
    port map (
            O => \N__28979\,
            I => \N__28973\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__28976\,
            I => \N__28969\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__28973\,
            I => \N__28966\
        );

    \I__4251\ : InMux
    port map (
            O => \N__28972\,
            I => \N__28963\
        );

    \I__4250\ : Span4Mux_v
    port map (
            O => \N__28969\,
            I => \N__28960\
        );

    \I__4249\ : Span4Mux_s2_h
    port map (
            O => \N__28966\,
            I => \N__28957\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__28963\,
            I => \N__28954\
        );

    \I__4247\ : Odrv4
    port map (
            O => \N__28960\,
            I => n2318
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__28957\,
            I => n2318
        );

    \I__4245\ : Odrv4
    port map (
            O => \N__28954\,
            I => n2318
        );

    \I__4244\ : CascadeMux
    port map (
            O => \N__28947\,
            I => \N__28944\
        );

    \I__4243\ : InMux
    port map (
            O => \N__28944\,
            I => \N__28941\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__28941\,
            I => \N__28938\
        );

    \I__4241\ : Span4Mux_h
    port map (
            O => \N__28938\,
            I => \N__28935\
        );

    \I__4240\ : Odrv4
    port map (
            O => \N__28935\,
            I => n2385
        );

    \I__4239\ : InMux
    port map (
            O => \N__28932\,
            I => \N__28929\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__28929\,
            I => \N__28926\
        );

    \I__4237\ : Odrv12
    port map (
            O => \N__28926\,
            I => n2390
        );

    \I__4236\ : CascadeMux
    port map (
            O => \N__28923\,
            I => \N__28919\
        );

    \I__4235\ : CascadeMux
    port map (
            O => \N__28922\,
            I => \N__28916\
        );

    \I__4234\ : InMux
    port map (
            O => \N__28919\,
            I => \N__28913\
        );

    \I__4233\ : InMux
    port map (
            O => \N__28916\,
            I => \N__28910\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__28913\,
            I => \N__28907\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__28910\,
            I => \N__28904\
        );

    \I__4230\ : Span4Mux_v
    port map (
            O => \N__28907\,
            I => \N__28899\
        );

    \I__4229\ : Span4Mux_v
    port map (
            O => \N__28904\,
            I => \N__28899\
        );

    \I__4228\ : Odrv4
    port map (
            O => \N__28899\,
            I => n2323
        );

    \I__4227\ : CascadeMux
    port map (
            O => \N__28896\,
            I => \N__28892\
        );

    \I__4226\ : InMux
    port map (
            O => \N__28895\,
            I => \N__28888\
        );

    \I__4225\ : InMux
    port map (
            O => \N__28892\,
            I => \N__28885\
        );

    \I__4224\ : InMux
    port map (
            O => \N__28891\,
            I => \N__28882\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__28888\,
            I => \N__28879\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__28885\,
            I => n2118
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__28882\,
            I => n2118
        );

    \I__4220\ : Odrv4
    port map (
            O => \N__28879\,
            I => n2118
        );

    \I__4219\ : InMux
    port map (
            O => \N__28872\,
            I => \N__28869\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__28869\,
            I => \N__28866\
        );

    \I__4217\ : Odrv12
    port map (
            O => \N__28866\,
            I => n2393
        );

    \I__4216\ : CascadeMux
    port map (
            O => \N__28863\,
            I => \N__28860\
        );

    \I__4215\ : InMux
    port map (
            O => \N__28860\,
            I => \N__28856\
        );

    \I__4214\ : CascadeMux
    port map (
            O => \N__28859\,
            I => \N__28853\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__28856\,
            I => \N__28850\
        );

    \I__4212\ : InMux
    port map (
            O => \N__28853\,
            I => \N__28846\
        );

    \I__4211\ : Span4Mux_v
    port map (
            O => \N__28850\,
            I => \N__28843\
        );

    \I__4210\ : InMux
    port map (
            O => \N__28849\,
            I => \N__28840\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__28846\,
            I => n2326
        );

    \I__4208\ : Odrv4
    port map (
            O => \N__28843\,
            I => n2326
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__28840\,
            I => n2326
        );

    \I__4206\ : InMux
    port map (
            O => \N__28833\,
            I => \N__28828\
        );

    \I__4205\ : CascadeMux
    port map (
            O => \N__28832\,
            I => \N__28825\
        );

    \I__4204\ : CascadeMux
    port map (
            O => \N__28831\,
            I => \N__28822\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__28828\,
            I => \N__28819\
        );

    \I__4202\ : InMux
    port map (
            O => \N__28825\,
            I => \N__28816\
        );

    \I__4201\ : InMux
    port map (
            O => \N__28822\,
            I => \N__28813\
        );

    \I__4200\ : Span4Mux_v
    port map (
            O => \N__28819\,
            I => \N__28808\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__28816\,
            I => \N__28808\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__28813\,
            I => n2330
        );

    \I__4197\ : Odrv4
    port map (
            O => \N__28808\,
            I => n2330
        );

    \I__4196\ : InMux
    port map (
            O => \N__28803\,
            I => \N__28800\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__28800\,
            I => \N__28797\
        );

    \I__4194\ : Span12Mux_v
    port map (
            O => \N__28797\,
            I => \N__28794\
        );

    \I__4193\ : Odrv12
    port map (
            O => \N__28794\,
            I => n2397
        );

    \I__4192\ : CascadeMux
    port map (
            O => \N__28791\,
            I => \N__28787\
        );

    \I__4191\ : InMux
    port map (
            O => \N__28790\,
            I => \N__28784\
        );

    \I__4190\ : InMux
    port map (
            O => \N__28787\,
            I => \N__28781\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__28784\,
            I => \N__28778\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__28781\,
            I => \N__28775\
        );

    \I__4187\ : Span4Mux_h
    port map (
            O => \N__28778\,
            I => \N__28769\
        );

    \I__4186\ : Span4Mux_s2_h
    port map (
            O => \N__28775\,
            I => \N__28769\
        );

    \I__4185\ : InMux
    port map (
            O => \N__28774\,
            I => \N__28766\
        );

    \I__4184\ : Odrv4
    port map (
            O => \N__28769\,
            I => n2322
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__28766\,
            I => n2322
        );

    \I__4182\ : CascadeMux
    port map (
            O => \N__28761\,
            I => \N__28758\
        );

    \I__4181\ : InMux
    port map (
            O => \N__28758\,
            I => \N__28755\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__28755\,
            I => \N__28752\
        );

    \I__4179\ : Odrv12
    port map (
            O => \N__28752\,
            I => n2389
        );

    \I__4178\ : InMux
    port map (
            O => \N__28749\,
            I => \N__28746\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__28746\,
            I => \N__28743\
        );

    \I__4176\ : Span4Mux_v
    port map (
            O => \N__28743\,
            I => \N__28740\
        );

    \I__4175\ : Odrv4
    port map (
            O => \N__28740\,
            I => n2399
        );

    \I__4174\ : CascadeMux
    port map (
            O => \N__28737\,
            I => \N__28733\
        );

    \I__4173\ : InMux
    port map (
            O => \N__28736\,
            I => \N__28730\
        );

    \I__4172\ : InMux
    port map (
            O => \N__28733\,
            I => \N__28727\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__28730\,
            I => \N__28724\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__28727\,
            I => \N__28721\
        );

    \I__4169\ : Span4Mux_v
    port map (
            O => \N__28724\,
            I => \N__28717\
        );

    \I__4168\ : Span4Mux_s2_h
    port map (
            O => \N__28721\,
            I => \N__28714\
        );

    \I__4167\ : InMux
    port map (
            O => \N__28720\,
            I => \N__28711\
        );

    \I__4166\ : Odrv4
    port map (
            O => \N__28717\,
            I => n2332
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__28714\,
            I => n2332
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__28711\,
            I => n2332
        );

    \I__4163\ : InMux
    port map (
            O => \N__28704\,
            I => \N__28701\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__28701\,
            I => \N__28698\
        );

    \I__4161\ : Span4Mux_v
    port map (
            O => \N__28698\,
            I => \N__28695\
        );

    \I__4160\ : Odrv4
    port map (
            O => \N__28695\,
            I => n2388
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__28692\,
            I => \N__28689\
        );

    \I__4158\ : InMux
    port map (
            O => \N__28689\,
            I => \N__28685\
        );

    \I__4157\ : InMux
    port map (
            O => \N__28688\,
            I => \N__28682\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__28685\,
            I => \N__28678\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__28682\,
            I => \N__28675\
        );

    \I__4154\ : InMux
    port map (
            O => \N__28681\,
            I => \N__28672\
        );

    \I__4153\ : Span4Mux_v
    port map (
            O => \N__28678\,
            I => \N__28669\
        );

    \I__4152\ : Span4Mux_s3_h
    port map (
            O => \N__28675\,
            I => \N__28664\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__28672\,
            I => \N__28664\
        );

    \I__4150\ : Odrv4
    port map (
            O => \N__28669\,
            I => n2321
        );

    \I__4149\ : Odrv4
    port map (
            O => \N__28664\,
            I => n2321
        );

    \I__4148\ : CascadeMux
    port map (
            O => \N__28659\,
            I => \n2420_cascade_\
        );

    \I__4147\ : InMux
    port map (
            O => \N__28656\,
            I => \N__28653\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__28653\,
            I => n14622
        );

    \I__4145\ : InMux
    port map (
            O => \N__28650\,
            I => \N__28647\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__28647\,
            I => \N__28644\
        );

    \I__4143\ : Span4Mux_v
    port map (
            O => \N__28644\,
            I => \N__28641\
        );

    \I__4142\ : Odrv4
    port map (
            O => \N__28641\,
            I => n2398
        );

    \I__4141\ : CascadeMux
    port map (
            O => \N__28638\,
            I => \N__28634\
        );

    \I__4140\ : CascadeMux
    port map (
            O => \N__28637\,
            I => \N__28631\
        );

    \I__4139\ : InMux
    port map (
            O => \N__28634\,
            I => \N__28628\
        );

    \I__4138\ : InMux
    port map (
            O => \N__28631\,
            I => \N__28625\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__28628\,
            I => \N__28622\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__28625\,
            I => \N__28619\
        );

    \I__4135\ : Span4Mux_v
    port map (
            O => \N__28622\,
            I => \N__28614\
        );

    \I__4134\ : Span4Mux_v
    port map (
            O => \N__28619\,
            I => \N__28614\
        );

    \I__4133\ : Odrv4
    port map (
            O => \N__28614\,
            I => n2331
        );

    \I__4132\ : CascadeMux
    port map (
            O => \N__28611\,
            I => \N__28608\
        );

    \I__4131\ : InMux
    port map (
            O => \N__28608\,
            I => \N__28604\
        );

    \I__4130\ : CascadeMux
    port map (
            O => \N__28607\,
            I => \N__28601\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__28604\,
            I => \N__28597\
        );

    \I__4128\ : InMux
    port map (
            O => \N__28601\,
            I => \N__28594\
        );

    \I__4127\ : InMux
    port map (
            O => \N__28600\,
            I => \N__28591\
        );

    \I__4126\ : Odrv4
    port map (
            O => \N__28597\,
            I => n2126
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__28594\,
            I => n2126
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__28591\,
            I => n2126
        );

    \I__4123\ : CascadeMux
    port map (
            O => \N__28584\,
            I => \n2128_cascade_\
        );

    \I__4122\ : InMux
    port map (
            O => \N__28581\,
            I => \N__28578\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__28578\,
            I => n14316
        );

    \I__4120\ : CascadeMux
    port map (
            O => \N__28575\,
            I => \N__28570\
        );

    \I__4119\ : CascadeMux
    port map (
            O => \N__28574\,
            I => \N__28567\
        );

    \I__4118\ : InMux
    port map (
            O => \N__28573\,
            I => \N__28564\
        );

    \I__4117\ : InMux
    port map (
            O => \N__28570\,
            I => \N__28561\
        );

    \I__4116\ : InMux
    port map (
            O => \N__28567\,
            I => \N__28558\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__28564\,
            I => \N__28555\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__28561\,
            I => n2125
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__28558\,
            I => n2125
        );

    \I__4112\ : Odrv4
    port map (
            O => \N__28555\,
            I => n2125
        );

    \I__4111\ : InMux
    port map (
            O => \N__28548\,
            I => \N__28545\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__28545\,
            I => \N__28542\
        );

    \I__4109\ : Odrv4
    port map (
            O => \N__28542\,
            I => n2185
        );

    \I__4108\ : CascadeMux
    port map (
            O => \N__28539\,
            I => \N__28536\
        );

    \I__4107\ : InMux
    port map (
            O => \N__28536\,
            I => \N__28532\
        );

    \I__4106\ : CascadeMux
    port map (
            O => \N__28535\,
            I => \N__28528\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__28532\,
            I => \N__28525\
        );

    \I__4104\ : InMux
    port map (
            O => \N__28531\,
            I => \N__28522\
        );

    \I__4103\ : InMux
    port map (
            O => \N__28528\,
            I => \N__28519\
        );

    \I__4102\ : Span4Mux_h
    port map (
            O => \N__28525\,
            I => \N__28516\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__28522\,
            I => \N__28513\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__28519\,
            I => n2217
        );

    \I__4099\ : Odrv4
    port map (
            O => \N__28516\,
            I => n2217
        );

    \I__4098\ : Odrv4
    port map (
            O => \N__28513\,
            I => n2217
        );

    \I__4097\ : InMux
    port map (
            O => \N__28506\,
            I => \N__28503\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__28503\,
            I => n2183
        );

    \I__4095\ : InMux
    port map (
            O => \N__28500\,
            I => \N__28496\
        );

    \I__4094\ : InMux
    port map (
            O => \N__28499\,
            I => \N__28493\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__28496\,
            I => n2116
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__28493\,
            I => n2116
        );

    \I__4091\ : InMux
    port map (
            O => \N__28488\,
            I => \N__28485\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__28485\,
            I => \N__28480\
        );

    \I__4089\ : InMux
    port map (
            O => \N__28484\,
            I => \N__28477\
        );

    \I__4088\ : InMux
    port map (
            O => \N__28483\,
            I => \N__28474\
        );

    \I__4087\ : Span4Mux_h
    port map (
            O => \N__28480\,
            I => \N__28471\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__28477\,
            I => \N__28468\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__28474\,
            I => n2215
        );

    \I__4084\ : Odrv4
    port map (
            O => \N__28471\,
            I => n2215
        );

    \I__4083\ : Odrv4
    port map (
            O => \N__28468\,
            I => n2215
        );

    \I__4082\ : InMux
    port map (
            O => \N__28461\,
            I => \N__28458\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__28458\,
            I => n2184
        );

    \I__4080\ : InMux
    port map (
            O => \N__28455\,
            I => \N__28452\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__28452\,
            I => \N__28447\
        );

    \I__4078\ : CascadeMux
    port map (
            O => \N__28451\,
            I => \N__28444\
        );

    \I__4077\ : InMux
    port map (
            O => \N__28450\,
            I => \N__28441\
        );

    \I__4076\ : Span4Mux_v
    port map (
            O => \N__28447\,
            I => \N__28438\
        );

    \I__4075\ : InMux
    port map (
            O => \N__28444\,
            I => \N__28435\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__28441\,
            I => \N__28432\
        );

    \I__4073\ : Odrv4
    port map (
            O => \N__28438\,
            I => n2122
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__28435\,
            I => n2122
        );

    \I__4071\ : Odrv4
    port map (
            O => \N__28432\,
            I => n2122
        );

    \I__4070\ : CascadeMux
    port map (
            O => \N__28425\,
            I => \N__28422\
        );

    \I__4069\ : InMux
    port map (
            O => \N__28422\,
            I => \N__28417\
        );

    \I__4068\ : InMux
    port map (
            O => \N__28421\,
            I => \N__28412\
        );

    \I__4067\ : InMux
    port map (
            O => \N__28420\,
            I => \N__28412\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__28417\,
            I => n2124
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__28412\,
            I => n2124
        );

    \I__4064\ : InMux
    port map (
            O => \N__28407\,
            I => \N__28404\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__28404\,
            I => \N__28401\
        );

    \I__4062\ : Span4Mux_h
    port map (
            O => \N__28401\,
            I => \N__28398\
        );

    \I__4061\ : Odrv4
    port map (
            O => \N__28398\,
            I => n2401
        );

    \I__4060\ : InMux
    port map (
            O => \N__28395\,
            I => \N__28392\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__28392\,
            I => n2198
        );

    \I__4058\ : CascadeMux
    port map (
            O => \N__28389\,
            I => \n2131_cascade_\
        );

    \I__4057\ : CascadeMux
    port map (
            O => \N__28386\,
            I => \N__28381\
        );

    \I__4056\ : InMux
    port map (
            O => \N__28385\,
            I => \N__28376\
        );

    \I__4055\ : InMux
    port map (
            O => \N__28384\,
            I => \N__28376\
        );

    \I__4054\ : InMux
    port map (
            O => \N__28381\,
            I => \N__28373\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__28376\,
            I => \N__28370\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__28373\,
            I => \N__28367\
        );

    \I__4051\ : Span4Mux_h
    port map (
            O => \N__28370\,
            I => \N__28364\
        );

    \I__4050\ : Span4Mux_h
    port map (
            O => \N__28367\,
            I => \N__28361\
        );

    \I__4049\ : Odrv4
    port map (
            O => \N__28364\,
            I => n2230
        );

    \I__4048\ : Odrv4
    port map (
            O => \N__28361\,
            I => n2230
        );

    \I__4047\ : InMux
    port map (
            O => \N__28356\,
            I => \N__28353\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__28353\,
            I => n14584
        );

    \I__4045\ : CascadeMux
    port map (
            O => \N__28350\,
            I => \N__28347\
        );

    \I__4044\ : InMux
    port map (
            O => \N__28347\,
            I => \N__28344\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__28344\,
            I => n2191
        );

    \I__4042\ : CascadeMux
    port map (
            O => \N__28341\,
            I => \N__28337\
        );

    \I__4041\ : CascadeMux
    port map (
            O => \N__28340\,
            I => \N__28333\
        );

    \I__4040\ : InMux
    port map (
            O => \N__28337\,
            I => \N__28330\
        );

    \I__4039\ : InMux
    port map (
            O => \N__28336\,
            I => \N__28327\
        );

    \I__4038\ : InMux
    port map (
            O => \N__28333\,
            I => \N__28324\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__28330\,
            I => \N__28319\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__28327\,
            I => \N__28319\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__28324\,
            I => \N__28314\
        );

    \I__4034\ : Span4Mux_v
    port map (
            O => \N__28319\,
            I => \N__28314\
        );

    \I__4033\ : Odrv4
    port map (
            O => \N__28314\,
            I => n2223
        );

    \I__4032\ : InMux
    port map (
            O => \N__28311\,
            I => \N__28308\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__28308\,
            I => n2192
        );

    \I__4030\ : CascadeMux
    port map (
            O => \N__28305\,
            I => \N__28301\
        );

    \I__4029\ : CascadeMux
    port map (
            O => \N__28304\,
            I => \N__28298\
        );

    \I__4028\ : InMux
    port map (
            O => \N__28301\,
            I => \N__28295\
        );

    \I__4027\ : InMux
    port map (
            O => \N__28298\,
            I => \N__28292\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__28295\,
            I => \N__28289\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__28292\,
            I => \N__28285\
        );

    \I__4024\ : Span4Mux_h
    port map (
            O => \N__28289\,
            I => \N__28282\
        );

    \I__4023\ : InMux
    port map (
            O => \N__28288\,
            I => \N__28279\
        );

    \I__4022\ : Odrv4
    port map (
            O => \N__28285\,
            I => n2224
        );

    \I__4021\ : Odrv4
    port map (
            O => \N__28282\,
            I => n2224
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__28279\,
            I => n2224
        );

    \I__4019\ : InMux
    port map (
            O => \N__28272\,
            I => \N__28269\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__28269\,
            I => n14330
        );

    \I__4017\ : CascadeMux
    port map (
            O => \N__28266\,
            I => \n2116_cascade_\
        );

    \I__4016\ : CascadeMux
    port map (
            O => \N__28263\,
            I => \n2148_cascade_\
        );

    \I__4015\ : InMux
    port map (
            O => \N__28260\,
            I => \N__28257\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__28257\,
            I => n2195
        );

    \I__4013\ : CascadeMux
    port map (
            O => \N__28254\,
            I => \N__28251\
        );

    \I__4012\ : InMux
    port map (
            O => \N__28251\,
            I => \N__28248\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__28248\,
            I => \N__28243\
        );

    \I__4010\ : CascadeMux
    port map (
            O => \N__28247\,
            I => \N__28240\
        );

    \I__4009\ : InMux
    port map (
            O => \N__28246\,
            I => \N__28237\
        );

    \I__4008\ : Span4Mux_h
    port map (
            O => \N__28243\,
            I => \N__28234\
        );

    \I__4007\ : InMux
    port map (
            O => \N__28240\,
            I => \N__28231\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__28237\,
            I => n2227
        );

    \I__4005\ : Odrv4
    port map (
            O => \N__28234\,
            I => n2227
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__28231\,
            I => n2227
        );

    \I__4003\ : CascadeMux
    port map (
            O => \N__28224\,
            I => \N__28220\
        );

    \I__4002\ : InMux
    port map (
            O => \N__28223\,
            I => \N__28217\
        );

    \I__4001\ : InMux
    port map (
            O => \N__28220\,
            I => \N__28214\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__28217\,
            I => n2128
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__28214\,
            I => n2128
        );

    \I__3998\ : InMux
    port map (
            O => \N__28209\,
            I => \N__28205\
        );

    \I__3997\ : InMux
    port map (
            O => \N__28208\,
            I => \N__28202\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__28205\,
            I => \N__28197\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__28202\,
            I => \N__28197\
        );

    \I__3994\ : Span4Mux_s3_v
    port map (
            O => \N__28197\,
            I => \N__28193\
        );

    \I__3993\ : InMux
    port map (
            O => \N__28196\,
            I => \N__28190\
        );

    \I__3992\ : Odrv4
    port map (
            O => \N__28193\,
            I => n3010
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__28190\,
            I => n3010
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__28185\,
            I => \N__28182\
        );

    \I__3989\ : InMux
    port map (
            O => \N__28182\,
            I => \N__28179\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__28179\,
            I => n3077
        );

    \I__3987\ : InMux
    port map (
            O => \N__28176\,
            I => \N__28173\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__28173\,
            I => \N__28170\
        );

    \I__3985\ : Odrv4
    port map (
            O => \N__28170\,
            I => n14264
        );

    \I__3984\ : CascadeMux
    port map (
            O => \N__28167\,
            I => \N__28164\
        );

    \I__3983\ : InMux
    port map (
            O => \N__28164\,
            I => \N__28161\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__28161\,
            I => \N__28158\
        );

    \I__3981\ : Odrv4
    port map (
            O => \N__28158\,
            I => n14260
        );

    \I__3980\ : CascadeMux
    port map (
            O => \N__28155\,
            I => \N__28152\
        );

    \I__3979\ : InMux
    port map (
            O => \N__28152\,
            I => \N__28147\
        );

    \I__3978\ : InMux
    port map (
            O => \N__28151\,
            I => \N__28142\
        );

    \I__3977\ : InMux
    port map (
            O => \N__28150\,
            I => \N__28142\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__28147\,
            I => n2130
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__28142\,
            I => n2130
        );

    \I__3974\ : CascadeMux
    port map (
            O => \N__28137\,
            I => \n14324_cascade_\
        );

    \I__3973\ : InMux
    port map (
            O => \N__28134\,
            I => \N__28131\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__28131\,
            I => n13787
        );

    \I__3971\ : CascadeMux
    port map (
            O => \N__28128\,
            I => \N__28124\
        );

    \I__3970\ : CascadeMux
    port map (
            O => \N__28127\,
            I => \N__28121\
        );

    \I__3969\ : InMux
    port map (
            O => \N__28124\,
            I => \N__28118\
        );

    \I__3968\ : InMux
    port map (
            O => \N__28121\,
            I => \N__28115\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__28118\,
            I => n2127
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__28115\,
            I => n2127
        );

    \I__3965\ : CascadeMux
    port map (
            O => \N__28110\,
            I => \n2127_cascade_\
        );

    \I__3964\ : InMux
    port map (
            O => \N__28107\,
            I => \N__28104\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__28104\,
            I => n14318
        );

    \I__3962\ : CascadeMux
    port map (
            O => \N__28101\,
            I => \N__28098\
        );

    \I__3961\ : InMux
    port map (
            O => \N__28098\,
            I => \N__28094\
        );

    \I__3960\ : InMux
    port map (
            O => \N__28097\,
            I => \N__28091\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__28094\,
            I => n2131
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__28091\,
            I => n2131
        );

    \I__3957\ : CascadeMux
    port map (
            O => \N__28086\,
            I => \n3212_cascade_\
        );

    \I__3956\ : InMux
    port map (
            O => \N__28083\,
            I => \N__28080\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__28080\,
            I => n14798
        );

    \I__3954\ : InMux
    port map (
            O => \N__28077\,
            I => \N__28072\
        );

    \I__3953\ : InMux
    port map (
            O => \N__28076\,
            I => \N__28069\
        );

    \I__3952\ : InMux
    port map (
            O => \N__28075\,
            I => \N__28066\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__28072\,
            I => n3107
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__28069\,
            I => n3107
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__28066\,
            I => n3107
        );

    \I__3948\ : InMux
    port map (
            O => \N__28059\,
            I => \N__28054\
        );

    \I__3947\ : InMux
    port map (
            O => \N__28058\,
            I => \N__28051\
        );

    \I__3946\ : InMux
    port map (
            O => \N__28057\,
            I => \N__28048\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__28054\,
            I => n3106
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__28051\,
            I => n3106
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__28048\,
            I => n3106
        );

    \I__3942\ : CascadeMux
    port map (
            O => \N__28041\,
            I => \N__28037\
        );

    \I__3941\ : InMux
    port map (
            O => \N__28040\,
            I => \N__28034\
        );

    \I__3940\ : InMux
    port map (
            O => \N__28037\,
            I => \N__28031\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__28034\,
            I => n3105
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__28031\,
            I => n3105
        );

    \I__3937\ : InMux
    port map (
            O => \N__28026\,
            I => \N__28023\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__28023\,
            I => \N__28020\
        );

    \I__3935\ : Span4Mux_h
    port map (
            O => \N__28020\,
            I => \N__28017\
        );

    \I__3934\ : Odrv4
    port map (
            O => \N__28017\,
            I => n3195
        );

    \I__3933\ : CascadeMux
    port map (
            O => \N__28014\,
            I => \n3138_cascade_\
        );

    \I__3932\ : InMux
    port map (
            O => \N__28011\,
            I => \N__28008\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__28008\,
            I => \N__28004\
        );

    \I__3930\ : CascadeMux
    port map (
            O => \N__28007\,
            I => \N__28001\
        );

    \I__3929\ : Span4Mux_h
    port map (
            O => \N__28004\,
            I => \N__27998\
        );

    \I__3928\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27995\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__27998\,
            I => n3128
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__27995\,
            I => n3128
        );

    \I__3925\ : CascadeMux
    port map (
            O => \N__27990\,
            I => \N__27987\
        );

    \I__3924\ : InMux
    port map (
            O => \N__27987\,
            I => \N__27984\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__27984\,
            I => \N__27981\
        );

    \I__3922\ : Odrv4
    port map (
            O => \N__27981\,
            I => n3181
        );

    \I__3921\ : InMux
    port map (
            O => \N__27978\,
            I => \N__27975\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__27975\,
            I => \N__27972\
        );

    \I__3919\ : Odrv4
    port map (
            O => \N__27972\,
            I => n3184
        );

    \I__3918\ : InMux
    port map (
            O => \N__27969\,
            I => \N__27964\
        );

    \I__3917\ : InMux
    port map (
            O => \N__27968\,
            I => \N__27961\
        );

    \I__3916\ : InMux
    port map (
            O => \N__27967\,
            I => \N__27958\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__27964\,
            I => \N__27955\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__27961\,
            I => \N__27952\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__27958\,
            I => \N__27949\
        );

    \I__3912\ : Span4Mux_s3_v
    port map (
            O => \N__27955\,
            I => \N__27944\
        );

    \I__3911\ : Span4Mux_v
    port map (
            O => \N__27952\,
            I => \N__27944\
        );

    \I__3910\ : Odrv4
    port map (
            O => \N__27949\,
            I => n3117
        );

    \I__3909\ : Odrv4
    port map (
            O => \N__27944\,
            I => n3117
        );

    \I__3908\ : CascadeMux
    port map (
            O => \N__27939\,
            I => \N__27936\
        );

    \I__3907\ : InMux
    port map (
            O => \N__27936\,
            I => \N__27933\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__27933\,
            I => \N__27930\
        );

    \I__3905\ : Span4Mux_s2_v
    port map (
            O => \N__27930\,
            I => \N__27927\
        );

    \I__3904\ : Odrv4
    port map (
            O => \N__27927\,
            I => n3083
        );

    \I__3903\ : InMux
    port map (
            O => \N__27924\,
            I => \N__27921\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__27921\,
            I => \N__27918\
        );

    \I__3901\ : Odrv4
    port map (
            O => \N__27918\,
            I => n13831
        );

    \I__3900\ : InMux
    port map (
            O => \N__27915\,
            I => \N__27910\
        );

    \I__3899\ : InMux
    port map (
            O => \N__27914\,
            I => \N__27907\
        );

    \I__3898\ : InMux
    port map (
            O => \N__27913\,
            I => \N__27904\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__27910\,
            I => n3114
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__27907\,
            I => n3114
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__27904\,
            I => n3114
        );

    \I__3894\ : CascadeMux
    port map (
            O => \N__27897\,
            I => \n3115_cascade_\
        );

    \I__3893\ : InMux
    port map (
            O => \N__27894\,
            I => \N__27891\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__27891\,
            I => \N__27888\
        );

    \I__3891\ : Span4Mux_v
    port map (
            O => \N__27888\,
            I => \N__27885\
        );

    \I__3890\ : Odrv4
    port map (
            O => \N__27885\,
            I => n14156
        );

    \I__3889\ : InMux
    port map (
            O => \N__27882\,
            I => \N__27878\
        );

    \I__3888\ : InMux
    port map (
            O => \N__27881\,
            I => \N__27874\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__27878\,
            I => \N__27871\
        );

    \I__3886\ : InMux
    port map (
            O => \N__27877\,
            I => \N__27868\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__27874\,
            I => \N__27863\
        );

    \I__3884\ : Span4Mux_s3_h
    port map (
            O => \N__27871\,
            I => \N__27863\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__27868\,
            I => \N__27860\
        );

    \I__3882\ : Span4Mux_v
    port map (
            O => \N__27863\,
            I => \N__27857\
        );

    \I__3881\ : Span12Mux_s2_v
    port map (
            O => \N__27860\,
            I => \N__27854\
        );

    \I__3880\ : Odrv4
    port map (
            O => \N__27857\,
            I => n3113
        );

    \I__3879\ : Odrv12
    port map (
            O => \N__27854\,
            I => n3113
        );

    \I__3878\ : CascadeMux
    port map (
            O => \N__27849\,
            I => \n14162_cascade_\
        );

    \I__3877\ : CascadeMux
    port map (
            O => \N__27846\,
            I => \n14168_cascade_\
        );

    \I__3876\ : InMux
    port map (
            O => \N__27843\,
            I => \N__27839\
        );

    \I__3875\ : InMux
    port map (
            O => \N__27842\,
            I => \N__27836\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__27839\,
            I => n3108
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__27836\,
            I => n3108
        );

    \I__3872\ : InMux
    port map (
            O => \N__27831\,
            I => \N__27828\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__27828\,
            I => n14174
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__27825\,
            I => \N__27822\
        );

    \I__3869\ : InMux
    port map (
            O => \N__27822\,
            I => \N__27819\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__27819\,
            I => \N__27816\
        );

    \I__3867\ : Odrv4
    port map (
            O => \N__27816\,
            I => n3190
        );

    \I__3866\ : InMux
    port map (
            O => \N__27813\,
            I => \N__27810\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__27810\,
            I => \N__27806\
        );

    \I__3864\ : InMux
    port map (
            O => \N__27809\,
            I => \N__27803\
        );

    \I__3863\ : Span4Mux_h
    port map (
            O => \N__27806\,
            I => \N__27799\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__27803\,
            I => \N__27796\
        );

    \I__3861\ : InMux
    port map (
            O => \N__27802\,
            I => \N__27793\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__27799\,
            I => n3121
        );

    \I__3859\ : Odrv4
    port map (
            O => \N__27796\,
            I => n3121
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__27793\,
            I => n3121
        );

    \I__3857\ : InMux
    port map (
            O => \N__27786\,
            I => \N__27783\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__27783\,
            I => \N__27780\
        );

    \I__3855\ : Odrv12
    port map (
            O => \N__27780\,
            I => n3188
        );

    \I__3854\ : InMux
    port map (
            O => \N__27777\,
            I => \N__27774\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__27774\,
            I => \N__27771\
        );

    \I__3852\ : Odrv4
    port map (
            O => \N__27771\,
            I => n3192
        );

    \I__3851\ : CascadeMux
    port map (
            O => \N__27768\,
            I => \N__27765\
        );

    \I__3850\ : InMux
    port map (
            O => \N__27765\,
            I => \N__27761\
        );

    \I__3849\ : CascadeMux
    port map (
            O => \N__27764\,
            I => \N__27758\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__27761\,
            I => \N__27755\
        );

    \I__3847\ : InMux
    port map (
            O => \N__27758\,
            I => \N__27752\
        );

    \I__3846\ : Span4Mux_h
    port map (
            O => \N__27755\,
            I => \N__27748\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__27752\,
            I => \N__27745\
        );

    \I__3844\ : InMux
    port map (
            O => \N__27751\,
            I => \N__27742\
        );

    \I__3843\ : Odrv4
    port map (
            O => \N__27748\,
            I => n3125
        );

    \I__3842\ : Odrv4
    port map (
            O => \N__27745\,
            I => n3125
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__27742\,
            I => n3125
        );

    \I__3840\ : InMux
    port map (
            O => \N__27735\,
            I => \N__27730\
        );

    \I__3839\ : InMux
    port map (
            O => \N__27734\,
            I => \N__27727\
        );

    \I__3838\ : InMux
    port map (
            O => \N__27733\,
            I => \N__27724\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__27730\,
            I => \N__27721\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__27727\,
            I => \N__27718\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__27724\,
            I => \N__27715\
        );

    \I__3834\ : Span4Mux_s2_h
    port map (
            O => \N__27721\,
            I => \N__27712\
        );

    \I__3833\ : Odrv4
    port map (
            O => \N__27718\,
            I => n3127
        );

    \I__3832\ : Odrv4
    port map (
            O => \N__27715\,
            I => n3127
        );

    \I__3831\ : Odrv4
    port map (
            O => \N__27712\,
            I => n3127
        );

    \I__3830\ : CascadeMux
    port map (
            O => \N__27705\,
            I => \N__27702\
        );

    \I__3829\ : InMux
    port map (
            O => \N__27702\,
            I => \N__27699\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__27699\,
            I => \N__27696\
        );

    \I__3827\ : Span4Mux_h
    port map (
            O => \N__27696\,
            I => \N__27693\
        );

    \I__3826\ : Odrv4
    port map (
            O => \N__27693\,
            I => n3194
        );

    \I__3825\ : CascadeMux
    port map (
            O => \N__27690\,
            I => \n3226_cascade_\
        );

    \I__3824\ : InMux
    port map (
            O => \N__27687\,
            I => \N__27684\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__27684\,
            I => \N__27680\
        );

    \I__3822\ : InMux
    port map (
            O => \N__27683\,
            I => \N__27677\
        );

    \I__3821\ : Span4Mux_h
    port map (
            O => \N__27680\,
            I => \N__27671\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__27677\,
            I => \N__27671\
        );

    \I__3819\ : InMux
    port map (
            O => \N__27676\,
            I => \N__27668\
        );

    \I__3818\ : Odrv4
    port map (
            O => \N__27671\,
            I => n3119
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__27668\,
            I => n3119
        );

    \I__3816\ : CascadeMux
    port map (
            O => \N__27663\,
            I => \N__27660\
        );

    \I__3815\ : InMux
    port map (
            O => \N__27660\,
            I => \N__27657\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__27657\,
            I => \N__27654\
        );

    \I__3813\ : Span4Mux_s2_v
    port map (
            O => \N__27654\,
            I => \N__27651\
        );

    \I__3812\ : Odrv4
    port map (
            O => \N__27651\,
            I => n3186
        );

    \I__3811\ : CascadeMux
    port map (
            O => \N__27648\,
            I => \n3218_cascade_\
        );

    \I__3810\ : CascadeMux
    port map (
            O => \N__27645\,
            I => \N__27642\
        );

    \I__3809\ : InMux
    port map (
            O => \N__27642\,
            I => \N__27639\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__27639\,
            I => \N__27636\
        );

    \I__3807\ : Odrv4
    port map (
            O => \N__27636\,
            I => n3180
        );

    \I__3806\ : CascadeMux
    port map (
            O => \N__27633\,
            I => \N__27630\
        );

    \I__3805\ : InMux
    port map (
            O => \N__27630\,
            I => \N__27627\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__27627\,
            I => n3098
        );

    \I__3803\ : CascadeMux
    port map (
            O => \N__27624\,
            I => \n3130_cascade_\
        );

    \I__3802\ : InMux
    port map (
            O => \N__27621\,
            I => \N__27618\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__27618\,
            I => n3101
        );

    \I__3800\ : InMux
    port map (
            O => \N__27615\,
            I => \N__27612\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__27612\,
            I => n3097
        );

    \I__3798\ : InMux
    port map (
            O => \N__27609\,
            I => \N__27606\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__27606\,
            I => n3100
        );

    \I__3796\ : CascadeMux
    port map (
            O => \N__27603\,
            I => \n3132_cascade_\
        );

    \I__3795\ : InMux
    port map (
            O => \N__27600\,
            I => \N__27597\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__27597\,
            I => n11945
        );

    \I__3793\ : InMux
    port map (
            O => \N__27594\,
            I => \N__27591\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__27591\,
            I => n3080
        );

    \I__3791\ : CascadeMux
    port map (
            O => \N__27588\,
            I => \N__27584\
        );

    \I__3790\ : InMux
    port map (
            O => \N__27587\,
            I => \N__27581\
        );

    \I__3789\ : InMux
    port map (
            O => \N__27584\,
            I => \N__27578\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__27581\,
            I => \N__27575\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__27578\,
            I => \N__27571\
        );

    \I__3786\ : Span4Mux_v
    port map (
            O => \N__27575\,
            I => \N__27568\
        );

    \I__3785\ : InMux
    port map (
            O => \N__27574\,
            I => \N__27565\
        );

    \I__3784\ : Odrv4
    port map (
            O => \N__27571\,
            I => n3013
        );

    \I__3783\ : Odrv4
    port map (
            O => \N__27568\,
            I => n3013
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__27565\,
            I => n3013
        );

    \I__3781\ : CascadeMux
    port map (
            O => \N__27558\,
            I => \n23_adj_715_cascade_\
        );

    \I__3780\ : InMux
    port map (
            O => \N__27555\,
            I => \N__27552\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__27552\,
            I => \N__27548\
        );

    \I__3778\ : CascadeMux
    port map (
            O => \N__27551\,
            I => \N__27545\
        );

    \I__3777\ : Span4Mux_h
    port map (
            O => \N__27548\,
            I => \N__27541\
        );

    \I__3776\ : InMux
    port map (
            O => \N__27545\,
            I => \N__27538\
        );

    \I__3775\ : InMux
    port map (
            O => \N__27544\,
            I => \N__27535\
        );

    \I__3774\ : Odrv4
    port map (
            O => \N__27541\,
            I => n3123
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__27538\,
            I => n3123
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__27535\,
            I => n3123
        );

    \I__3771\ : CascadeMux
    port map (
            O => \N__27528\,
            I => \N__27525\
        );

    \I__3770\ : InMux
    port map (
            O => \N__27525\,
            I => \N__27522\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__27522\,
            I => \N__27519\
        );

    \I__3768\ : Span4Mux_h
    port map (
            O => \N__27519\,
            I => \N__27516\
        );

    \I__3767\ : Odrv4
    port map (
            O => \N__27516\,
            I => n2995
        );

    \I__3766\ : CascadeMux
    port map (
            O => \N__27513\,
            I => \N__27510\
        );

    \I__3765\ : InMux
    port map (
            O => \N__27510\,
            I => \N__27507\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__27507\,
            I => \N__27504\
        );

    \I__3763\ : Span4Mux_v
    port map (
            O => \N__27504\,
            I => \N__27501\
        );

    \I__3762\ : Odrv4
    port map (
            O => \N__27501\,
            I => n3000
        );

    \I__3761\ : InMux
    port map (
            O => \N__27498\,
            I => \N__27495\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__27495\,
            I => \N__27491\
        );

    \I__3759\ : InMux
    port map (
            O => \N__27494\,
            I => \N__27488\
        );

    \I__3758\ : Span4Mux_s2_v
    port map (
            O => \N__27491\,
            I => \N__27482\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__27488\,
            I => \N__27482\
        );

    \I__3756\ : InMux
    port map (
            O => \N__27487\,
            I => \N__27479\
        );

    \I__3755\ : Odrv4
    port map (
            O => \N__27482\,
            I => n3015
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__27479\,
            I => n3015
        );

    \I__3753\ : InMux
    port map (
            O => \N__27474\,
            I => \N__27471\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__27471\,
            I => \N__27468\
        );

    \I__3751\ : Span4Mux_v
    port map (
            O => \N__27468\,
            I => \N__27465\
        );

    \I__3750\ : Odrv4
    port map (
            O => \N__27465\,
            I => n14736
        );

    \I__3749\ : InMux
    port map (
            O => \N__27462\,
            I => \N__27458\
        );

    \I__3748\ : CascadeMux
    port map (
            O => \N__27461\,
            I => \N__27454\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__27458\,
            I => \N__27451\
        );

    \I__3746\ : InMux
    port map (
            O => \N__27457\,
            I => \N__27448\
        );

    \I__3745\ : InMux
    port map (
            O => \N__27454\,
            I => \N__27445\
        );

    \I__3744\ : Span4Mux_s3_v
    port map (
            O => \N__27451\,
            I => \N__27440\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__27448\,
            I => \N__27440\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__27445\,
            I => n3014
        );

    \I__3741\ : Odrv4
    port map (
            O => \N__27440\,
            I => n3014
        );

    \I__3740\ : CascadeMux
    port map (
            O => \N__27435\,
            I => \n14742_cascade_\
        );

    \I__3739\ : InMux
    port map (
            O => \N__27432\,
            I => \N__27428\
        );

    \I__3738\ : CascadeMux
    port map (
            O => \N__27431\,
            I => \N__27425\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__27428\,
            I => \N__27422\
        );

    \I__3736\ : InMux
    port map (
            O => \N__27425\,
            I => \N__27419\
        );

    \I__3735\ : Span4Mux_s2_v
    port map (
            O => \N__27422\,
            I => \N__27413\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__27419\,
            I => \N__27413\
        );

    \I__3733\ : InMux
    port map (
            O => \N__27418\,
            I => \N__27410\
        );

    \I__3732\ : Odrv4
    port map (
            O => \N__27413\,
            I => n3011
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__27410\,
            I => n3011
        );

    \I__3730\ : InMux
    port map (
            O => \N__27405\,
            I => \N__27401\
        );

    \I__3729\ : InMux
    port map (
            O => \N__27404\,
            I => \N__27398\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__27401\,
            I => \N__27395\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__27398\,
            I => \N__27391\
        );

    \I__3726\ : Span4Mux_h
    port map (
            O => \N__27395\,
            I => \N__27388\
        );

    \I__3725\ : InMux
    port map (
            O => \N__27394\,
            I => \N__27385\
        );

    \I__3724\ : Span4Mux_h
    port map (
            O => \N__27391\,
            I => \N__27382\
        );

    \I__3723\ : Span4Mux_v
    port map (
            O => \N__27388\,
            I => \N__27377\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__27385\,
            I => \N__27377\
        );

    \I__3721\ : Odrv4
    port map (
            O => \N__27382\,
            I => n3009
        );

    \I__3720\ : Odrv4
    port map (
            O => \N__27377\,
            I => n3009
        );

    \I__3719\ : CascadeMux
    port map (
            O => \N__27372\,
            I => \n14748_cascade_\
        );

    \I__3718\ : CascadeMux
    port map (
            O => \N__27369\,
            I => \N__27366\
        );

    \I__3717\ : InMux
    port map (
            O => \N__27366\,
            I => \N__27362\
        );

    \I__3716\ : InMux
    port map (
            O => \N__27365\,
            I => \N__27359\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__27362\,
            I => \N__27356\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__27359\,
            I => \N__27353\
        );

    \I__3713\ : Odrv4
    port map (
            O => \N__27356\,
            I => n3006
        );

    \I__3712\ : Odrv4
    port map (
            O => \N__27353\,
            I => n3006
        );

    \I__3711\ : InMux
    port map (
            O => \N__27348\,
            I => \N__27342\
        );

    \I__3710\ : InMux
    port map (
            O => \N__27347\,
            I => \N__27342\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__27342\,
            I => \N__27338\
        );

    \I__3708\ : InMux
    port map (
            O => \N__27341\,
            I => \N__27335\
        );

    \I__3707\ : Sp12to4
    port map (
            O => \N__27338\,
            I => \N__27330\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__27335\,
            I => \N__27330\
        );

    \I__3705\ : Odrv12
    port map (
            O => \N__27330\,
            I => n3008
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__27327\,
            I => \n14754_cascade_\
        );

    \I__3703\ : InMux
    port map (
            O => \N__27324\,
            I => \N__27318\
        );

    \I__3702\ : InMux
    port map (
            O => \N__27323\,
            I => \N__27318\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__27318\,
            I => \N__27315\
        );

    \I__3700\ : Span4Mux_s2_v
    port map (
            O => \N__27315\,
            I => \N__27312\
        );

    \I__3699\ : IoSpan4Mux
    port map (
            O => \N__27312\,
            I => \N__27308\
        );

    \I__3698\ : InMux
    port map (
            O => \N__27311\,
            I => \N__27305\
        );

    \I__3697\ : IoSpan4Mux
    port map (
            O => \N__27308\,
            I => \N__27302\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__27305\,
            I => \N__27299\
        );

    \I__3695\ : Span4Mux_s0_h
    port map (
            O => \N__27302\,
            I => \N__27294\
        );

    \I__3694\ : Span4Mux_v
    port map (
            O => \N__27299\,
            I => \N__27294\
        );

    \I__3693\ : Odrv4
    port map (
            O => \N__27294\,
            I => n3007
        );

    \I__3692\ : InMux
    port map (
            O => \N__27291\,
            I => \N__27288\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__27288\,
            I => n3099
        );

    \I__3690\ : CascadeMux
    port map (
            O => \N__27285\,
            I => \n3039_cascade_\
        );

    \I__3689\ : InMux
    port map (
            O => \N__27282\,
            I => \N__27279\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__27279\,
            I => \N__27274\
        );

    \I__3687\ : InMux
    port map (
            O => \N__27278\,
            I => \N__27271\
        );

    \I__3686\ : InMux
    port map (
            O => \N__27277\,
            I => \N__27268\
        );

    \I__3685\ : Span4Mux_h
    port map (
            O => \N__27274\,
            I => \N__27263\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__27271\,
            I => \N__27263\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__27268\,
            I => \N__27260\
        );

    \I__3682\ : Span4Mux_v
    port map (
            O => \N__27263\,
            I => \N__27257\
        );

    \I__3681\ : Odrv4
    port map (
            O => \N__27260\,
            I => n3018
        );

    \I__3680\ : Odrv4
    port map (
            O => \N__27257\,
            I => n3018
        );

    \I__3679\ : CascadeMux
    port map (
            O => \N__27252\,
            I => \N__27249\
        );

    \I__3678\ : InMux
    port map (
            O => \N__27249\,
            I => \N__27246\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__27246\,
            I => n3085
        );

    \I__3676\ : InMux
    port map (
            O => \N__27243\,
            I => \N__27240\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__27240\,
            I => \N__27236\
        );

    \I__3674\ : InMux
    port map (
            O => \N__27239\,
            I => \N__27232\
        );

    \I__3673\ : Span4Mux_h
    port map (
            O => \N__27236\,
            I => \N__27229\
        );

    \I__3672\ : InMux
    port map (
            O => \N__27235\,
            I => \N__27226\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__27232\,
            I => \N__27223\
        );

    \I__3670\ : Odrv4
    port map (
            O => \N__27229\,
            I => n2817
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__27226\,
            I => n2817
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__27223\,
            I => n2817
        );

    \I__3667\ : InMux
    port map (
            O => \N__27216\,
            I => \N__27213\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__27213\,
            I => \N__27210\
        );

    \I__3665\ : Span4Mux_h
    port map (
            O => \N__27210\,
            I => \N__27207\
        );

    \I__3664\ : Odrv4
    port map (
            O => \N__27207\,
            I => n2884
        );

    \I__3663\ : InMux
    port map (
            O => \N__27204\,
            I => \N__27201\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__27201\,
            I => \N__27197\
        );

    \I__3661\ : InMux
    port map (
            O => \N__27200\,
            I => \N__27193\
        );

    \I__3660\ : Span4Mux_s3_h
    port map (
            O => \N__27197\,
            I => \N__27190\
        );

    \I__3659\ : InMux
    port map (
            O => \N__27196\,
            I => \N__27187\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__27193\,
            I => n2916
        );

    \I__3657\ : Odrv4
    port map (
            O => \N__27190\,
            I => n2916
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__27187\,
            I => n2916
        );

    \I__3655\ : CascadeMux
    port map (
            O => \N__27180\,
            I => \N__27177\
        );

    \I__3654\ : InMux
    port map (
            O => \N__27177\,
            I => \N__27174\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__27174\,
            I => \N__27171\
        );

    \I__3652\ : Odrv4
    port map (
            O => \N__27171\,
            I => n2981
        );

    \I__3651\ : CascadeMux
    port map (
            O => \N__27168\,
            I => \N__27163\
        );

    \I__3650\ : CascadeMux
    port map (
            O => \N__27167\,
            I => \N__27160\
        );

    \I__3649\ : CascadeMux
    port map (
            O => \N__27166\,
            I => \N__27157\
        );

    \I__3648\ : InMux
    port map (
            O => \N__27163\,
            I => \N__27154\
        );

    \I__3647\ : InMux
    port map (
            O => \N__27160\,
            I => \N__27151\
        );

    \I__3646\ : InMux
    port map (
            O => \N__27157\,
            I => \N__27148\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__27154\,
            I => \N__27145\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__27151\,
            I => \N__27142\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__27148\,
            I => \N__27139\
        );

    \I__3642\ : Span4Mux_v
    port map (
            O => \N__27145\,
            I => \N__27134\
        );

    \I__3641\ : Span4Mux_s3_h
    port map (
            O => \N__27142\,
            I => \N__27134\
        );

    \I__3640\ : Odrv12
    port map (
            O => \N__27139\,
            I => n2929
        );

    \I__3639\ : Odrv4
    port map (
            O => \N__27134\,
            I => n2929
        );

    \I__3638\ : InMux
    port map (
            O => \N__27129\,
            I => \N__27126\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__27126\,
            I => n14222
        );

    \I__3636\ : InMux
    port map (
            O => \N__27123\,
            I => \N__27120\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__27120\,
            I => \N__27115\
        );

    \I__3634\ : InMux
    port map (
            O => \N__27119\,
            I => \N__27112\
        );

    \I__3633\ : InMux
    port map (
            O => \N__27118\,
            I => \N__27109\
        );

    \I__3632\ : Span4Mux_v
    port map (
            O => \N__27115\,
            I => \N__27106\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__27112\,
            I => \N__27103\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__27109\,
            I => n2915
        );

    \I__3629\ : Odrv4
    port map (
            O => \N__27106\,
            I => n2915
        );

    \I__3628\ : Odrv4
    port map (
            O => \N__27103\,
            I => n2915
        );

    \I__3627\ : CascadeMux
    port map (
            O => \N__27096\,
            I => \n14224_cascade_\
        );

    \I__3626\ : InMux
    port map (
            O => \N__27093\,
            I => \N__27088\
        );

    \I__3625\ : InMux
    port map (
            O => \N__27092\,
            I => \N__27083\
        );

    \I__3624\ : InMux
    port map (
            O => \N__27091\,
            I => \N__27083\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__27088\,
            I => \N__27078\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__27083\,
            I => \N__27078\
        );

    \I__3621\ : Span4Mux_h
    port map (
            O => \N__27078\,
            I => \N__27075\
        );

    \I__3620\ : Odrv4
    port map (
            O => \N__27075\,
            I => n2914
        );

    \I__3619\ : InMux
    port map (
            O => \N__27072\,
            I => \N__27068\
        );

    \I__3618\ : InMux
    port map (
            O => \N__27071\,
            I => \N__27065\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__27068\,
            I => \N__27059\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__27065\,
            I => \N__27059\
        );

    \I__3615\ : InMux
    port map (
            O => \N__27064\,
            I => \N__27056\
        );

    \I__3614\ : Span12Mux_s3_h
    port map (
            O => \N__27059\,
            I => \N__27053\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__27056\,
            I => \N__27050\
        );

    \I__3612\ : Odrv12
    port map (
            O => \N__27053\,
            I => n2910
        );

    \I__3611\ : Odrv4
    port map (
            O => \N__27050\,
            I => n2910
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__27045\,
            I => \n14230_cascade_\
        );

    \I__3609\ : InMux
    port map (
            O => \N__27042\,
            I => \N__27038\
        );

    \I__3608\ : InMux
    port map (
            O => \N__27041\,
            I => \N__27035\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__27038\,
            I => n2912
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__27035\,
            I => n2912
        );

    \I__3605\ : CascadeMux
    port map (
            O => \N__27030\,
            I => \N__27027\
        );

    \I__3604\ : InMux
    port map (
            O => \N__27027\,
            I => \N__27023\
        );

    \I__3603\ : InMux
    port map (
            O => \N__27026\,
            I => \N__27020\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__27023\,
            I => \N__27017\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__27020\,
            I => \N__27014\
        );

    \I__3600\ : Span4Mux_h
    port map (
            O => \N__27017\,
            I => \N__27011\
        );

    \I__3599\ : Span4Mux_h
    port map (
            O => \N__27014\,
            I => \N__27008\
        );

    \I__3598\ : Odrv4
    port map (
            O => \N__27011\,
            I => n2908
        );

    \I__3597\ : Odrv4
    port map (
            O => \N__27008\,
            I => n2908
        );

    \I__3596\ : InMux
    port map (
            O => \N__27003\,
            I => \N__26999\
        );

    \I__3595\ : InMux
    port map (
            O => \N__27002\,
            I => \N__26996\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__26999\,
            I => \N__26993\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__26996\,
            I => \N__26990\
        );

    \I__3592\ : Span4Mux_v
    port map (
            O => \N__26993\,
            I => \N__26987\
        );

    \I__3591\ : Odrv4
    port map (
            O => \N__26990\,
            I => n2907
        );

    \I__3590\ : Odrv4
    port map (
            O => \N__26987\,
            I => n2907
        );

    \I__3589\ : CascadeMux
    port map (
            O => \N__26982\,
            I => \n14236_cascade_\
        );

    \I__3588\ : CascadeMux
    port map (
            O => \N__26979\,
            I => \N__26976\
        );

    \I__3587\ : InMux
    port map (
            O => \N__26976\,
            I => \N__26973\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__26973\,
            I => \N__26968\
        );

    \I__3585\ : InMux
    port map (
            O => \N__26972\,
            I => \N__26965\
        );

    \I__3584\ : InMux
    port map (
            O => \N__26971\,
            I => \N__26962\
        );

    \I__3583\ : Span4Mux_s3_h
    port map (
            O => \N__26968\,
            I => \N__26957\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__26965\,
            I => \N__26957\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__26962\,
            I => n2909
        );

    \I__3580\ : Odrv4
    port map (
            O => \N__26957\,
            I => n2909
        );

    \I__3579\ : CascadeMux
    port map (
            O => \N__26952\,
            I => \n2940_cascade_\
        );

    \I__3578\ : InMux
    port map (
            O => \N__26949\,
            I => \N__26946\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__26946\,
            I => \N__26943\
        );

    \I__3576\ : Span4Mux_h
    port map (
            O => \N__26943\,
            I => \N__26940\
        );

    \I__3575\ : Odrv4
    port map (
            O => \N__26940\,
            I => n2997
        );

    \I__3574\ : InMux
    port map (
            O => \N__26937\,
            I => \N__26932\
        );

    \I__3573\ : InMux
    port map (
            O => \N__26936\,
            I => \N__26927\
        );

    \I__3572\ : InMux
    port map (
            O => \N__26935\,
            I => \N__26927\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__26932\,
            I => n2911
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__26927\,
            I => n2911
        );

    \I__3569\ : InMux
    port map (
            O => \N__26922\,
            I => \N__26919\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__26919\,
            I => \N__26916\
        );

    \I__3567\ : Odrv4
    port map (
            O => \N__26916\,
            I => n2978
        );

    \I__3566\ : InMux
    port map (
            O => \N__26913\,
            I => \N__26910\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__26910\,
            I => \N__26907\
        );

    \I__3564\ : Span4Mux_v
    port map (
            O => \N__26907\,
            I => \N__26904\
        );

    \I__3563\ : Odrv4
    port map (
            O => \N__26904\,
            I => n3081
        );

    \I__3562\ : InMux
    port map (
            O => \N__26901\,
            I => \N__26898\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__26898\,
            I => \N__26895\
        );

    \I__3560\ : Span4Mux_s2_h
    port map (
            O => \N__26895\,
            I => \N__26890\
        );

    \I__3559\ : InMux
    port map (
            O => \N__26894\,
            I => \N__26885\
        );

    \I__3558\ : InMux
    port map (
            O => \N__26893\,
            I => \N__26885\
        );

    \I__3557\ : Odrv4
    port map (
            O => \N__26890\,
            I => n2810
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__26885\,
            I => n2810
        );

    \I__3555\ : InMux
    port map (
            O => \N__26880\,
            I => \N__26877\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__26877\,
            I => \N__26874\
        );

    \I__3553\ : Odrv12
    port map (
            O => \N__26874\,
            I => n2877
        );

    \I__3552\ : CascadeMux
    port map (
            O => \N__26871\,
            I => \N__26868\
        );

    \I__3551\ : InMux
    port map (
            O => \N__26868\,
            I => \N__26865\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__26865\,
            I => \N__26862\
        );

    \I__3549\ : Span4Mux_v
    port map (
            O => \N__26862\,
            I => \N__26859\
        );

    \I__3548\ : Odrv4
    port map (
            O => \N__26859\,
            I => n2976
        );

    \I__3547\ : InMux
    port map (
            O => \N__26856\,
            I => \N__26853\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__26853\,
            I => \N__26850\
        );

    \I__3545\ : Span4Mux_h
    port map (
            O => \N__26850\,
            I => \N__26847\
        );

    \I__3544\ : Odrv4
    port map (
            O => \N__26847\,
            I => n2886
        );

    \I__3543\ : InMux
    port map (
            O => \N__26844\,
            I => \N__26840\
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__26843\,
            I => \N__26837\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__26840\,
            I => \N__26834\
        );

    \I__3540\ : InMux
    port map (
            O => \N__26837\,
            I => \N__26830\
        );

    \I__3539\ : Span4Mux_s2_h
    port map (
            O => \N__26834\,
            I => \N__26827\
        );

    \I__3538\ : InMux
    port map (
            O => \N__26833\,
            I => \N__26824\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__26830\,
            I => n2819
        );

    \I__3536\ : Odrv4
    port map (
            O => \N__26827\,
            I => n2819
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__26824\,
            I => n2819
        );

    \I__3534\ : InMux
    port map (
            O => \N__26817\,
            I => \N__26814\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__26814\,
            I => \N__26810\
        );

    \I__3532\ : InMux
    port map (
            O => \N__26813\,
            I => \N__26807\
        );

    \I__3531\ : IoSpan4Mux
    port map (
            O => \N__26810\,
            I => \N__26802\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__26807\,
            I => \N__26802\
        );

    \I__3529\ : Span4Mux_s3_h
    port map (
            O => \N__26802\,
            I => \N__26799\
        );

    \I__3528\ : Odrv4
    port map (
            O => \N__26799\,
            I => n2918
        );

    \I__3527\ : InMux
    port map (
            O => \N__26796\,
            I => \N__26792\
        );

    \I__3526\ : InMux
    port map (
            O => \N__26795\,
            I => \N__26789\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__26792\,
            I => \N__26786\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__26789\,
            I => n2927
        );

    \I__3523\ : Odrv4
    port map (
            O => \N__26786\,
            I => n2927
        );

    \I__3522\ : InMux
    port map (
            O => \N__26781\,
            I => \N__26778\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__26778\,
            I => \N__26775\
        );

    \I__3520\ : Span4Mux_s2_h
    port map (
            O => \N__26775\,
            I => \N__26770\
        );

    \I__3519\ : InMux
    port map (
            O => \N__26774\,
            I => \N__26767\
        );

    \I__3518\ : InMux
    port map (
            O => \N__26773\,
            I => \N__26764\
        );

    \I__3517\ : Odrv4
    port map (
            O => \N__26770\,
            I => n2926
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__26767\,
            I => n2926
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__26764\,
            I => n2926
        );

    \I__3514\ : CascadeMux
    port map (
            O => \N__26757\,
            I => \n2918_cascade_\
        );

    \I__3513\ : InMux
    port map (
            O => \N__26754\,
            I => \N__26751\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__26751\,
            I => \N__26747\
        );

    \I__3511\ : CascadeMux
    port map (
            O => \N__26750\,
            I => \N__26744\
        );

    \I__3510\ : Span4Mux_v
    port map (
            O => \N__26747\,
            I => \N__26741\
        );

    \I__3509\ : InMux
    port map (
            O => \N__26744\,
            I => \N__26737\
        );

    \I__3508\ : IoSpan4Mux
    port map (
            O => \N__26741\,
            I => \N__26734\
        );

    \I__3507\ : InMux
    port map (
            O => \N__26740\,
            I => \N__26731\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__26737\,
            I => \N__26728\
        );

    \I__3505\ : Span4Mux_s1_h
    port map (
            O => \N__26734\,
            I => \N__26723\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__26731\,
            I => \N__26723\
        );

    \I__3503\ : Span4Mux_v
    port map (
            O => \N__26728\,
            I => \N__26720\
        );

    \I__3502\ : Odrv4
    port map (
            O => \N__26723\,
            I => n2825
        );

    \I__3501\ : Odrv4
    port map (
            O => \N__26720\,
            I => n2825
        );

    \I__3500\ : CascadeMux
    port map (
            O => \N__26715\,
            I => \N__26712\
        );

    \I__3499\ : InMux
    port map (
            O => \N__26712\,
            I => \N__26709\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__26709\,
            I => \N__26706\
        );

    \I__3497\ : Span4Mux_v
    port map (
            O => \N__26706\,
            I => \N__26703\
        );

    \I__3496\ : Odrv4
    port map (
            O => \N__26703\,
            I => n2892
        );

    \I__3495\ : InMux
    port map (
            O => \N__26700\,
            I => \N__26695\
        );

    \I__3494\ : InMux
    port map (
            O => \N__26699\,
            I => \N__26692\
        );

    \I__3493\ : InMux
    port map (
            O => \N__26698\,
            I => \N__26689\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__26695\,
            I => n2921
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__26692\,
            I => n2921
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__26689\,
            I => n2921
        );

    \I__3489\ : InMux
    port map (
            O => \N__26682\,
            I => \N__26679\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__26679\,
            I => \N__26676\
        );

    \I__3487\ : Span4Mux_s2_h
    port map (
            O => \N__26676\,
            I => \N__26671\
        );

    \I__3486\ : InMux
    port map (
            O => \N__26675\,
            I => \N__26668\
        );

    \I__3485\ : InMux
    port map (
            O => \N__26674\,
            I => \N__26665\
        );

    \I__3484\ : Odrv4
    port map (
            O => \N__26671\,
            I => n2922
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__26668\,
            I => n2922
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__26665\,
            I => n2922
        );

    \I__3481\ : CascadeMux
    port map (
            O => \N__26658\,
            I => \n2924_cascade_\
        );

    \I__3480\ : InMux
    port map (
            O => \N__26655\,
            I => \N__26650\
        );

    \I__3479\ : InMux
    port map (
            O => \N__26654\,
            I => \N__26647\
        );

    \I__3478\ : InMux
    port map (
            O => \N__26653\,
            I => \N__26644\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__26650\,
            I => n2919
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__26647\,
            I => n2919
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__26644\,
            I => n2919
        );

    \I__3474\ : CascadeMux
    port map (
            O => \N__26637\,
            I => \n14212_cascade_\
        );

    \I__3473\ : InMux
    port map (
            O => \N__26634\,
            I => \N__26631\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__26631\,
            I => n14216
        );

    \I__3471\ : CascadeMux
    port map (
            O => \N__26628\,
            I => \N__26625\
        );

    \I__3470\ : InMux
    port map (
            O => \N__26625\,
            I => \N__26622\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__26622\,
            I => \N__26619\
        );

    \I__3468\ : Span4Mux_v
    port map (
            O => \N__26619\,
            I => \N__26615\
        );

    \I__3467\ : InMux
    port map (
            O => \N__26618\,
            I => \N__26611\
        );

    \I__3466\ : Span4Mux_s2_h
    port map (
            O => \N__26615\,
            I => \N__26608\
        );

    \I__3465\ : InMux
    port map (
            O => \N__26614\,
            I => \N__26605\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__26611\,
            I => n2733
        );

    \I__3463\ : Odrv4
    port map (
            O => \N__26608\,
            I => n2733
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__26605\,
            I => n2733
        );

    \I__3461\ : CascadeMux
    port map (
            O => \N__26598\,
            I => \N__26595\
        );

    \I__3460\ : InMux
    port map (
            O => \N__26595\,
            I => \N__26592\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__26592\,
            I => \N__26589\
        );

    \I__3458\ : Span4Mux_v
    port map (
            O => \N__26589\,
            I => \N__26586\
        );

    \I__3457\ : Span4Mux_v
    port map (
            O => \N__26586\,
            I => \N__26583\
        );

    \I__3456\ : Odrv4
    port map (
            O => \N__26583\,
            I => n2800
        );

    \I__3455\ : CascadeMux
    port map (
            O => \N__26580\,
            I => \n2832_cascade_\
        );

    \I__3454\ : CascadeMux
    port map (
            O => \N__26577\,
            I => \N__26574\
        );

    \I__3453\ : InMux
    port map (
            O => \N__26574\,
            I => \N__26569\
        );

    \I__3452\ : InMux
    port map (
            O => \N__26573\,
            I => \N__26566\
        );

    \I__3451\ : InMux
    port map (
            O => \N__26572\,
            I => \N__26563\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__26569\,
            I => \N__26560\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__26566\,
            I => \N__26557\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__26563\,
            I => \N__26552\
        );

    \I__3447\ : Span4Mux_s1_h
    port map (
            O => \N__26560\,
            I => \N__26552\
        );

    \I__3446\ : Span4Mux_v
    port map (
            O => \N__26557\,
            I => \N__26549\
        );

    \I__3445\ : Odrv4
    port map (
            O => \N__26552\,
            I => n2833
        );

    \I__3444\ : Odrv4
    port map (
            O => \N__26549\,
            I => n2833
        );

    \I__3443\ : CascadeMux
    port map (
            O => \N__26544\,
            I => \N__26541\
        );

    \I__3442\ : InMux
    port map (
            O => \N__26541\,
            I => \N__26537\
        );

    \I__3441\ : CascadeMux
    port map (
            O => \N__26540\,
            I => \N__26534\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__26537\,
            I => \N__26530\
        );

    \I__3439\ : InMux
    port map (
            O => \N__26534\,
            I => \N__26525\
        );

    \I__3438\ : InMux
    port map (
            O => \N__26533\,
            I => \N__26525\
        );

    \I__3437\ : Span4Mux_s2_h
    port map (
            O => \N__26530\,
            I => \N__26522\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__26525\,
            I => n2830
        );

    \I__3435\ : Odrv4
    port map (
            O => \N__26522\,
            I => n2830
        );

    \I__3434\ : CascadeMux
    port map (
            O => \N__26517\,
            I => \n11953_cascade_\
        );

    \I__3433\ : InMux
    port map (
            O => \N__26514\,
            I => \N__26511\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__26511\,
            I => n13857
        );

    \I__3431\ : CascadeMux
    port map (
            O => \N__26508\,
            I => \N__26505\
        );

    \I__3430\ : InMux
    port map (
            O => \N__26505\,
            I => \N__26501\
        );

    \I__3429\ : CascadeMux
    port map (
            O => \N__26504\,
            I => \N__26497\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__26501\,
            I => \N__26494\
        );

    \I__3427\ : InMux
    port map (
            O => \N__26500\,
            I => \N__26491\
        );

    \I__3426\ : InMux
    port map (
            O => \N__26497\,
            I => \N__26488\
        );

    \I__3425\ : Span4Mux_h
    port map (
            O => \N__26494\,
            I => \N__26485\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__26491\,
            I => n2815
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__26488\,
            I => n2815
        );

    \I__3422\ : Odrv4
    port map (
            O => \N__26485\,
            I => n2815
        );

    \I__3421\ : InMux
    port map (
            O => \N__26478\,
            I => \N__26475\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__26475\,
            I => n14702
        );

    \I__3419\ : InMux
    port map (
            O => \N__26472\,
            I => \N__26468\
        );

    \I__3418\ : InMux
    port map (
            O => \N__26471\,
            I => \N__26465\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__26468\,
            I => \N__26461\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__26465\,
            I => \N__26458\
        );

    \I__3415\ : InMux
    port map (
            O => \N__26464\,
            I => \N__26455\
        );

    \I__3414\ : Odrv4
    port map (
            O => \N__26461\,
            I => n2812
        );

    \I__3413\ : Odrv4
    port map (
            O => \N__26458\,
            I => n2812
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__26455\,
            I => n2812
        );

    \I__3411\ : CascadeMux
    port map (
            O => \N__26448\,
            I => \N__26444\
        );

    \I__3410\ : InMux
    port map (
            O => \N__26447\,
            I => \N__26441\
        );

    \I__3409\ : InMux
    port map (
            O => \N__26444\,
            I => \N__26438\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__26441\,
            I => \N__26435\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__26438\,
            I => \N__26429\
        );

    \I__3406\ : Span4Mux_s2_h
    port map (
            O => \N__26435\,
            I => \N__26429\
        );

    \I__3405\ : InMux
    port map (
            O => \N__26434\,
            I => \N__26426\
        );

    \I__3404\ : Odrv4
    port map (
            O => \N__26429\,
            I => n2813
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__26426\,
            I => n2813
        );

    \I__3402\ : CascadeMux
    port map (
            O => \N__26421\,
            I => \n14708_cascade_\
        );

    \I__3401\ : InMux
    port map (
            O => \N__26418\,
            I => \N__26415\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__26415\,
            I => \N__26411\
        );

    \I__3399\ : InMux
    port map (
            O => \N__26414\,
            I => \N__26408\
        );

    \I__3398\ : Odrv4
    port map (
            O => \N__26411\,
            I => n2811
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__26408\,
            I => n2811
        );

    \I__3396\ : InMux
    port map (
            O => \N__26403\,
            I => \N__26399\
        );

    \I__3395\ : InMux
    port map (
            O => \N__26402\,
            I => \N__26396\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__26399\,
            I => \N__26392\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__26396\,
            I => \N__26389\
        );

    \I__3392\ : InMux
    port map (
            O => \N__26395\,
            I => \N__26386\
        );

    \I__3391\ : Span4Mux_v
    port map (
            O => \N__26392\,
            I => \N__26383\
        );

    \I__3390\ : Span4Mux_s2_h
    port map (
            O => \N__26389\,
            I => \N__26380\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__26386\,
            I => \N__26377\
        );

    \I__3388\ : Odrv4
    port map (
            O => \N__26383\,
            I => n2809
        );

    \I__3387\ : Odrv4
    port map (
            O => \N__26380\,
            I => n2809
        );

    \I__3386\ : Odrv4
    port map (
            O => \N__26377\,
            I => n2809
        );

    \I__3385\ : CascadeMux
    port map (
            O => \N__26370\,
            I => \n14714_cascade_\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__26367\,
            I => \N__26363\
        );

    \I__3383\ : InMux
    port map (
            O => \N__26366\,
            I => \N__26360\
        );

    \I__3382\ : InMux
    port map (
            O => \N__26363\,
            I => \N__26357\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__26360\,
            I => \N__26354\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__26357\,
            I => \N__26351\
        );

    \I__3379\ : Span4Mux_v
    port map (
            O => \N__26354\,
            I => \N__26348\
        );

    \I__3378\ : Span4Mux_v
    port map (
            O => \N__26351\,
            I => \N__26345\
        );

    \I__3377\ : Span4Mux_v
    port map (
            O => \N__26348\,
            I => \N__26342\
        );

    \I__3376\ : Odrv4
    port map (
            O => \N__26345\,
            I => n2808
        );

    \I__3375\ : Odrv4
    port map (
            O => \N__26342\,
            I => n2808
        );

    \I__3374\ : InMux
    port map (
            O => \N__26337\,
            I => \N__26334\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__26334\,
            I => \N__26329\
        );

    \I__3372\ : InMux
    port map (
            O => \N__26333\,
            I => \N__26324\
        );

    \I__3371\ : InMux
    port map (
            O => \N__26332\,
            I => \N__26324\
        );

    \I__3370\ : Odrv4
    port map (
            O => \N__26329\,
            I => n2816
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__26324\,
            I => n2816
        );

    \I__3368\ : CascadeMux
    port map (
            O => \N__26319\,
            I => \n2841_cascade_\
        );

    \I__3367\ : InMux
    port map (
            O => \N__26316\,
            I => \N__26313\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__26313\,
            I => \N__26310\
        );

    \I__3365\ : Span4Mux_h
    port map (
            O => \N__26310\,
            I => \N__26307\
        );

    \I__3364\ : Odrv4
    port map (
            O => \N__26307\,
            I => n2883
        );

    \I__3363\ : InMux
    port map (
            O => \N__26304\,
            I => \N__26301\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__26301\,
            I => \N__26298\
        );

    \I__3361\ : Span4Mux_h
    port map (
            O => \N__26298\,
            I => \N__26295\
        );

    \I__3360\ : Odrv4
    port map (
            O => \N__26295\,
            I => n2885
        );

    \I__3359\ : InMux
    port map (
            O => \N__26292\,
            I => \N__26288\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__26291\,
            I => \N__26285\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__26288\,
            I => \N__26282\
        );

    \I__3356\ : InMux
    port map (
            O => \N__26285\,
            I => \N__26278\
        );

    \I__3355\ : Span4Mux_s1_h
    port map (
            O => \N__26282\,
            I => \N__26275\
        );

    \I__3354\ : InMux
    port map (
            O => \N__26281\,
            I => \N__26272\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__26278\,
            I => n2818
        );

    \I__3352\ : Odrv4
    port map (
            O => \N__26275\,
            I => n2818
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__26272\,
            I => n2818
        );

    \I__3350\ : InMux
    port map (
            O => \N__26265\,
            I => \N__26262\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__26262\,
            I => \N__26258\
        );

    \I__3348\ : InMux
    port map (
            O => \N__26261\,
            I => \N__26255\
        );

    \I__3347\ : Span12Mux_s3_h
    port map (
            O => \N__26258\,
            I => \N__26252\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__26255\,
            I => n2633
        );

    \I__3345\ : Odrv12
    port map (
            O => \N__26252\,
            I => n2633
        );

    \I__3344\ : CascadeMux
    port map (
            O => \N__26247\,
            I => \n2633_cascade_\
        );

    \I__3343\ : CascadeMux
    port map (
            O => \N__26244\,
            I => \N__26241\
        );

    \I__3342\ : InMux
    port map (
            O => \N__26241\,
            I => \N__26238\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__26238\,
            I => n12059
        );

    \I__3340\ : InMux
    port map (
            O => \N__26235\,
            I => \N__26232\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__26232\,
            I => \N__26227\
        );

    \I__3338\ : CascadeMux
    port map (
            O => \N__26231\,
            I => \N__26224\
        );

    \I__3337\ : InMux
    port map (
            O => \N__26230\,
            I => \N__26221\
        );

    \I__3336\ : Span12Mux_s3_h
    port map (
            O => \N__26227\,
            I => \N__26218\
        );

    \I__3335\ : InMux
    port map (
            O => \N__26224\,
            I => \N__26215\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__26221\,
            I => n2618
        );

    \I__3333\ : Odrv12
    port map (
            O => \N__26218\,
            I => n2618
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__26215\,
            I => n2618
        );

    \I__3331\ : InMux
    port map (
            O => \N__26208\,
            I => \N__26204\
        );

    \I__3330\ : InMux
    port map (
            O => \N__26207\,
            I => \N__26201\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__26204\,
            I => \N__26198\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__26201\,
            I => \N__26195\
        );

    \I__3327\ : Span4Mux_s3_h
    port map (
            O => \N__26198\,
            I => \N__26192\
        );

    \I__3326\ : Span4Mux_s3_h
    port map (
            O => \N__26195\,
            I => \N__26188\
        );

    \I__3325\ : Span4Mux_v
    port map (
            O => \N__26192\,
            I => \N__26185\
        );

    \I__3324\ : InMux
    port map (
            O => \N__26191\,
            I => \N__26182\
        );

    \I__3323\ : Odrv4
    port map (
            O => \N__26188\,
            I => n2614
        );

    \I__3322\ : Odrv4
    port map (
            O => \N__26185\,
            I => n2614
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__26182\,
            I => n2614
        );

    \I__3320\ : InMux
    port map (
            O => \N__26175\,
            I => \N__26172\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__26172\,
            I => \N__26169\
        );

    \I__3318\ : Span4Mux_s3_h
    port map (
            O => \N__26169\,
            I => \N__26165\
        );

    \I__3317\ : InMux
    port map (
            O => \N__26168\,
            I => \N__26161\
        );

    \I__3316\ : Sp12to4
    port map (
            O => \N__26165\,
            I => \N__26158\
        );

    \I__3315\ : InMux
    port map (
            O => \N__26164\,
            I => \N__26155\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__26161\,
            I => n2613
        );

    \I__3313\ : Odrv12
    port map (
            O => \N__26158\,
            I => n2613
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__26155\,
            I => n2613
        );

    \I__3311\ : CascadeMux
    port map (
            O => \N__26148\,
            I => \N__26145\
        );

    \I__3310\ : InMux
    port map (
            O => \N__26145\,
            I => \N__26142\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__26142\,
            I => \N__26139\
        );

    \I__3308\ : Span4Mux_s3_h
    port map (
            O => \N__26139\,
            I => \N__26136\
        );

    \I__3307\ : Span4Mux_v
    port map (
            O => \N__26136\,
            I => \N__26131\
        );

    \I__3306\ : InMux
    port map (
            O => \N__26135\,
            I => \N__26126\
        );

    \I__3305\ : InMux
    port map (
            O => \N__26134\,
            I => \N__26126\
        );

    \I__3304\ : Span4Mux_v
    port map (
            O => \N__26131\,
            I => \N__26123\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__26126\,
            I => n2619
        );

    \I__3302\ : Odrv4
    port map (
            O => \N__26123\,
            I => n2619
        );

    \I__3301\ : InMux
    port map (
            O => \N__26118\,
            I => \N__26115\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__26115\,
            I => \N__26112\
        );

    \I__3299\ : Span4Mux_h
    port map (
            O => \N__26112\,
            I => \N__26109\
        );

    \I__3298\ : Odrv4
    port map (
            O => \N__26109\,
            I => n2897
        );

    \I__3297\ : InMux
    port map (
            O => \N__26106\,
            I => \N__26103\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__26103\,
            I => \N__26099\
        );

    \I__3295\ : InMux
    port map (
            O => \N__26102\,
            I => \N__26095\
        );

    \I__3294\ : Span12Mux_s2_h
    port map (
            O => \N__26099\,
            I => \N__26092\
        );

    \I__3293\ : InMux
    port map (
            O => \N__26098\,
            I => \N__26089\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__26095\,
            I => n2712
        );

    \I__3291\ : Odrv12
    port map (
            O => \N__26092\,
            I => n2712
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__26089\,
            I => n2712
        );

    \I__3289\ : CascadeMux
    port map (
            O => \N__26082\,
            I => \N__26079\
        );

    \I__3288\ : InMux
    port map (
            O => \N__26079\,
            I => \N__26076\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__26076\,
            I => \N__26073\
        );

    \I__3286\ : Span12Mux_v
    port map (
            O => \N__26073\,
            I => \N__26070\
        );

    \I__3285\ : Odrv12
    port map (
            O => \N__26070\,
            I => n2779
        );

    \I__3284\ : InMux
    port map (
            O => \N__26067\,
            I => \N__26064\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__26064\,
            I => \N__26061\
        );

    \I__3282\ : Odrv12
    port map (
            O => \N__26061\,
            I => n2878
        );

    \I__3281\ : CascadeMux
    port map (
            O => \N__26058\,
            I => \n2811_cascade_\
        );

    \I__3280\ : CascadeMux
    port map (
            O => \N__26055\,
            I => \n2524_cascade_\
        );

    \I__3279\ : CascadeMux
    port map (
            O => \N__26052\,
            I => \n14574_cascade_\
        );

    \I__3278\ : CascadeMux
    port map (
            O => \N__26049\,
            I => \n2523_cascade_\
        );

    \I__3277\ : InMux
    port map (
            O => \N__26046\,
            I => \N__26043\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__26043\,
            I => n14576
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__26040\,
            I => \n2527_cascade_\
        );

    \I__3274\ : CascadeMux
    port map (
            O => \N__26037\,
            I => \N__26034\
        );

    \I__3273\ : InMux
    port map (
            O => \N__26034\,
            I => \N__26030\
        );

    \I__3272\ : CascadeMux
    port map (
            O => \N__26033\,
            I => \N__26027\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__26030\,
            I => \N__26024\
        );

    \I__3270\ : InMux
    port map (
            O => \N__26027\,
            I => \N__26021\
        );

    \I__3269\ : Span4Mux_s2_h
    port map (
            O => \N__26024\,
            I => \N__26018\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__26021\,
            I => \N__26014\
        );

    \I__3267\ : Span4Mux_v
    port map (
            O => \N__26018\,
            I => \N__26011\
        );

    \I__3266\ : InMux
    port map (
            O => \N__26017\,
            I => \N__26008\
        );

    \I__3265\ : Span4Mux_s2_h
    port map (
            O => \N__26014\,
            I => \N__26003\
        );

    \I__3264\ : Span4Mux_v
    port map (
            O => \N__26011\,
            I => \N__26003\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__26008\,
            I => n2626
        );

    \I__3262\ : Odrv4
    port map (
            O => \N__26003\,
            I => n2626
        );

    \I__3261\ : CascadeMux
    port map (
            O => \N__25998\,
            I => \N__25994\
        );

    \I__3260\ : InMux
    port map (
            O => \N__25997\,
            I => \N__25991\
        );

    \I__3259\ : InMux
    port map (
            O => \N__25994\,
            I => \N__25988\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__25991\,
            I => \N__25985\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__25988\,
            I => \N__25982\
        );

    \I__3256\ : Span4Mux_s3_h
    port map (
            O => \N__25985\,
            I => \N__25979\
        );

    \I__3255\ : Span4Mux_s3_h
    port map (
            O => \N__25982\,
            I => \N__25974\
        );

    \I__3254\ : Span4Mux_v
    port map (
            O => \N__25979\,
            I => \N__25974\
        );

    \I__3253\ : Odrv4
    port map (
            O => \N__25974\,
            I => n2617
        );

    \I__3252\ : CascadeMux
    port map (
            O => \N__25971\,
            I => \N__25968\
        );

    \I__3251\ : InMux
    port map (
            O => \N__25968\,
            I => \N__25965\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__25965\,
            I => \N__25960\
        );

    \I__3249\ : CascadeMux
    port map (
            O => \N__25964\,
            I => \N__25957\
        );

    \I__3248\ : InMux
    port map (
            O => \N__25963\,
            I => \N__25954\
        );

    \I__3247\ : Span4Mux_s3_h
    port map (
            O => \N__25960\,
            I => \N__25951\
        );

    \I__3246\ : InMux
    port map (
            O => \N__25957\,
            I => \N__25948\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__25954\,
            I => \N__25945\
        );

    \I__3244\ : Span4Mux_v
    port map (
            O => \N__25951\,
            I => \N__25942\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__25948\,
            I => n2625
        );

    \I__3242\ : Odrv4
    port map (
            O => \N__25945\,
            I => n2625
        );

    \I__3241\ : Odrv4
    port map (
            O => \N__25942\,
            I => n2625
        );

    \I__3240\ : CascadeMux
    port map (
            O => \N__25935\,
            I => \n2617_cascade_\
        );

    \I__3239\ : InMux
    port map (
            O => \N__25932\,
            I => \N__25929\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__25929\,
            I => n14812
        );

    \I__3237\ : InMux
    port map (
            O => \N__25926\,
            I => \N__25923\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__25923\,
            I => \N__25920\
        );

    \I__3235\ : Odrv4
    port map (
            O => \N__25920\,
            I => n2382
        );

    \I__3234\ : InMux
    port map (
            O => \N__25917\,
            I => \N__25914\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__25914\,
            I => \N__25911\
        );

    \I__3232\ : Span4Mux_h
    port map (
            O => \N__25911\,
            I => \N__25908\
        );

    \I__3231\ : Odrv4
    port map (
            O => \N__25908\,
            I => n2396
        );

    \I__3230\ : CascadeMux
    port map (
            O => \N__25905\,
            I => \N__25901\
        );

    \I__3229\ : CascadeMux
    port map (
            O => \N__25904\,
            I => \N__25898\
        );

    \I__3228\ : InMux
    port map (
            O => \N__25901\,
            I => \N__25895\
        );

    \I__3227\ : InMux
    port map (
            O => \N__25898\,
            I => \N__25891\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__25895\,
            I => \N__25888\
        );

    \I__3225\ : InMux
    port map (
            O => \N__25894\,
            I => \N__25885\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__25891\,
            I => \N__25882\
        );

    \I__3223\ : Odrv4
    port map (
            O => \N__25888\,
            I => n2329
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__25885\,
            I => n2329
        );

    \I__3221\ : Odrv4
    port map (
            O => \N__25882\,
            I => n2329
        );

    \I__3220\ : CascadeMux
    port map (
            O => \N__25875\,
            I => \N__25871\
        );

    \I__3219\ : InMux
    port map (
            O => \N__25874\,
            I => \N__25868\
        );

    \I__3218\ : InMux
    port map (
            O => \N__25871\,
            I => \N__25865\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__25868\,
            I => \N__25861\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__25865\,
            I => \N__25858\
        );

    \I__3215\ : InMux
    port map (
            O => \N__25864\,
            I => \N__25855\
        );

    \I__3214\ : Odrv4
    port map (
            O => \N__25861\,
            I => n2328
        );

    \I__3213\ : Odrv4
    port map (
            O => \N__25858\,
            I => n2328
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__25855\,
            I => n2328
        );

    \I__3211\ : InMux
    port map (
            O => \N__25848\,
            I => \N__25845\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__25845\,
            I => \N__25842\
        );

    \I__3209\ : Span4Mux_h
    port map (
            O => \N__25842\,
            I => \N__25839\
        );

    \I__3208\ : Odrv4
    port map (
            O => \N__25839\,
            I => n2395
        );

    \I__3207\ : CascadeMux
    port map (
            O => \N__25836\,
            I => \n2427_cascade_\
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__25833\,
            I => \n14620_cascade_\
        );

    \I__3205\ : CascadeMux
    port map (
            O => \N__25830\,
            I => \n2526_cascade_\
        );

    \I__3204\ : InMux
    port map (
            O => \N__25827\,
            I => \N__25824\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__25824\,
            I => \N__25821\
        );

    \I__3202\ : Odrv4
    port map (
            O => \N__25821\,
            I => n14816
        );

    \I__3201\ : InMux
    port map (
            O => \N__25818\,
            I => \N__25815\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__25815\,
            I => n14392
        );

    \I__3199\ : CascadeMux
    port map (
            O => \N__25812\,
            I => \N__25809\
        );

    \I__3198\ : InMux
    port map (
            O => \N__25809\,
            I => \N__25806\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__25806\,
            I => \N__25802\
        );

    \I__3196\ : InMux
    port map (
            O => \N__25805\,
            I => \N__25799\
        );

    \I__3195\ : Span4Mux_v
    port map (
            O => \N__25802\,
            I => \N__25796\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__25799\,
            I => \N__25793\
        );

    \I__3193\ : Span4Mux_v
    port map (
            O => \N__25796\,
            I => \N__25788\
        );

    \I__3192\ : Span4Mux_v
    port map (
            O => \N__25793\,
            I => \N__25788\
        );

    \I__3191\ : Odrv4
    port map (
            O => \N__25788\,
            I => n2313
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__25785\,
            I => \n14398_cascade_\
        );

    \I__3189\ : CascadeMux
    port map (
            O => \N__25782\,
            I => \N__25779\
        );

    \I__3188\ : InMux
    port map (
            O => \N__25779\,
            I => \N__25775\
        );

    \I__3187\ : InMux
    port map (
            O => \N__25778\,
            I => \N__25771\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__25775\,
            I => \N__25768\
        );

    \I__3185\ : InMux
    port map (
            O => \N__25774\,
            I => \N__25765\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__25771\,
            I => n2327
        );

    \I__3183\ : Odrv4
    port map (
            O => \N__25768\,
            I => n2327
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__25765\,
            I => n2327
        );

    \I__3181\ : CascadeMux
    port map (
            O => \N__25758\,
            I => \n2346_cascade_\
        );

    \I__3180\ : InMux
    port map (
            O => \N__25755\,
            I => \N__25752\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__25752\,
            I => \N__25749\
        );

    \I__3178\ : Span4Mux_h
    port map (
            O => \N__25749\,
            I => \N__25746\
        );

    \I__3177\ : Odrv4
    port map (
            O => \N__25746\,
            I => n2394
        );

    \I__3176\ : InMux
    port map (
            O => \N__25743\,
            I => \N__25740\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__25740\,
            I => \N__25737\
        );

    \I__3174\ : Span4Mux_v
    port map (
            O => \N__25737\,
            I => \N__25734\
        );

    \I__3173\ : Odrv4
    port map (
            O => \N__25734\,
            I => n2284
        );

    \I__3172\ : InMux
    port map (
            O => \N__25731\,
            I => \N__25728\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__25728\,
            I => \N__25724\
        );

    \I__3170\ : InMux
    port map (
            O => \N__25727\,
            I => \N__25720\
        );

    \I__3169\ : Span4Mux_h
    port map (
            O => \N__25724\,
            I => \N__25717\
        );

    \I__3168\ : InMux
    port map (
            O => \N__25723\,
            I => \N__25714\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__25720\,
            I => n2316
        );

    \I__3166\ : Odrv4
    port map (
            O => \N__25717\,
            I => n2316
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__25714\,
            I => n2316
        );

    \I__3164\ : InMux
    port map (
            O => \N__25707\,
            I => \N__25704\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__25704\,
            I => \N__25701\
        );

    \I__3162\ : Span4Mux_v
    port map (
            O => \N__25701\,
            I => \N__25698\
        );

    \I__3161\ : Odrv4
    port map (
            O => \N__25698\,
            I => n2282
        );

    \I__3160\ : InMux
    port map (
            O => \N__25695\,
            I => \N__25692\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__25692\,
            I => \N__25689\
        );

    \I__3158\ : Span4Mux_v
    port map (
            O => \N__25689\,
            I => \N__25685\
        );

    \I__3157\ : InMux
    port map (
            O => \N__25688\,
            I => \N__25682\
        );

    \I__3156\ : Odrv4
    port map (
            O => \N__25685\,
            I => n2314
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__25682\,
            I => n2314
        );

    \I__3154\ : CascadeMux
    port map (
            O => \N__25677\,
            I => \n2314_cascade_\
        );

    \I__3153\ : InMux
    port map (
            O => \N__25674\,
            I => \N__25671\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__25671\,
            I => \N__25668\
        );

    \I__3151\ : Span4Mux_h
    port map (
            O => \N__25668\,
            I => \N__25665\
        );

    \I__3150\ : Odrv4
    port map (
            O => \N__25665\,
            I => n2381
        );

    \I__3149\ : InMux
    port map (
            O => \N__25662\,
            I => \N__25659\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__25659\,
            I => \N__25656\
        );

    \I__3147\ : Odrv4
    port map (
            O => \N__25656\,
            I => n2392
        );

    \I__3146\ : CascadeMux
    port map (
            O => \N__25653\,
            I => \N__25649\
        );

    \I__3145\ : CascadeMux
    port map (
            O => \N__25652\,
            I => \N__25646\
        );

    \I__3144\ : InMux
    port map (
            O => \N__25649\,
            I => \N__25643\
        );

    \I__3143\ : InMux
    port map (
            O => \N__25646\,
            I => \N__25640\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__25643\,
            I => \N__25637\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__25640\,
            I => \N__25631\
        );

    \I__3140\ : Span4Mux_s3_h
    port map (
            O => \N__25637\,
            I => \N__25631\
        );

    \I__3139\ : InMux
    port map (
            O => \N__25636\,
            I => \N__25628\
        );

    \I__3138\ : Odrv4
    port map (
            O => \N__25631\,
            I => n2325
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__25628\,
            I => n2325
        );

    \I__3136\ : InMux
    port map (
            O => \N__25623\,
            I => \N__25619\
        );

    \I__3135\ : InMux
    port map (
            O => \N__25622\,
            I => \N__25615\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__25619\,
            I => \N__25612\
        );

    \I__3133\ : InMux
    port map (
            O => \N__25618\,
            I => \N__25609\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__25615\,
            I => n2320
        );

    \I__3131\ : Odrv4
    port map (
            O => \N__25612\,
            I => n2320
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__25609\,
            I => n2320
        );

    \I__3129\ : InMux
    port map (
            O => \N__25602\,
            I => \N__25599\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__25599\,
            I => \N__25596\
        );

    \I__3127\ : Odrv12
    port map (
            O => \N__25596\,
            I => n2387
        );

    \I__3126\ : InMux
    port map (
            O => \N__25593\,
            I => n12671
        );

    \I__3125\ : InMux
    port map (
            O => \N__25590\,
            I => \bfn_4_19_0_\
        );

    \I__3124\ : InMux
    port map (
            O => \N__25587\,
            I => n12673
        );

    \I__3123\ : InMux
    port map (
            O => \N__25584\,
            I => n12674
        );

    \I__3122\ : InMux
    port map (
            O => \N__25581\,
            I => n12675
        );

    \I__3121\ : InMux
    port map (
            O => \N__25578\,
            I => \N__25575\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__25575\,
            I => \N__25571\
        );

    \I__3119\ : InMux
    port map (
            O => \N__25574\,
            I => \N__25568\
        );

    \I__3118\ : Odrv4
    port map (
            O => \N__25571\,
            I => n2214
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__25568\,
            I => n2214
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__25563\,
            I => \N__25560\
        );

    \I__3115\ : InMux
    port map (
            O => \N__25560\,
            I => \N__25557\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__25557\,
            I => \N__25554\
        );

    \I__3113\ : Span4Mux_v
    port map (
            O => \N__25554\,
            I => \N__25551\
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__25551\,
            I => n2294
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__25548\,
            I => \N__25545\
        );

    \I__3110\ : InMux
    port map (
            O => \N__25545\,
            I => \N__25542\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__25542\,
            I => n2186
        );

    \I__3108\ : CascadeMux
    port map (
            O => \N__25539\,
            I => \N__25536\
        );

    \I__3107\ : InMux
    port map (
            O => \N__25536\,
            I => \N__25533\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__25533\,
            I => \N__25530\
        );

    \I__3105\ : Span4Mux_v
    port map (
            O => \N__25530\,
            I => \N__25526\
        );

    \I__3104\ : InMux
    port map (
            O => \N__25529\,
            I => \N__25523\
        );

    \I__3103\ : Odrv4
    port map (
            O => \N__25526\,
            I => n2218
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__25523\,
            I => n2218
        );

    \I__3101\ : InMux
    port map (
            O => \N__25518\,
            I => \N__25515\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__25515\,
            I => \N__25512\
        );

    \I__3099\ : Span4Mux_v
    port map (
            O => \N__25512\,
            I => \N__25509\
        );

    \I__3098\ : Odrv4
    port map (
            O => \N__25509\,
            I => n2285
        );

    \I__3097\ : CascadeMux
    port map (
            O => \N__25506\,
            I => \n2218_cascade_\
        );

    \I__3096\ : CascadeMux
    port map (
            O => \N__25503\,
            I => \N__25500\
        );

    \I__3095\ : InMux
    port map (
            O => \N__25500\,
            I => \N__25497\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__25497\,
            I => n2188
        );

    \I__3093\ : InMux
    port map (
            O => \N__25494\,
            I => \N__25491\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__25491\,
            I => \N__25487\
        );

    \I__3091\ : InMux
    port map (
            O => \N__25490\,
            I => \N__25483\
        );

    \I__3090\ : Span4Mux_v
    port map (
            O => \N__25487\,
            I => \N__25480\
        );

    \I__3089\ : InMux
    port map (
            O => \N__25486\,
            I => \N__25477\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__25483\,
            I => n2220
        );

    \I__3087\ : Odrv4
    port map (
            O => \N__25480\,
            I => n2220
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__25477\,
            I => n2220
        );

    \I__3085\ : InMux
    port map (
            O => \N__25470\,
            I => n12662
        );

    \I__3084\ : InMux
    port map (
            O => \N__25467\,
            I => \N__25464\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__25464\,
            I => n2194
        );

    \I__3082\ : InMux
    port map (
            O => \N__25461\,
            I => n12663
        );

    \I__3081\ : InMux
    port map (
            O => \N__25458\,
            I => \N__25455\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__25455\,
            I => \N__25452\
        );

    \I__3079\ : Odrv4
    port map (
            O => \N__25452\,
            I => n2193
        );

    \I__3078\ : InMux
    port map (
            O => \N__25449\,
            I => \bfn_4_18_0_\
        );

    \I__3077\ : InMux
    port map (
            O => \N__25446\,
            I => n12665
        );

    \I__3076\ : InMux
    port map (
            O => \N__25443\,
            I => n12666
        );

    \I__3075\ : InMux
    port map (
            O => \N__25440\,
            I => \N__25437\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__25437\,
            I => n2190
        );

    \I__3073\ : InMux
    port map (
            O => \N__25434\,
            I => n12667
        );

    \I__3072\ : InMux
    port map (
            O => \N__25431\,
            I => \N__25428\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__25428\,
            I => \N__25425\
        );

    \I__3070\ : Odrv4
    port map (
            O => \N__25425\,
            I => n2189
        );

    \I__3069\ : InMux
    port map (
            O => \N__25422\,
            I => n12668
        );

    \I__3068\ : InMux
    port map (
            O => \N__25419\,
            I => n12669
        );

    \I__3067\ : InMux
    port map (
            O => \N__25416\,
            I => \N__25413\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__25413\,
            I => n2187
        );

    \I__3065\ : InMux
    port map (
            O => \N__25410\,
            I => n12670
        );

    \I__3064\ : CascadeMux
    port map (
            O => \N__25407\,
            I => \n2129_cascade_\
        );

    \I__3063\ : CascadeMux
    port map (
            O => \N__25404\,
            I => \N__25401\
        );

    \I__3062\ : InMux
    port map (
            O => \N__25401\,
            I => \N__25397\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__25400\,
            I => \N__25394\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__25397\,
            I => \N__25391\
        );

    \I__3059\ : InMux
    port map (
            O => \N__25394\,
            I => \N__25388\
        );

    \I__3058\ : Span4Mux_s3_h
    port map (
            O => \N__25391\,
            I => \N__25385\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__25388\,
            I => \N__25382\
        );

    \I__3056\ : Odrv4
    port map (
            O => \N__25385\,
            I => n2228
        );

    \I__3055\ : Odrv4
    port map (
            O => \N__25382\,
            I => n2228
        );

    \I__3054\ : InMux
    port map (
            O => \N__25377\,
            I => \N__25373\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__25376\,
            I => \N__25370\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__25373\,
            I => \N__25366\
        );

    \I__3051\ : InMux
    port map (
            O => \N__25370\,
            I => \N__25363\
        );

    \I__3050\ : InMux
    port map (
            O => \N__25369\,
            I => \N__25360\
        );

    \I__3049\ : Odrv4
    port map (
            O => \N__25366\,
            I => n2226
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__25363\,
            I => n2226
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__25360\,
            I => n2226
        );

    \I__3046\ : InMux
    port map (
            O => \N__25353\,
            I => \N__25350\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__25350\,
            I => \N__25346\
        );

    \I__3044\ : CascadeMux
    port map (
            O => \N__25349\,
            I => \N__25343\
        );

    \I__3043\ : Span4Mux_v
    port map (
            O => \N__25346\,
            I => \N__25339\
        );

    \I__3042\ : InMux
    port map (
            O => \N__25343\,
            I => \N__25336\
        );

    \I__3041\ : InMux
    port map (
            O => \N__25342\,
            I => \N__25333\
        );

    \I__3040\ : Odrv4
    port map (
            O => \N__25339\,
            I => n2225
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__25336\,
            I => n2225
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__25333\,
            I => n2225
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__25326\,
            I => \n2228_cascade_\
        );

    \I__3036\ : InMux
    port map (
            O => \N__25323\,
            I => \N__25320\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__25320\,
            I => n14588
        );

    \I__3034\ : InMux
    port map (
            O => \N__25317\,
            I => \N__25314\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__25314\,
            I => n2201
        );

    \I__3032\ : InMux
    port map (
            O => \N__25311\,
            I => \bfn_4_17_0_\
        );

    \I__3031\ : InMux
    port map (
            O => \N__25308\,
            I => \N__25305\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__25305\,
            I => \N__25302\
        );

    \I__3029\ : Odrv4
    port map (
            O => \N__25302\,
            I => n2200
        );

    \I__3028\ : InMux
    port map (
            O => \N__25299\,
            I => n12657
        );

    \I__3027\ : InMux
    port map (
            O => \N__25296\,
            I => \N__25293\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__25293\,
            I => \N__25290\
        );

    \I__3025\ : Odrv4
    port map (
            O => \N__25290\,
            I => n2199
        );

    \I__3024\ : InMux
    port map (
            O => \N__25287\,
            I => n12658
        );

    \I__3023\ : InMux
    port map (
            O => \N__25284\,
            I => n12659
        );

    \I__3022\ : InMux
    port map (
            O => \N__25281\,
            I => \N__25278\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__25278\,
            I => n2197
        );

    \I__3020\ : InMux
    port map (
            O => \N__25275\,
            I => n12660
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__25272\,
            I => \N__25268\
        );

    \I__3018\ : CascadeMux
    port map (
            O => \N__25271\,
            I => \N__25265\
        );

    \I__3017\ : InMux
    port map (
            O => \N__25268\,
            I => \N__25262\
        );

    \I__3016\ : InMux
    port map (
            O => \N__25265\,
            I => \N__25259\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__25262\,
            I => n2129
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__25259\,
            I => n2129
        );

    \I__3013\ : InMux
    port map (
            O => \N__25254\,
            I => \N__25251\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__25251\,
            I => n2196
        );

    \I__3011\ : InMux
    port map (
            O => \N__25248\,
            I => n12661
        );

    \I__3010\ : InMux
    port map (
            O => \N__25245\,
            I => \N__25242\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__25242\,
            I => n3175
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__25239\,
            I => \n3108_cascade_\
        );

    \I__3007\ : InMux
    port map (
            O => \N__25236\,
            I => \N__25232\
        );

    \I__3006\ : CascadeMux
    port map (
            O => \N__25235\,
            I => \N__25228\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__25232\,
            I => \N__25225\
        );

    \I__3004\ : InMux
    port map (
            O => \N__25231\,
            I => \N__25222\
        );

    \I__3003\ : InMux
    port map (
            O => \N__25228\,
            I => \N__25219\
        );

    \I__3002\ : Odrv4
    port map (
            O => \N__25225\,
            I => n2232
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__25222\,
            I => n2232
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__25219\,
            I => n2232
        );

    \I__2999\ : InMux
    port map (
            O => \N__25212\,
            I => \N__25209\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__25209\,
            I => \N__25205\
        );

    \I__2997\ : CascadeMux
    port map (
            O => \N__25208\,
            I => \N__25202\
        );

    \I__2996\ : Span4Mux_v
    port map (
            O => \N__25205\,
            I => \N__25198\
        );

    \I__2995\ : InMux
    port map (
            O => \N__25202\,
            I => \N__25195\
        );

    \I__2994\ : InMux
    port map (
            O => \N__25201\,
            I => \N__25192\
        );

    \I__2993\ : Odrv4
    port map (
            O => \N__25198\,
            I => n2231
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__25195\,
            I => n2231
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__25192\,
            I => n2231
        );

    \I__2990\ : CascadeMux
    port map (
            O => \N__25185\,
            I => \N__25182\
        );

    \I__2989\ : InMux
    port map (
            O => \N__25182\,
            I => \N__25179\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__25179\,
            I => \N__25174\
        );

    \I__2987\ : CascadeMux
    port map (
            O => \N__25178\,
            I => \N__25171\
        );

    \I__2986\ : CascadeMux
    port map (
            O => \N__25177\,
            I => \N__25168\
        );

    \I__2985\ : Span4Mux_v
    port map (
            O => \N__25174\,
            I => \N__25165\
        );

    \I__2984\ : InMux
    port map (
            O => \N__25171\,
            I => \N__25162\
        );

    \I__2983\ : InMux
    port map (
            O => \N__25168\,
            I => \N__25159\
        );

    \I__2982\ : Odrv4
    port map (
            O => \N__25165\,
            I => n2221
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__25162\,
            I => n2221
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__25159\,
            I => n2221
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__25152\,
            I => \N__25147\
        );

    \I__2978\ : InMux
    port map (
            O => \N__25151\,
            I => \N__25142\
        );

    \I__2977\ : InMux
    port map (
            O => \N__25150\,
            I => \N__25142\
        );

    \I__2976\ : InMux
    port map (
            O => \N__25147\,
            I => \N__25139\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__25142\,
            I => \N__25136\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__25139\,
            I => \N__25133\
        );

    \I__2973\ : Odrv4
    port map (
            O => \N__25136\,
            I => n2229
        );

    \I__2972\ : Odrv4
    port map (
            O => \N__25133\,
            I => n2229
        );

    \I__2971\ : InMux
    port map (
            O => \N__25128\,
            I => n12891
        );

    \I__2970\ : CascadeMux
    port map (
            O => \N__25125\,
            I => \N__25122\
        );

    \I__2969\ : InMux
    port map (
            O => \N__25122\,
            I => \N__25119\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__25119\,
            I => n3075
        );

    \I__2967\ : InMux
    port map (
            O => \N__25116\,
            I => \N__25113\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__25113\,
            I => n3082
        );

    \I__2965\ : CascadeMux
    port map (
            O => \N__25110\,
            I => \N__25107\
        );

    \I__2964\ : InMux
    port map (
            O => \N__25107\,
            I => \N__25104\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__25104\,
            I => n3074
        );

    \I__2962\ : InMux
    port map (
            O => \N__25101\,
            I => \N__25098\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__25098\,
            I => n3173
        );

    \I__2960\ : InMux
    port map (
            O => \N__25095\,
            I => \N__25092\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__25092\,
            I => n3174
        );

    \I__2958\ : InMux
    port map (
            O => \N__25089\,
            I => \N__25086\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__25086\,
            I => \N__25083\
        );

    \I__2956\ : Odrv4
    port map (
            O => \N__25083\,
            I => n3079
        );

    \I__2955\ : CascadeMux
    port map (
            O => \N__25080\,
            I => \N__25077\
        );

    \I__2954\ : InMux
    port map (
            O => \N__25077\,
            I => \N__25074\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__25074\,
            I => \N__25071\
        );

    \I__2952\ : Odrv4
    port map (
            O => \N__25071\,
            I => n3078
        );

    \I__2951\ : InMux
    port map (
            O => \N__25068\,
            I => \N__25065\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__25065\,
            I => n3076
        );

    \I__2949\ : InMux
    port map (
            O => \N__25062\,
            I => n12882
        );

    \I__2948\ : InMux
    port map (
            O => \N__25059\,
            I => n12883
        );

    \I__2947\ : InMux
    port map (
            O => \N__25056\,
            I => n12884
        );

    \I__2946\ : InMux
    port map (
            O => \N__25053\,
            I => n12885
        );

    \I__2945\ : InMux
    port map (
            O => \N__25050\,
            I => n12886
        );

    \I__2944\ : InMux
    port map (
            O => \N__25047\,
            I => \bfn_3_31_0_\
        );

    \I__2943\ : InMux
    port map (
            O => \N__25044\,
            I => n12888
        );

    \I__2942\ : InMux
    port map (
            O => \N__25041\,
            I => n12889
        );

    \I__2941\ : InMux
    port map (
            O => \N__25038\,
            I => n12890
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__25035\,
            I => \N__25032\
        );

    \I__2939\ : InMux
    port map (
            O => \N__25032\,
            I => \N__25029\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__25029\,
            I => \N__25026\
        );

    \I__2937\ : Span4Mux_s2_h
    port map (
            O => \N__25026\,
            I => \N__25023\
        );

    \I__2936\ : Odrv4
    port map (
            O => \N__25023\,
            I => n3090
        );

    \I__2935\ : InMux
    port map (
            O => \N__25020\,
            I => n12874
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__25017\,
            I => \N__25014\
        );

    \I__2933\ : InMux
    port map (
            O => \N__25014\,
            I => \N__25011\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__25011\,
            I => \N__25007\
        );

    \I__2931\ : InMux
    port map (
            O => \N__25010\,
            I => \N__25003\
        );

    \I__2930\ : Span4Mux_h
    port map (
            O => \N__25007\,
            I => \N__25000\
        );

    \I__2929\ : InMux
    port map (
            O => \N__25006\,
            I => \N__24997\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__25003\,
            I => n3022
        );

    \I__2927\ : Odrv4
    port map (
            O => \N__25000\,
            I => n3022
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__24997\,
            I => n3022
        );

    \I__2925\ : CascadeMux
    port map (
            O => \N__24990\,
            I => \N__24987\
        );

    \I__2924\ : InMux
    port map (
            O => \N__24987\,
            I => \N__24984\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__24984\,
            I => n3089
        );

    \I__2922\ : InMux
    port map (
            O => \N__24981\,
            I => n12875
        );

    \I__2921\ : CascadeMux
    port map (
            O => \N__24978\,
            I => \N__24974\
        );

    \I__2920\ : CascadeMux
    port map (
            O => \N__24977\,
            I => \N__24971\
        );

    \I__2919\ : InMux
    port map (
            O => \N__24974\,
            I => \N__24968\
        );

    \I__2918\ : InMux
    port map (
            O => \N__24971\,
            I => \N__24965\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__24968\,
            I => \N__24962\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__24965\,
            I => \N__24959\
        );

    \I__2915\ : Span4Mux_s1_h
    port map (
            O => \N__24962\,
            I => \N__24954\
        );

    \I__2914\ : Span4Mux_h
    port map (
            O => \N__24959\,
            I => \N__24954\
        );

    \I__2913\ : Odrv4
    port map (
            O => \N__24954\,
            I => n3021
        );

    \I__2912\ : InMux
    port map (
            O => \N__24951\,
            I => \N__24948\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__24948\,
            I => \N__24945\
        );

    \I__2910\ : Odrv4
    port map (
            O => \N__24945\,
            I => n3088
        );

    \I__2909\ : InMux
    port map (
            O => \N__24942\,
            I => n12876
        );

    \I__2908\ : CascadeMux
    port map (
            O => \N__24939\,
            I => \N__24936\
        );

    \I__2907\ : InMux
    port map (
            O => \N__24936\,
            I => \N__24931\
        );

    \I__2906\ : InMux
    port map (
            O => \N__24935\,
            I => \N__24928\
        );

    \I__2905\ : InMux
    port map (
            O => \N__24934\,
            I => \N__24925\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__24931\,
            I => \N__24922\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__24928\,
            I => \N__24919\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__24925\,
            I => n3020
        );

    \I__2901\ : Odrv4
    port map (
            O => \N__24922\,
            I => n3020
        );

    \I__2900\ : Odrv12
    port map (
            O => \N__24919\,
            I => n3020
        );

    \I__2899\ : InMux
    port map (
            O => \N__24912\,
            I => \N__24909\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__24909\,
            I => n3087
        );

    \I__2897\ : InMux
    port map (
            O => \N__24906\,
            I => n12877
        );

    \I__2896\ : InMux
    port map (
            O => \N__24903\,
            I => \N__24900\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__24900\,
            I => \N__24897\
        );

    \I__2894\ : Odrv4
    port map (
            O => \N__24897\,
            I => n3086
        );

    \I__2893\ : InMux
    port map (
            O => \N__24894\,
            I => n12878
        );

    \I__2892\ : InMux
    port map (
            O => \N__24891\,
            I => \bfn_3_30_0_\
        );

    \I__2891\ : InMux
    port map (
            O => \N__24888\,
            I => \N__24885\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__24885\,
            I => \N__24881\
        );

    \I__2889\ : InMux
    port map (
            O => \N__24884\,
            I => \N__24877\
        );

    \I__2888\ : Span4Mux_h
    port map (
            O => \N__24881\,
            I => \N__24874\
        );

    \I__2887\ : InMux
    port map (
            O => \N__24880\,
            I => \N__24871\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__24877\,
            I => n3017
        );

    \I__2885\ : Odrv4
    port map (
            O => \N__24874\,
            I => n3017
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__24871\,
            I => n3017
        );

    \I__2883\ : InMux
    port map (
            O => \N__24864\,
            I => \N__24861\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__24861\,
            I => \N__24858\
        );

    \I__2881\ : Odrv4
    port map (
            O => \N__24858\,
            I => n3084
        );

    \I__2880\ : InMux
    port map (
            O => \N__24855\,
            I => n12880
        );

    \I__2879\ : InMux
    port map (
            O => \N__24852\,
            I => n12881
        );

    \I__2878\ : InMux
    port map (
            O => \N__24849\,
            I => n12866
        );

    \I__2877\ : InMux
    port map (
            O => \N__24846\,
            I => n12867
        );

    \I__2876\ : InMux
    port map (
            O => \N__24843\,
            I => \N__24840\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__24840\,
            I => \N__24837\
        );

    \I__2874\ : Odrv12
    port map (
            O => \N__24837\,
            I => n3096
        );

    \I__2873\ : InMux
    port map (
            O => \N__24834\,
            I => n12868
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__24831\,
            I => \N__24827\
        );

    \I__2871\ : InMux
    port map (
            O => \N__24830\,
            I => \N__24824\
        );

    \I__2870\ : InMux
    port map (
            O => \N__24827\,
            I => \N__24821\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__24824\,
            I => \N__24818\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__24821\,
            I => n3028
        );

    \I__2867\ : Odrv12
    port map (
            O => \N__24818\,
            I => n3028
        );

    \I__2866\ : InMux
    port map (
            O => \N__24813\,
            I => \N__24810\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__24810\,
            I => n3095
        );

    \I__2864\ : InMux
    port map (
            O => \N__24807\,
            I => n12869
        );

    \I__2863\ : InMux
    port map (
            O => \N__24804\,
            I => \N__24801\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__24801\,
            I => \N__24798\
        );

    \I__2861\ : Odrv12
    port map (
            O => \N__24798\,
            I => n3094
        );

    \I__2860\ : InMux
    port map (
            O => \N__24795\,
            I => n12870
        );

    \I__2859\ : CascadeMux
    port map (
            O => \N__24792\,
            I => \N__24789\
        );

    \I__2858\ : InMux
    port map (
            O => \N__24789\,
            I => \N__24785\
        );

    \I__2857\ : InMux
    port map (
            O => \N__24788\,
            I => \N__24782\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__24785\,
            I => \N__24779\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__24782\,
            I => \N__24775\
        );

    \I__2854\ : Span4Mux_h
    port map (
            O => \N__24779\,
            I => \N__24772\
        );

    \I__2853\ : InMux
    port map (
            O => \N__24778\,
            I => \N__24769\
        );

    \I__2852\ : Odrv4
    port map (
            O => \N__24775\,
            I => n3026
        );

    \I__2851\ : Odrv4
    port map (
            O => \N__24772\,
            I => n3026
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__24769\,
            I => n3026
        );

    \I__2849\ : CascadeMux
    port map (
            O => \N__24762\,
            I => \N__24759\
        );

    \I__2848\ : InMux
    port map (
            O => \N__24759\,
            I => \N__24756\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__24756\,
            I => n3093
        );

    \I__2846\ : InMux
    port map (
            O => \N__24753\,
            I => \bfn_3_29_0_\
        );

    \I__2845\ : CascadeMux
    port map (
            O => \N__24750\,
            I => \N__24747\
        );

    \I__2844\ : InMux
    port map (
            O => \N__24747\,
            I => \N__24743\
        );

    \I__2843\ : InMux
    port map (
            O => \N__24746\,
            I => \N__24740\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__24743\,
            I => \N__24737\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__24740\,
            I => \N__24731\
        );

    \I__2840\ : Span4Mux_h
    port map (
            O => \N__24737\,
            I => \N__24731\
        );

    \I__2839\ : InMux
    port map (
            O => \N__24736\,
            I => \N__24728\
        );

    \I__2838\ : Odrv4
    port map (
            O => \N__24731\,
            I => n3025
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__24728\,
            I => n3025
        );

    \I__2836\ : InMux
    port map (
            O => \N__24723\,
            I => \N__24720\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__24720\,
            I => \N__24717\
        );

    \I__2834\ : Odrv4
    port map (
            O => \N__24717\,
            I => n3092
        );

    \I__2833\ : InMux
    port map (
            O => \N__24714\,
            I => n12872
        );

    \I__2832\ : CascadeMux
    port map (
            O => \N__24711\,
            I => \N__24708\
        );

    \I__2831\ : InMux
    port map (
            O => \N__24708\,
            I => \N__24704\
        );

    \I__2830\ : InMux
    port map (
            O => \N__24707\,
            I => \N__24701\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__24704\,
            I => \N__24698\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__24701\,
            I => \N__24695\
        );

    \I__2827\ : Span4Mux_v
    port map (
            O => \N__24698\,
            I => \N__24692\
        );

    \I__2826\ : Odrv12
    port map (
            O => \N__24695\,
            I => n3024
        );

    \I__2825\ : Odrv4
    port map (
            O => \N__24692\,
            I => n3024
        );

    \I__2824\ : CascadeMux
    port map (
            O => \N__24687\,
            I => \N__24684\
        );

    \I__2823\ : InMux
    port map (
            O => \N__24684\,
            I => \N__24681\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__24681\,
            I => \N__24678\
        );

    \I__2821\ : Odrv4
    port map (
            O => \N__24678\,
            I => n3091
        );

    \I__2820\ : InMux
    port map (
            O => \N__24675\,
            I => n12873
        );

    \I__2819\ : CascadeMux
    port map (
            O => \N__24672\,
            I => \n3028_cascade_\
        );

    \I__2818\ : CascadeMux
    port map (
            O => \N__24669\,
            I => \N__24666\
        );

    \I__2817\ : InMux
    port map (
            O => \N__24666\,
            I => \N__24663\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__24663\,
            I => n2988
        );

    \I__2815\ : InMux
    port map (
            O => \N__24660\,
            I => \N__24657\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__24657\,
            I => \N__24654\
        );

    \I__2813\ : Span4Mux_v
    port map (
            O => \N__24654\,
            I => \N__24651\
        );

    \I__2812\ : Odrv4
    port map (
            O => \N__24651\,
            I => n2880
        );

    \I__2811\ : InMux
    port map (
            O => \N__24648\,
            I => \N__24645\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__24645\,
            I => n2979
        );

    \I__2809\ : CascadeMux
    port map (
            O => \N__24642\,
            I => \n2912_cascade_\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__24639\,
            I => \N__24636\
        );

    \I__2807\ : InMux
    port map (
            O => \N__24636\,
            I => \N__24633\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__24633\,
            I => n2983
        );

    \I__2805\ : InMux
    port map (
            O => \N__24630\,
            I => \bfn_3_28_0_\
        );

    \I__2804\ : InMux
    port map (
            O => \N__24627\,
            I => n12864
        );

    \I__2803\ : InMux
    port map (
            O => \N__24624\,
            I => n12865
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__24621\,
            I => \N__24618\
        );

    \I__2801\ : InMux
    port map (
            O => \N__24618\,
            I => \N__24613\
        );

    \I__2800\ : InMux
    port map (
            O => \N__24617\,
            I => \N__24608\
        );

    \I__2799\ : InMux
    port map (
            O => \N__24616\,
            I => \N__24608\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__24613\,
            I => n2823
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__24608\,
            I => n2823
        );

    \I__2796\ : CascadeMux
    port map (
            O => \N__24603\,
            I => \N__24600\
        );

    \I__2795\ : InMux
    port map (
            O => \N__24600\,
            I => \N__24597\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__24597\,
            I => \N__24594\
        );

    \I__2793\ : Span4Mux_v
    port map (
            O => \N__24594\,
            I => \N__24591\
        );

    \I__2792\ : Odrv4
    port map (
            O => \N__24591\,
            I => n2890
        );

    \I__2791\ : InMux
    port map (
            O => \N__24588\,
            I => \N__24585\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__24585\,
            I => \N__24581\
        );

    \I__2789\ : CascadeMux
    port map (
            O => \N__24584\,
            I => \N__24578\
        );

    \I__2788\ : Span4Mux_v
    port map (
            O => \N__24581\,
            I => \N__24574\
        );

    \I__2787\ : InMux
    port map (
            O => \N__24578\,
            I => \N__24571\
        );

    \I__2786\ : InMux
    port map (
            O => \N__24577\,
            I => \N__24568\
        );

    \I__2785\ : Odrv4
    port map (
            O => \N__24574\,
            I => n2827
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__24571\,
            I => n2827
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__24568\,
            I => n2827
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__24561\,
            I => \N__24558\
        );

    \I__2781\ : InMux
    port map (
            O => \N__24558\,
            I => \N__24555\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__24555\,
            I => \N__24552\
        );

    \I__2779\ : Span4Mux_v
    port map (
            O => \N__24552\,
            I => \N__24549\
        );

    \I__2778\ : Odrv4
    port map (
            O => \N__24549\,
            I => n2894
        );

    \I__2777\ : InMux
    port map (
            O => \N__24546\,
            I => \N__24543\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__24543\,
            I => \N__24539\
        );

    \I__2775\ : CascadeMux
    port map (
            O => \N__24542\,
            I => \N__24536\
        );

    \I__2774\ : Span4Mux_v
    port map (
            O => \N__24539\,
            I => \N__24532\
        );

    \I__2773\ : InMux
    port map (
            O => \N__24536\,
            I => \N__24529\
        );

    \I__2772\ : InMux
    port map (
            O => \N__24535\,
            I => \N__24526\
        );

    \I__2771\ : Odrv4
    port map (
            O => \N__24532\,
            I => n2822
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__24529\,
            I => n2822
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__24526\,
            I => n2822
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__24519\,
            I => \N__24516\
        );

    \I__2767\ : InMux
    port map (
            O => \N__24516\,
            I => \N__24513\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__24513\,
            I => \N__24510\
        );

    \I__2765\ : Span4Mux_h
    port map (
            O => \N__24510\,
            I => \N__24507\
        );

    \I__2764\ : Odrv4
    port map (
            O => \N__24507\,
            I => n2889
        );

    \I__2763\ : CascadeMux
    port map (
            O => \N__24504\,
            I => \N__24501\
        );

    \I__2762\ : InMux
    port map (
            O => \N__24501\,
            I => \N__24498\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__24498\,
            I => n2982
        );

    \I__2760\ : CascadeMux
    port map (
            O => \N__24495\,
            I => \N__24492\
        );

    \I__2759\ : InMux
    port map (
            O => \N__24492\,
            I => \N__24489\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__24489\,
            I => n2986
        );

    \I__2757\ : InMux
    port map (
            O => \N__24486\,
            I => \N__24483\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__24483\,
            I => \N__24480\
        );

    \I__2755\ : Span4Mux_h
    port map (
            O => \N__24480\,
            I => \N__24477\
        );

    \I__2754\ : Span4Mux_s0_h
    port map (
            O => \N__24477\,
            I => \N__24474\
        );

    \I__2753\ : Odrv4
    port map (
            O => \N__24474\,
            I => n2879
        );

    \I__2752\ : InMux
    port map (
            O => \N__24471\,
            I => \N__24468\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__24468\,
            I => \N__24464\
        );

    \I__2750\ : InMux
    port map (
            O => \N__24467\,
            I => \N__24460\
        );

    \I__2749\ : Span4Mux_v
    port map (
            O => \N__24464\,
            I => \N__24457\
        );

    \I__2748\ : InMux
    port map (
            O => \N__24463\,
            I => \N__24454\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__24460\,
            I => \N__24451\
        );

    \I__2746\ : Odrv4
    port map (
            O => \N__24457\,
            I => n2710
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__24454\,
            I => n2710
        );

    \I__2744\ : Odrv12
    port map (
            O => \N__24451\,
            I => n2710
        );

    \I__2743\ : CascadeMux
    port map (
            O => \N__24444\,
            I => \N__24441\
        );

    \I__2742\ : InMux
    port map (
            O => \N__24441\,
            I => \N__24438\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__24438\,
            I => \N__24435\
        );

    \I__2740\ : Span4Mux_v
    port map (
            O => \N__24435\,
            I => \N__24432\
        );

    \I__2739\ : Span4Mux_v
    port map (
            O => \N__24432\,
            I => \N__24429\
        );

    \I__2738\ : Odrv4
    port map (
            O => \N__24429\,
            I => n2777
        );

    \I__2737\ : InMux
    port map (
            O => \N__24426\,
            I => \N__24423\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__24423\,
            I => \N__24420\
        );

    \I__2735\ : Odrv4
    port map (
            O => \N__24420\,
            I => n2996
        );

    \I__2734\ : InMux
    port map (
            O => \N__24417\,
            I => \N__24412\
        );

    \I__2733\ : InMux
    port map (
            O => \N__24416\,
            I => \N__24409\
        );

    \I__2732\ : InMux
    port map (
            O => \N__24415\,
            I => \N__24406\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__24412\,
            I => \N__24403\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__24409\,
            I => \N__24398\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__24406\,
            I => \N__24398\
        );

    \I__2728\ : Odrv4
    port map (
            O => \N__24403\,
            I => n2713
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__24398\,
            I => n2713
        );

    \I__2726\ : InMux
    port map (
            O => \N__24393\,
            I => \N__24390\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__24390\,
            I => \N__24387\
        );

    \I__2724\ : Span4Mux_v
    port map (
            O => \N__24387\,
            I => \N__24384\
        );

    \I__2723\ : Odrv4
    port map (
            O => \N__24384\,
            I => n2780
        );

    \I__2722\ : InMux
    port map (
            O => \N__24381\,
            I => \N__24378\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__24378\,
            I => \N__24375\
        );

    \I__2720\ : Span4Mux_v
    port map (
            O => \N__24375\,
            I => \N__24372\
        );

    \I__2719\ : Odrv4
    port map (
            O => \N__24372\,
            I => n2798
        );

    \I__2718\ : CascadeMux
    port map (
            O => \N__24369\,
            I => \N__24365\
        );

    \I__2717\ : CascadeMux
    port map (
            O => \N__24368\,
            I => \N__24362\
        );

    \I__2716\ : InMux
    port map (
            O => \N__24365\,
            I => \N__24359\
        );

    \I__2715\ : InMux
    port map (
            O => \N__24362\,
            I => \N__24356\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__24359\,
            I => \N__24353\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__24356\,
            I => \N__24349\
        );

    \I__2712\ : Span12Mux_s2_h
    port map (
            O => \N__24353\,
            I => \N__24346\
        );

    \I__2711\ : InMux
    port map (
            O => \N__24352\,
            I => \N__24343\
        );

    \I__2710\ : Odrv4
    port map (
            O => \N__24349\,
            I => n2731
        );

    \I__2709\ : Odrv12
    port map (
            O => \N__24346\,
            I => n2731
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__24343\,
            I => n2731
        );

    \I__2707\ : InMux
    port map (
            O => \N__24336\,
            I => \N__24333\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__24333\,
            I => \N__24330\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__24330\,
            I => \N__24327\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__24327\,
            I => \N__24324\
        );

    \I__2703\ : Odrv4
    port map (
            O => \N__24324\,
            I => n2680
        );

    \I__2702\ : InMux
    port map (
            O => \N__24321\,
            I => \N__24318\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__24318\,
            I => \N__24315\
        );

    \I__2700\ : Span4Mux_h
    port map (
            O => \N__24315\,
            I => \N__24312\
        );

    \I__2699\ : Odrv4
    port map (
            O => \N__24312\,
            I => n2887
        );

    \I__2698\ : InMux
    port map (
            O => \N__24309\,
            I => \N__24304\
        );

    \I__2697\ : InMux
    port map (
            O => \N__24308\,
            I => \N__24299\
        );

    \I__2696\ : InMux
    port map (
            O => \N__24307\,
            I => \N__24299\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__24304\,
            I => n2820
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__24299\,
            I => n2820
        );

    \I__2693\ : CascadeMux
    port map (
            O => \N__24294\,
            I => \n14690_cascade_\
        );

    \I__2692\ : InMux
    port map (
            O => \N__24291\,
            I => \N__24288\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__24288\,
            I => \N__24285\
        );

    \I__2690\ : Odrv4
    port map (
            O => \N__24285\,
            I => n14688
        );

    \I__2689\ : CascadeMux
    port map (
            O => \N__24282\,
            I => \n14696_cascade_\
        );

    \I__2688\ : InMux
    port map (
            O => \N__24279\,
            I => \N__24274\
        );

    \I__2687\ : InMux
    port map (
            O => \N__24278\,
            I => \N__24271\
        );

    \I__2686\ : InMux
    port map (
            O => \N__24277\,
            I => \N__24268\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__24274\,
            I => \N__24265\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__24271\,
            I => \N__24262\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__24268\,
            I => \N__24259\
        );

    \I__2682\ : Span4Mux_v
    port map (
            O => \N__24265\,
            I => \N__24256\
        );

    \I__2681\ : Span4Mux_h
    port map (
            O => \N__24262\,
            I => \N__24253\
        );

    \I__2680\ : Odrv4
    port map (
            O => \N__24259\,
            I => n2714
        );

    \I__2679\ : Odrv4
    port map (
            O => \N__24256\,
            I => n2714
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__24253\,
            I => n2714
        );

    \I__2677\ : CascadeMux
    port map (
            O => \N__24246\,
            I => \N__24243\
        );

    \I__2676\ : InMux
    port map (
            O => \N__24243\,
            I => \N__24240\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__24240\,
            I => \N__24237\
        );

    \I__2674\ : Span4Mux_v
    port map (
            O => \N__24237\,
            I => \N__24234\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__24234\,
            I => n2781
        );

    \I__2672\ : InMux
    port map (
            O => \N__24231\,
            I => \N__24228\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__24228\,
            I => \N__24224\
        );

    \I__2670\ : InMux
    port map (
            O => \N__24227\,
            I => \N__24221\
        );

    \I__2669\ : Span4Mux_v
    port map (
            O => \N__24224\,
            I => \N__24217\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__24221\,
            I => \N__24214\
        );

    \I__2667\ : InMux
    port map (
            O => \N__24220\,
            I => \N__24211\
        );

    \I__2666\ : Odrv4
    port map (
            O => \N__24217\,
            I => n2720
        );

    \I__2665\ : Odrv4
    port map (
            O => \N__24214\,
            I => n2720
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__24211\,
            I => n2720
        );

    \I__2663\ : CascadeMux
    port map (
            O => \N__24204\,
            I => \N__24201\
        );

    \I__2662\ : InMux
    port map (
            O => \N__24201\,
            I => \N__24198\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__24198\,
            I => \N__24195\
        );

    \I__2660\ : Span4Mux_v
    port map (
            O => \N__24195\,
            I => \N__24192\
        );

    \I__2659\ : Odrv4
    port map (
            O => \N__24192\,
            I => n2787
        );

    \I__2658\ : CascadeMux
    port map (
            O => \N__24189\,
            I => \n14660_cascade_\
        );

    \I__2657\ : InMux
    port map (
            O => \N__24186\,
            I => \N__24183\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__24183\,
            I => n14674
        );

    \I__2655\ : CascadeMux
    port map (
            O => \N__24180\,
            I => \n2643_cascade_\
        );

    \I__2654\ : InMux
    port map (
            O => \N__24177\,
            I => \N__24174\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__24174\,
            I => \N__24171\
        );

    \I__2652\ : Span12Mux_v
    port map (
            O => \N__24171\,
            I => \N__24168\
        );

    \I__2651\ : Odrv12
    port map (
            O => \N__24168\,
            I => n2686
        );

    \I__2650\ : InMux
    port map (
            O => \N__24165\,
            I => \N__24162\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__24162\,
            I => \N__24159\
        );

    \I__2648\ : Span4Mux_v
    port map (
            O => \N__24159\,
            I => \N__24154\
        );

    \I__2647\ : InMux
    port map (
            O => \N__24158\,
            I => \N__24149\
        );

    \I__2646\ : InMux
    port map (
            O => \N__24157\,
            I => \N__24149\
        );

    \I__2645\ : Odrv4
    port map (
            O => \N__24154\,
            I => n2718
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__24149\,
            I => n2718
        );

    \I__2643\ : InMux
    port map (
            O => \N__24144\,
            I => \N__24141\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__24141\,
            I => \N__24138\
        );

    \I__2641\ : Span4Mux_v
    port map (
            O => \N__24138\,
            I => \N__24135\
        );

    \I__2640\ : Span4Mux_v
    port map (
            O => \N__24135\,
            I => \N__24132\
        );

    \I__2639\ : Odrv4
    port map (
            O => \N__24132\,
            I => n2690
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__24129\,
            I => \N__24125\
        );

    \I__2637\ : InMux
    port map (
            O => \N__24128\,
            I => \N__24121\
        );

    \I__2636\ : InMux
    port map (
            O => \N__24125\,
            I => \N__24116\
        );

    \I__2635\ : InMux
    port map (
            O => \N__24124\,
            I => \N__24116\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__24121\,
            I => \N__24113\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__24116\,
            I => \N__24110\
        );

    \I__2632\ : Span4Mux_v
    port map (
            O => \N__24113\,
            I => \N__24107\
        );

    \I__2631\ : Odrv4
    port map (
            O => \N__24110\,
            I => n2623
        );

    \I__2630\ : Odrv4
    port map (
            O => \N__24107\,
            I => n2623
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__24102\,
            I => \N__24099\
        );

    \I__2628\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24096\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__24096\,
            I => \N__24093\
        );

    \I__2626\ : Span12Mux_s2_h
    port map (
            O => \N__24093\,
            I => \N__24088\
        );

    \I__2625\ : InMux
    port map (
            O => \N__24092\,
            I => \N__24083\
        );

    \I__2624\ : InMux
    port map (
            O => \N__24091\,
            I => \N__24083\
        );

    \I__2623\ : Odrv12
    port map (
            O => \N__24088\,
            I => n2722
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__24083\,
            I => n2722
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__24078\,
            I => \N__24075\
        );

    \I__2620\ : InMux
    port map (
            O => \N__24075\,
            I => \N__24071\
        );

    \I__2619\ : InMux
    port map (
            O => \N__24074\,
            I => \N__24068\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__24071\,
            I => \N__24065\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__24068\,
            I => \N__24062\
        );

    \I__2616\ : Span4Mux_v
    port map (
            O => \N__24065\,
            I => \N__24059\
        );

    \I__2615\ : Odrv4
    port map (
            O => \N__24062\,
            I => n2732
        );

    \I__2614\ : Odrv4
    port map (
            O => \N__24059\,
            I => n2732
        );

    \I__2613\ : CascadeMux
    port map (
            O => \N__24054\,
            I => \N__24051\
        );

    \I__2612\ : InMux
    port map (
            O => \N__24051\,
            I => \N__24048\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__24048\,
            I => \N__24045\
        );

    \I__2610\ : Span4Mux_v
    port map (
            O => \N__24045\,
            I => \N__24042\
        );

    \I__2609\ : Odrv4
    port map (
            O => \N__24042\,
            I => n2799
        );

    \I__2608\ : InMux
    port map (
            O => \N__24039\,
            I => \N__24036\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__24036\,
            I => \N__24032\
        );

    \I__2606\ : InMux
    port map (
            O => \N__24035\,
            I => \N__24029\
        );

    \I__2605\ : Span4Mux_v
    port map (
            O => \N__24032\,
            I => \N__24026\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__24029\,
            I => n2711
        );

    \I__2603\ : Odrv4
    port map (
            O => \N__24026\,
            I => n2711
        );

    \I__2602\ : InMux
    port map (
            O => \N__24021\,
            I => \N__24018\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__24018\,
            I => \N__24015\
        );

    \I__2600\ : Span4Mux_h
    port map (
            O => \N__24015\,
            I => \N__24012\
        );

    \I__2599\ : Span4Mux_s1_h
    port map (
            O => \N__24012\,
            I => \N__24009\
        );

    \I__2598\ : Span4Mux_v
    port map (
            O => \N__24009\,
            I => \N__24006\
        );

    \I__2597\ : Odrv4
    port map (
            O => \N__24006\,
            I => n2778
        );

    \I__2596\ : InMux
    port map (
            O => \N__24003\,
            I => \N__24000\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__24000\,
            I => \N__23997\
        );

    \I__2594\ : Span4Mux_v
    port map (
            O => \N__23997\,
            I => \N__23994\
        );

    \I__2593\ : Odrv4
    port map (
            O => \N__23994\,
            I => n2786
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__23991\,
            I => \N__23987\
        );

    \I__2591\ : InMux
    port map (
            O => \N__23990\,
            I => \N__23984\
        );

    \I__2590\ : InMux
    port map (
            O => \N__23987\,
            I => \N__23980\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__23984\,
            I => \N__23977\
        );

    \I__2588\ : InMux
    port map (
            O => \N__23983\,
            I => \N__23974\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__23980\,
            I => n2719
        );

    \I__2586\ : Odrv12
    port map (
            O => \N__23977\,
            I => n2719
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__23974\,
            I => n2719
        );

    \I__2584\ : InMux
    port map (
            O => \N__23967\,
            I => \N__23964\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__23964\,
            I => \N__23961\
        );

    \I__2582\ : Span4Mux_v
    port map (
            O => \N__23961\,
            I => \N__23958\
        );

    \I__2581\ : Span4Mux_v
    port map (
            O => \N__23958\,
            I => \N__23955\
        );

    \I__2580\ : Odrv4
    port map (
            O => \N__23955\,
            I => n2685
        );

    \I__2579\ : InMux
    port map (
            O => \N__23952\,
            I => \N__23949\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__23949\,
            I => \N__23946\
        );

    \I__2577\ : Span4Mux_v
    port map (
            O => \N__23946\,
            I => \N__23942\
        );

    \I__2576\ : InMux
    port map (
            O => \N__23945\,
            I => \N__23939\
        );

    \I__2575\ : Odrv4
    port map (
            O => \N__23942\,
            I => n2717
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__23939\,
            I => n2717
        );

    \I__2573\ : InMux
    port map (
            O => \N__23934\,
            I => \N__23931\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__23931\,
            I => \N__23928\
        );

    \I__2571\ : Span4Mux_v
    port map (
            O => \N__23928\,
            I => \N__23925\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__23925\,
            I => n2784
        );

    \I__2569\ : CascadeMux
    port map (
            O => \N__23922\,
            I => \n2717_cascade_\
        );

    \I__2568\ : CascadeMux
    port map (
            O => \N__23919\,
            I => \n2732_cascade_\
        );

    \I__2567\ : InMux
    port map (
            O => \N__23916\,
            I => \N__23912\
        );

    \I__2566\ : InMux
    port map (
            O => \N__23915\,
            I => \N__23909\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__23912\,
            I => \N__23906\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__23909\,
            I => \N__23902\
        );

    \I__2563\ : Span4Mux_v
    port map (
            O => \N__23906\,
            I => \N__23899\
        );

    \I__2562\ : InMux
    port map (
            O => \N__23905\,
            I => \N__23896\
        );

    \I__2561\ : Odrv4
    port map (
            O => \N__23902\,
            I => n2729
        );

    \I__2560\ : Odrv4
    port map (
            O => \N__23899\,
            I => n2729
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__23896\,
            I => n2729
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__23889\,
            I => \n11957_cascade_\
        );

    \I__2557\ : InMux
    port map (
            O => \N__23886\,
            I => \N__23883\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__23883\,
            I => n13808
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__23880\,
            I => \N__23877\
        );

    \I__2554\ : InMux
    port map (
            O => \N__23877\,
            I => \N__23874\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__23874\,
            I => \N__23871\
        );

    \I__2552\ : Span4Mux_v
    port map (
            O => \N__23871\,
            I => \N__23867\
        );

    \I__2551\ : InMux
    port map (
            O => \N__23870\,
            I => \N__23864\
        );

    \I__2550\ : Odrv4
    port map (
            O => \N__23867\,
            I => n2621
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__23864\,
            I => n2621
        );

    \I__2548\ : InMux
    port map (
            O => \N__23859\,
            I => \N__23856\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__23856\,
            I => n14668
        );

    \I__2546\ : InMux
    port map (
            O => \N__23853\,
            I => \N__23850\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__23850\,
            I => \N__23847\
        );

    \I__2544\ : Span4Mux_v
    port map (
            O => \N__23847\,
            I => \N__23844\
        );

    \I__2543\ : Span4Mux_v
    port map (
            O => \N__23844\,
            I => \N__23841\
        );

    \I__2542\ : Odrv4
    port map (
            O => \N__23841\,
            I => n2698
        );

    \I__2541\ : CascadeMux
    port map (
            O => \N__23838\,
            I => \N__23835\
        );

    \I__2540\ : InMux
    port map (
            O => \N__23835\,
            I => \N__23832\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__23832\,
            I => \N__23828\
        );

    \I__2538\ : InMux
    port map (
            O => \N__23831\,
            I => \N__23824\
        );

    \I__2537\ : Span4Mux_v
    port map (
            O => \N__23828\,
            I => \N__23821\
        );

    \I__2536\ : InMux
    port map (
            O => \N__23827\,
            I => \N__23818\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__23824\,
            I => n2730
        );

    \I__2534\ : Odrv4
    port map (
            O => \N__23821\,
            I => n2730
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__23818\,
            I => n2730
        );

    \I__2532\ : InMux
    port map (
            O => \N__23811\,
            I => \N__23808\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__23808\,
            I => \N__23805\
        );

    \I__2530\ : Span4Mux_v
    port map (
            O => \N__23805\,
            I => \N__23802\
        );

    \I__2529\ : Span4Mux_v
    port map (
            O => \N__23802\,
            I => \N__23799\
        );

    \I__2528\ : Odrv4
    port map (
            O => \N__23799\,
            I => n2699
        );

    \I__2527\ : InMux
    port map (
            O => \N__23796\,
            I => \N__23793\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__23793\,
            I => \N__23790\
        );

    \I__2525\ : Span4Mux_h
    port map (
            O => \N__23790\,
            I => \N__23787\
        );

    \I__2524\ : Span4Mux_v
    port map (
            O => \N__23787\,
            I => \N__23784\
        );

    \I__2523\ : Span4Mux_v
    port map (
            O => \N__23784\,
            I => \N__23781\
        );

    \I__2522\ : Odrv4
    port map (
            O => \N__23781\,
            I => n2701
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__23778\,
            I => \n14650_cascade_\
        );

    \I__2520\ : CascadeMux
    port map (
            O => \N__23775\,
            I => \n14654_cascade_\
        );

    \I__2519\ : InMux
    port map (
            O => \N__23772\,
            I => \N__23769\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__23769\,
            I => \N__23766\
        );

    \I__2517\ : Span4Mux_v
    port map (
            O => \N__23766\,
            I => \N__23763\
        );

    \I__2516\ : Odrv4
    port map (
            O => \N__23763\,
            I => n2689
        );

    \I__2515\ : CascadeMux
    port map (
            O => \N__23760\,
            I => \n2622_cascade_\
        );

    \I__2514\ : InMux
    port map (
            O => \N__23757\,
            I => \N__23753\
        );

    \I__2513\ : CascadeMux
    port map (
            O => \N__23756\,
            I => \N__23750\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__23753\,
            I => \N__23747\
        );

    \I__2511\ : InMux
    port map (
            O => \N__23750\,
            I => \N__23744\
        );

    \I__2510\ : Span4Mux_v
    port map (
            O => \N__23747\,
            I => \N__23741\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__23744\,
            I => \N__23738\
        );

    \I__2508\ : Odrv4
    port map (
            O => \N__23741\,
            I => n2721
        );

    \I__2507\ : Odrv4
    port map (
            O => \N__23738\,
            I => n2721
        );

    \I__2506\ : CascadeMux
    port map (
            O => \N__23733\,
            I => \N__23730\
        );

    \I__2505\ : InMux
    port map (
            O => \N__23730\,
            I => \N__23727\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__23727\,
            I => \N__23723\
        );

    \I__2503\ : InMux
    port map (
            O => \N__23726\,
            I => \N__23720\
        );

    \I__2502\ : Odrv12
    port map (
            O => \N__23723\,
            I => n2728
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__23720\,
            I => n2728
        );

    \I__2500\ : CascadeMux
    port map (
            O => \N__23715\,
            I => \N__23712\
        );

    \I__2499\ : InMux
    port map (
            O => \N__23712\,
            I => \N__23709\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__23709\,
            I => \N__23705\
        );

    \I__2497\ : InMux
    port map (
            O => \N__23708\,
            I => \N__23702\
        );

    \I__2496\ : Odrv4
    port map (
            O => \N__23705\,
            I => n2726
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__23702\,
            I => n2726
        );

    \I__2494\ : CascadeMux
    port map (
            O => \N__23697\,
            I => \n2721_cascade_\
        );

    \I__2493\ : InMux
    port map (
            O => \N__23694\,
            I => \N__23691\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__23691\,
            I => \N__23688\
        );

    \I__2491\ : Odrv4
    port map (
            O => \N__23688\,
            I => n14348
        );

    \I__2490\ : InMux
    port map (
            O => \N__23685\,
            I => \N__23682\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__23682\,
            I => \N__23679\
        );

    \I__2488\ : Odrv4
    port map (
            O => \N__23679\,
            I => n2383
        );

    \I__2487\ : CascadeMux
    port map (
            O => \N__23676\,
            I => \N__23673\
        );

    \I__2486\ : InMux
    port map (
            O => \N__23673\,
            I => \N__23670\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__23670\,
            I => \N__23667\
        );

    \I__2484\ : Span4Mux_v
    port map (
            O => \N__23667\,
            I => \N__23663\
        );

    \I__2483\ : InMux
    port map (
            O => \N__23666\,
            I => \N__23660\
        );

    \I__2482\ : Odrv4
    port map (
            O => \N__23663\,
            I => n2622
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__23660\,
            I => n2622
        );

    \I__2480\ : CascadeMux
    port map (
            O => \N__23655\,
            I => \n2628_cascade_\
        );

    \I__2479\ : InMux
    port map (
            O => \N__23652\,
            I => \N__23649\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__23649\,
            I => \N__23646\
        );

    \I__2477\ : Span4Mux_v
    port map (
            O => \N__23646\,
            I => \N__23643\
        );

    \I__2476\ : Span4Mux_v
    port map (
            O => \N__23643\,
            I => \N__23640\
        );

    \I__2475\ : Odrv4
    port map (
            O => \N__23640\,
            I => n2692
        );

    \I__2474\ : CascadeMux
    port map (
            O => \N__23637\,
            I => \N__23633\
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__23636\,
            I => \N__23630\
        );

    \I__2472\ : InMux
    port map (
            O => \N__23633\,
            I => \N__23627\
        );

    \I__2471\ : InMux
    port map (
            O => \N__23630\,
            I => \N__23624\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__23627\,
            I => \N__23621\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__23624\,
            I => \N__23617\
        );

    \I__2468\ : Span4Mux_s3_h
    port map (
            O => \N__23621\,
            I => \N__23614\
        );

    \I__2467\ : InMux
    port map (
            O => \N__23620\,
            I => \N__23611\
        );

    \I__2466\ : Odrv4
    port map (
            O => \N__23617\,
            I => n2724
        );

    \I__2465\ : Odrv4
    port map (
            O => \N__23614\,
            I => n2724
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__23611\,
            I => n2724
        );

    \I__2463\ : InMux
    port map (
            O => \N__23604\,
            I => \N__23601\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__23601\,
            I => \N__23598\
        );

    \I__2461\ : Span4Mux_v
    port map (
            O => \N__23598\,
            I => \N__23595\
        );

    \I__2460\ : Span4Mux_v
    port map (
            O => \N__23595\,
            I => \N__23592\
        );

    \I__2459\ : Odrv4
    port map (
            O => \N__23592\,
            I => n2695
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__23589\,
            I => \N__23586\
        );

    \I__2457\ : InMux
    port map (
            O => \N__23586\,
            I => \N__23583\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__23583\,
            I => \N__23579\
        );

    \I__2455\ : CascadeMux
    port map (
            O => \N__23582\,
            I => \N__23576\
        );

    \I__2454\ : Span4Mux_s3_h
    port map (
            O => \N__23579\,
            I => \N__23573\
        );

    \I__2453\ : InMux
    port map (
            O => \N__23576\,
            I => \N__23570\
        );

    \I__2452\ : Span4Mux_v
    port map (
            O => \N__23573\,
            I => \N__23567\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__23570\,
            I => n2628
        );

    \I__2450\ : Odrv4
    port map (
            O => \N__23567\,
            I => n2628
        );

    \I__2449\ : CascadeMux
    port map (
            O => \N__23562\,
            I => \N__23559\
        );

    \I__2448\ : InMux
    port map (
            O => \N__23559\,
            I => \N__23556\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__23556\,
            I => \N__23553\
        );

    \I__2446\ : Span4Mux_v
    port map (
            O => \N__23553\,
            I => \N__23548\
        );

    \I__2445\ : InMux
    port map (
            O => \N__23552\,
            I => \N__23543\
        );

    \I__2444\ : InMux
    port map (
            O => \N__23551\,
            I => \N__23543\
        );

    \I__2443\ : Odrv4
    port map (
            O => \N__23548\,
            I => n2727
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__23543\,
            I => n2727
        );

    \I__2441\ : InMux
    port map (
            O => \N__23538\,
            I => \N__23535\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__23535\,
            I => \N__23532\
        );

    \I__2439\ : Span4Mux_v
    port map (
            O => \N__23532\,
            I => \N__23529\
        );

    \I__2438\ : Span4Mux_v
    port map (
            O => \N__23529\,
            I => \N__23526\
        );

    \I__2437\ : Odrv4
    port map (
            O => \N__23526\,
            I => n2700
        );

    \I__2436\ : InMux
    port map (
            O => \N__23523\,
            I => \N__23520\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__23520\,
            I => \N__23517\
        );

    \I__2434\ : Odrv12
    port map (
            O => \N__23517\,
            I => n2288
        );

    \I__2433\ : InMux
    port map (
            O => \N__23514\,
            I => \N__23511\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__23511\,
            I => \N__23508\
        );

    \I__2431\ : Odrv4
    port map (
            O => \N__23508\,
            I => n2391
        );

    \I__2430\ : InMux
    port map (
            O => \N__23505\,
            I => \N__23502\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__23502\,
            I => \N__23499\
        );

    \I__2428\ : Odrv12
    port map (
            O => \N__23499\,
            I => n2287
        );

    \I__2427\ : InMux
    port map (
            O => \N__23496\,
            I => \N__23493\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__23493\,
            I => \N__23490\
        );

    \I__2425\ : Odrv4
    port map (
            O => \N__23490\,
            I => n2386
        );

    \I__2424\ : CascadeMux
    port map (
            O => \N__23487\,
            I => \n2319_cascade_\
        );

    \I__2423\ : InMux
    port map (
            O => \N__23484\,
            I => \N__23481\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__23481\,
            I => \N__23478\
        );

    \I__2421\ : Odrv4
    port map (
            O => \N__23478\,
            I => n11971
        );

    \I__2420\ : InMux
    port map (
            O => \N__23475\,
            I => \N__23472\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__23472\,
            I => \N__23469\
        );

    \I__2418\ : Span4Mux_v
    port map (
            O => \N__23469\,
            I => \N__23466\
        );

    \I__2417\ : Odrv4
    port map (
            O => \N__23466\,
            I => n2292
        );

    \I__2416\ : CascadeMux
    port map (
            O => \N__23463\,
            I => \N__23459\
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__23462\,
            I => \N__23456\
        );

    \I__2414\ : InMux
    port map (
            O => \N__23459\,
            I => \N__23453\
        );

    \I__2413\ : InMux
    port map (
            O => \N__23456\,
            I => \N__23450\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__23453\,
            I => \N__23447\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__23450\,
            I => n2324
        );

    \I__2410\ : Odrv4
    port map (
            O => \N__23447\,
            I => n2324
        );

    \I__2409\ : CascadeMux
    port map (
            O => \N__23442\,
            I => \n2324_cascade_\
        );

    \I__2408\ : InMux
    port map (
            O => \N__23439\,
            I => \N__23436\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__23436\,
            I => \N__23432\
        );

    \I__2406\ : InMux
    port map (
            O => \N__23435\,
            I => \N__23429\
        );

    \I__2405\ : Odrv4
    port map (
            O => \N__23432\,
            I => n2319
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__23429\,
            I => n2319
        );

    \I__2403\ : CascadeMux
    port map (
            O => \N__23424\,
            I => \n14384_cascade_\
        );

    \I__2402\ : InMux
    port map (
            O => \N__23421\,
            I => \N__23418\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__23418\,
            I => \N__23415\
        );

    \I__2400\ : Odrv4
    port map (
            O => \N__23415\,
            I => n14382
        );

    \I__2399\ : InMux
    port map (
            O => \N__23412\,
            I => \N__23409\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__23409\,
            I => n14390
        );

    \I__2397\ : InMux
    port map (
            O => \N__23406\,
            I => \N__23403\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__23403\,
            I => \N__23400\
        );

    \I__2395\ : Odrv12
    port map (
            O => \N__23400\,
            I => n2293
        );

    \I__2394\ : InMux
    port map (
            O => \N__23397\,
            I => \N__23394\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__23394\,
            I => \N__23391\
        );

    \I__2392\ : Odrv12
    port map (
            O => \N__23391\,
            I => n2298
        );

    \I__2391\ : InMux
    port map (
            O => \N__23388\,
            I => \N__23385\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__23385\,
            I => \N__23382\
        );

    \I__2389\ : Odrv12
    port map (
            O => \N__23382\,
            I => n2295
        );

    \I__2388\ : InMux
    port map (
            O => \N__23379\,
            I => \N__23376\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__23376\,
            I => \N__23373\
        );

    \I__2386\ : Odrv12
    port map (
            O => \N__23373\,
            I => n2296
        );

    \I__2385\ : InMux
    port map (
            O => \N__23370\,
            I => \N__23367\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__23367\,
            I => \N__23364\
        );

    \I__2383\ : Odrv4
    port map (
            O => \N__23364\,
            I => n11977
        );

    \I__2382\ : CascadeMux
    port map (
            O => \N__23361\,
            I => \n14808_cascade_\
        );

    \I__2381\ : InMux
    port map (
            O => \N__23358\,
            I => \N__23355\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__23355\,
            I => \N__23352\
        );

    \I__2379\ : Odrv4
    port map (
            O => \N__23352\,
            I => n14594
        );

    \I__2378\ : CascadeMux
    port map (
            O => \N__23349\,
            I => \N__23346\
        );

    \I__2377\ : InMux
    port map (
            O => \N__23346\,
            I => \N__23343\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__23343\,
            I => \N__23339\
        );

    \I__2375\ : InMux
    port map (
            O => \N__23342\,
            I => \N__23336\
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__23339\,
            I => n2219
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__23336\,
            I => n2219
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__23331\,
            I => \n14598_cascade_\
        );

    \I__2371\ : CascadeMux
    port map (
            O => \N__23328\,
            I => \n14604_cascade_\
        );

    \I__2370\ : CascadeMux
    port map (
            O => \N__23325\,
            I => \n2247_cascade_\
        );

    \I__2369\ : InMux
    port map (
            O => \N__23322\,
            I => \N__23319\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__23319\,
            I => \N__23316\
        );

    \I__2367\ : Span4Mux_v
    port map (
            O => \N__23316\,
            I => \N__23313\
        );

    \I__2366\ : Odrv4
    port map (
            O => \N__23313\,
            I => n2297
        );

    \I__2365\ : CascadeMux
    port map (
            O => \N__23310\,
            I => \N__23307\
        );

    \I__2364\ : InMux
    port map (
            O => \N__23307\,
            I => \N__23304\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__23304\,
            I => \N__23300\
        );

    \I__2362\ : InMux
    port map (
            O => \N__23303\,
            I => \N__23297\
        );

    \I__2361\ : Odrv4
    port map (
            O => \N__23300\,
            I => n2222
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__23297\,
            I => n2222
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__23292\,
            I => \n2222_cascade_\
        );

    \I__2358\ : InMux
    port map (
            O => \N__23289\,
            I => \N__23286\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__23286\,
            I => \N__23283\
        );

    \I__2356\ : Odrv4
    port map (
            O => \N__23283\,
            I => n2289
        );

    \I__2355\ : InMux
    port map (
            O => \N__23280\,
            I => \N__23277\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__23277\,
            I => \N__23274\
        );

    \I__2353\ : Odrv4
    port map (
            O => \N__23274\,
            I => n2291
        );

    \I__2352\ : CascadeMux
    port map (
            O => \N__23271\,
            I => \n2323_cascade_\
        );

    \I__2351\ : CascadeMux
    port map (
            O => \N__23268\,
            I => \n2219_cascade_\
        );

    \I__2350\ : InMux
    port map (
            O => \N__23265\,
            I => \N__23262\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__23262\,
            I => \N__23259\
        );

    \I__2348\ : Odrv12
    port map (
            O => \N__23259\,
            I => n2286
        );

    \I__2347\ : InMux
    port map (
            O => \N__23256\,
            I => \N__23253\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__23253\,
            I => \N__23250\
        );

    \I__2345\ : Odrv4
    port map (
            O => \N__23250\,
            I => n2290
        );

    \I__2344\ : InMux
    port map (
            O => \N__23247\,
            I => n12693
        );

    \I__2343\ : InMux
    port map (
            O => \N__23244\,
            I => n12694
        );

    \I__2342\ : InMux
    port map (
            O => \N__23241\,
            I => n12695
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__23238\,
            I => \N__23235\
        );

    \I__2340\ : InMux
    port map (
            O => \N__23235\,
            I => \N__23231\
        );

    \I__2339\ : CascadeMux
    port map (
            O => \N__23234\,
            I => \N__23228\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__23231\,
            I => \N__23225\
        );

    \I__2337\ : InMux
    port map (
            O => \N__23228\,
            I => \N__23222\
        );

    \I__2336\ : Odrv4
    port map (
            O => \N__23225\,
            I => n2233
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__23222\,
            I => n2233
        );

    \I__2334\ : InMux
    port map (
            O => \N__23217\,
            I => \N__23214\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__23214\,
            I => \N__23211\
        );

    \I__2332\ : Odrv12
    port map (
            O => \N__23211\,
            I => n2300
        );

    \I__2331\ : CascadeMux
    port map (
            O => \N__23208\,
            I => \n2233_cascade_\
        );

    \I__2330\ : InMux
    port map (
            O => \N__23205\,
            I => \N__23202\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__23202\,
            I => \N__23199\
        );

    \I__2328\ : Odrv4
    port map (
            O => \N__23199\,
            I => n2299
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__23196\,
            I => \n2331_cascade_\
        );

    \I__2326\ : InMux
    port map (
            O => \N__23193\,
            I => \N__23190\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__23190\,
            I => \N__23187\
        );

    \I__2324\ : Odrv12
    port map (
            O => \N__23187\,
            I => n2301
        );

    \I__2323\ : InMux
    port map (
            O => \N__23184\,
            I => n12684
        );

    \I__2322\ : InMux
    port map (
            O => \N__23181\,
            I => n12685
        );

    \I__2321\ : InMux
    port map (
            O => \N__23178\,
            I => n12686
        );

    \I__2320\ : InMux
    port map (
            O => \N__23175\,
            I => n12687
        );

    \I__2319\ : InMux
    port map (
            O => \N__23172\,
            I => n12688
        );

    \I__2318\ : InMux
    port map (
            O => \N__23169\,
            I => n12689
        );

    \I__2317\ : InMux
    port map (
            O => \N__23166\,
            I => n12690
        );

    \I__2316\ : InMux
    port map (
            O => \N__23163\,
            I => \bfn_3_16_0_\
        );

    \I__2315\ : InMux
    port map (
            O => \N__23160\,
            I => n12692
        );

    \I__2314\ : InMux
    port map (
            O => \N__23157\,
            I => \bfn_3_14_0_\
        );

    \I__2313\ : InMux
    port map (
            O => \N__23154\,
            I => n12676
        );

    \I__2312\ : InMux
    port map (
            O => \N__23151\,
            I => n12677
        );

    \I__2311\ : InMux
    port map (
            O => \N__23148\,
            I => n12678
        );

    \I__2310\ : InMux
    port map (
            O => \N__23145\,
            I => n12679
        );

    \I__2309\ : InMux
    port map (
            O => \N__23142\,
            I => n12680
        );

    \I__2308\ : InMux
    port map (
            O => \N__23139\,
            I => n12681
        );

    \I__2307\ : InMux
    port map (
            O => \N__23136\,
            I => n12682
        );

    \I__2306\ : InMux
    port map (
            O => \N__23133\,
            I => \bfn_3_15_0_\
        );

    \I__2305\ : InMux
    port map (
            O => \N__23130\,
            I => n12912
        );

    \I__2304\ : InMux
    port map (
            O => \N__23127\,
            I => n12913
        );

    \I__2303\ : InMux
    port map (
            O => \N__23124\,
            I => n12914
        );

    \I__2302\ : InMux
    port map (
            O => \N__23121\,
            I => \bfn_2_32_0_\
        );

    \I__2301\ : InMux
    port map (
            O => \N__23118\,
            I => n12916
        );

    \I__2300\ : InMux
    port map (
            O => \N__23115\,
            I => n12917
        );

    \I__2299\ : InMux
    port map (
            O => \N__23112\,
            I => n12918
        );

    \I__2298\ : InMux
    port map (
            O => \N__23109\,
            I => n12919
        );

    \I__2297\ : InMux
    port map (
            O => \N__23106\,
            I => n12920
        );

    \I__2296\ : InMux
    port map (
            O => \N__23103\,
            I => n12903
        );

    \I__2295\ : InMux
    port map (
            O => \N__23100\,
            I => n12904
        );

    \I__2294\ : InMux
    port map (
            O => \N__23097\,
            I => \N__23093\
        );

    \I__2293\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23090\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__23093\,
            I => n3120
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__23090\,
            I => n3120
        );

    \I__2290\ : InMux
    port map (
            O => \N__23085\,
            I => \N__23082\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__23082\,
            I => n3187
        );

    \I__2288\ : InMux
    port map (
            O => \N__23079\,
            I => n12905
        );

    \I__2287\ : InMux
    port map (
            O => \N__23076\,
            I => n12906
        );

    \I__2286\ : InMux
    port map (
            O => \N__23073\,
            I => \bfn_2_31_0_\
        );

    \I__2285\ : InMux
    port map (
            O => \N__23070\,
            I => n12908
        );

    \I__2284\ : InMux
    port map (
            O => \N__23067\,
            I => n12909
        );

    \I__2283\ : InMux
    port map (
            O => \N__23064\,
            I => n12910
        );

    \I__2282\ : InMux
    port map (
            O => \N__23061\,
            I => n12911
        );

    \I__2281\ : InMux
    port map (
            O => \N__23058\,
            I => n12894
        );

    \I__2280\ : InMux
    port map (
            O => \N__23055\,
            I => n12895
        );

    \I__2279\ : InMux
    port map (
            O => \N__23052\,
            I => n12896
        );

    \I__2278\ : InMux
    port map (
            O => \N__23049\,
            I => n12897
        );

    \I__2277\ : InMux
    port map (
            O => \N__23046\,
            I => n12898
        );

    \I__2276\ : InMux
    port map (
            O => \N__23043\,
            I => \bfn_2_30_0_\
        );

    \I__2275\ : InMux
    port map (
            O => \N__23040\,
            I => n12900
        );

    \I__2274\ : InMux
    port map (
            O => \N__23037\,
            I => n12901
        );

    \I__2273\ : InMux
    port map (
            O => \N__23034\,
            I => n12902
        );

    \I__2272\ : InMux
    port map (
            O => \N__23031\,
            I => n12861
        );

    \I__2271\ : InMux
    port map (
            O => \N__23028\,
            I => \N__23025\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__23025\,
            I => \N__23022\
        );

    \I__2269\ : Odrv4
    port map (
            O => \N__23022\,
            I => n2975
        );

    \I__2268\ : InMux
    port map (
            O => \N__23019\,
            I => n12862
        );

    \I__2267\ : InMux
    port map (
            O => \N__23016\,
            I => n12863
        );

    \I__2266\ : InMux
    port map (
            O => \N__23013\,
            I => \bfn_2_29_0_\
        );

    \I__2265\ : InMux
    port map (
            O => \N__23010\,
            I => n12892
        );

    \I__2264\ : InMux
    port map (
            O => \N__23007\,
            I => n12893
        );

    \I__2263\ : InMux
    port map (
            O => \N__23004\,
            I => \N__23001\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__23001\,
            I => n2985
        );

    \I__2261\ : InMux
    port map (
            O => \N__22998\,
            I => \bfn_2_27_0_\
        );

    \I__2260\ : InMux
    port map (
            O => \N__22995\,
            I => n12853
        );

    \I__2259\ : InMux
    port map (
            O => \N__22992\,
            I => n12854
        );

    \I__2258\ : InMux
    port map (
            O => \N__22989\,
            I => n12855
        );

    \I__2257\ : InMux
    port map (
            O => \N__22986\,
            I => n12856
        );

    \I__2256\ : InMux
    port map (
            O => \N__22983\,
            I => n12857
        );

    \I__2255\ : InMux
    port map (
            O => \N__22980\,
            I => n12858
        );

    \I__2254\ : InMux
    port map (
            O => \N__22977\,
            I => n12859
        );

    \I__2253\ : CascadeMux
    port map (
            O => \N__22974\,
            I => \N__22971\
        );

    \I__2252\ : InMux
    port map (
            O => \N__22971\,
            I => \N__22968\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__22968\,
            I => n2977
        );

    \I__2250\ : InMux
    port map (
            O => \N__22965\,
            I => \bfn_2_28_0_\
        );

    \I__2249\ : InMux
    port map (
            O => \N__22962\,
            I => \N__22959\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__22959\,
            I => n2993
        );

    \I__2247\ : InMux
    port map (
            O => \N__22956\,
            I => \bfn_2_26_0_\
        );

    \I__2246\ : InMux
    port map (
            O => \N__22953\,
            I => \N__22950\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__22950\,
            I => n2992
        );

    \I__2244\ : InMux
    port map (
            O => \N__22947\,
            I => n12845
        );

    \I__2243\ : InMux
    port map (
            O => \N__22944\,
            I => n12846
        );

    \I__2242\ : CascadeMux
    port map (
            O => \N__22941\,
            I => \N__22938\
        );

    \I__2241\ : InMux
    port map (
            O => \N__22938\,
            I => \N__22935\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__22935\,
            I => n2990
        );

    \I__2239\ : InMux
    port map (
            O => \N__22932\,
            I => n12847
        );

    \I__2238\ : InMux
    port map (
            O => \N__22929\,
            I => \N__22926\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__22926\,
            I => n2989
        );

    \I__2236\ : InMux
    port map (
            O => \N__22923\,
            I => n12848
        );

    \I__2235\ : InMux
    port map (
            O => \N__22920\,
            I => n12849
        );

    \I__2234\ : InMux
    port map (
            O => \N__22917\,
            I => n12850
        );

    \I__2233\ : InMux
    port map (
            O => \N__22914\,
            I => n12851
        );

    \I__2232\ : InMux
    port map (
            O => \N__22911\,
            I => \N__22908\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__22908\,
            I => \N__22905\
        );

    \I__2230\ : Odrv12
    port map (
            O => \N__22905\,
            I => n2791
        );

    \I__2229\ : InMux
    port map (
            O => \N__22902\,
            I => \bfn_2_25_0_\
        );

    \I__2228\ : InMux
    port map (
            O => \N__22899\,
            I => n12837
        );

    \I__2227\ : InMux
    port map (
            O => \N__22896\,
            I => n12838
        );

    \I__2226\ : InMux
    port map (
            O => \N__22893\,
            I => n12839
        );

    \I__2225\ : InMux
    port map (
            O => \N__22890\,
            I => n12840
        );

    \I__2224\ : InMux
    port map (
            O => \N__22887\,
            I => n12841
        );

    \I__2223\ : InMux
    port map (
            O => \N__22884\,
            I => n12842
        );

    \I__2222\ : InMux
    port map (
            O => \N__22881\,
            I => \N__22878\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__22878\,
            I => n2994
        );

    \I__2220\ : InMux
    port map (
            O => \N__22875\,
            I => n12843
        );

    \I__2219\ : InMux
    port map (
            O => \N__22872\,
            I => \N__22869\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__22869\,
            I => \N__22866\
        );

    \I__2217\ : Span4Mux_v
    port map (
            O => \N__22866\,
            I => \N__22863\
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__22863\,
            I => n2785
        );

    \I__2215\ : InMux
    port map (
            O => \N__22860\,
            I => \N__22857\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__22857\,
            I => \N__22854\
        );

    \I__2213\ : Span4Mux_v
    port map (
            O => \N__22854\,
            I => \N__22851\
        );

    \I__2212\ : Span4Mux_v
    port map (
            O => \N__22851\,
            I => \N__22848\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__22848\,
            I => n2684
        );

    \I__2210\ : InMux
    port map (
            O => \N__22845\,
            I => \N__22840\
        );

    \I__2209\ : InMux
    port map (
            O => \N__22844\,
            I => \N__22837\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__22843\,
            I => \N__22834\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__22840\,
            I => \N__22831\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__22837\,
            I => \N__22828\
        );

    \I__2205\ : InMux
    port map (
            O => \N__22834\,
            I => \N__22825\
        );

    \I__2204\ : Odrv4
    port map (
            O => \N__22831\,
            I => n2716
        );

    \I__2203\ : Odrv12
    port map (
            O => \N__22828\,
            I => n2716
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__22825\,
            I => n2716
        );

    \I__2201\ : CascadeMux
    port map (
            O => \N__22818\,
            I => \N__22815\
        );

    \I__2200\ : InMux
    port map (
            O => \N__22815\,
            I => \N__22812\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__22812\,
            I => \N__22809\
        );

    \I__2198\ : Span4Mux_v
    port map (
            O => \N__22809\,
            I => \N__22806\
        );

    \I__2197\ : Span4Mux_v
    port map (
            O => \N__22806\,
            I => \N__22803\
        );

    \I__2196\ : Odrv4
    port map (
            O => \N__22803\,
            I => n2679
        );

    \I__2195\ : InMux
    port map (
            O => \N__22800\,
            I => \N__22796\
        );

    \I__2194\ : InMux
    port map (
            O => \N__22799\,
            I => \N__22793\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__22796\,
            I => \N__22790\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__22793\,
            I => n2709
        );

    \I__2191\ : Odrv12
    port map (
            O => \N__22790\,
            I => n2709
        );

    \I__2190\ : CascadeMux
    port map (
            O => \N__22785\,
            I => \n2711_cascade_\
        );

    \I__2189\ : InMux
    port map (
            O => \N__22782\,
            I => \N__22779\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__22779\,
            I => n14368
        );

    \I__2187\ : InMux
    port map (
            O => \N__22776\,
            I => \N__22773\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__22773\,
            I => \N__22770\
        );

    \I__2185\ : Span4Mux_v
    port map (
            O => \N__22770\,
            I => \N__22767\
        );

    \I__2184\ : Odrv4
    port map (
            O => \N__22767\,
            I => n2796
        );

    \I__2183\ : CascadeMux
    port map (
            O => \N__22764\,
            I => \n2742_cascade_\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__22761\,
            I => \N__22758\
        );

    \I__2181\ : InMux
    port map (
            O => \N__22758\,
            I => \N__22753\
        );

    \I__2180\ : InMux
    port map (
            O => \N__22757\,
            I => \N__22750\
        );

    \I__2179\ : InMux
    port map (
            O => \N__22756\,
            I => \N__22747\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__22753\,
            I => \N__22744\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__22750\,
            I => \N__22741\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__22747\,
            I => \N__22738\
        );

    \I__2175\ : Odrv4
    port map (
            O => \N__22744\,
            I => n2828
        );

    \I__2174\ : Odrv4
    port map (
            O => \N__22741\,
            I => n2828
        );

    \I__2173\ : Odrv4
    port map (
            O => \N__22738\,
            I => n2828
        );

    \I__2172\ : InMux
    port map (
            O => \N__22731\,
            I => \N__22728\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__22728\,
            I => \N__22725\
        );

    \I__2170\ : Span4Mux_v
    port map (
            O => \N__22725\,
            I => \N__22722\
        );

    \I__2169\ : Odrv4
    port map (
            O => \N__22722\,
            I => n2788
        );

    \I__2168\ : InMux
    port map (
            O => \N__22719\,
            I => \N__22716\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__22716\,
            I => \N__22713\
        );

    \I__2166\ : Span12Mux_v
    port map (
            O => \N__22713\,
            I => \N__22710\
        );

    \I__2165\ : Odrv12
    port map (
            O => \N__22710\,
            I => n2687
        );

    \I__2164\ : InMux
    port map (
            O => \N__22707\,
            I => \N__22704\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__22704\,
            I => \N__22701\
        );

    \I__2162\ : Odrv12
    port map (
            O => \N__22701\,
            I => n2792
        );

    \I__2161\ : CascadeMux
    port map (
            O => \N__22698\,
            I => \N__22695\
        );

    \I__2160\ : InMux
    port map (
            O => \N__22695\,
            I => \N__22691\
        );

    \I__2159\ : InMux
    port map (
            O => \N__22694\,
            I => \N__22687\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__22691\,
            I => \N__22684\
        );

    \I__2157\ : CascadeMux
    port map (
            O => \N__22690\,
            I => \N__22681\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__22687\,
            I => \N__22678\
        );

    \I__2155\ : Span4Mux_s2_h
    port map (
            O => \N__22684\,
            I => \N__22675\
        );

    \I__2154\ : InMux
    port map (
            O => \N__22681\,
            I => \N__22672\
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__22678\,
            I => n2725
        );

    \I__2152\ : Odrv4
    port map (
            O => \N__22675\,
            I => n2725
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__22672\,
            I => n2725
        );

    \I__2150\ : CascadeMux
    port map (
            O => \N__22665\,
            I => \N__22662\
        );

    \I__2149\ : InMux
    port map (
            O => \N__22662\,
            I => \N__22659\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__22659\,
            I => \N__22656\
        );

    \I__2147\ : Span4Mux_v
    port map (
            O => \N__22656\,
            I => \N__22653\
        );

    \I__2146\ : Odrv4
    port map (
            O => \N__22653\,
            I => n2681
        );

    \I__2145\ : CascadeMux
    port map (
            O => \N__22650\,
            I => \N__22647\
        );

    \I__2144\ : InMux
    port map (
            O => \N__22647\,
            I => \N__22644\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__22644\,
            I => \N__22641\
        );

    \I__2142\ : Span4Mux_v
    port map (
            O => \N__22641\,
            I => \N__22638\
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__22638\,
            I => n2794
        );

    \I__2140\ : CascadeMux
    port map (
            O => \N__22635\,
            I => \n2826_cascade_\
        );

    \I__2139\ : CascadeMux
    port map (
            O => \N__22632\,
            I => \n14362_cascade_\
        );

    \I__2138\ : InMux
    port map (
            O => \N__22629\,
            I => \N__22626\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__22626\,
            I => \N__22623\
        );

    \I__2136\ : Span4Mux_v
    port map (
            O => \N__22623\,
            I => \N__22620\
        );

    \I__2135\ : Odrv4
    port map (
            O => \N__22620\,
            I => n2789
        );

    \I__2134\ : CascadeMux
    port map (
            O => \N__22617\,
            I => \N__22614\
        );

    \I__2133\ : InMux
    port map (
            O => \N__22614\,
            I => \N__22611\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__22611\,
            I => n14346
        );

    \I__2131\ : CascadeMux
    port map (
            O => \N__22608\,
            I => \n14350_cascade_\
        );

    \I__2130\ : InMux
    port map (
            O => \N__22605\,
            I => \N__22602\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__22602\,
            I => n14356
        );

    \I__2128\ : InMux
    port map (
            O => \N__22599\,
            I => \N__22596\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__22596\,
            I => \N__22593\
        );

    \I__2126\ : Span4Mux_v
    port map (
            O => \N__22593\,
            I => \N__22590\
        );

    \I__2125\ : Odrv4
    port map (
            O => \N__22590\,
            I => n2782
        );

    \I__2124\ : CascadeMux
    port map (
            O => \N__22587\,
            I => \N__22584\
        );

    \I__2123\ : InMux
    port map (
            O => \N__22584\,
            I => \N__22577\
        );

    \I__2122\ : InMux
    port map (
            O => \N__22583\,
            I => \N__22577\
        );

    \I__2121\ : InMux
    port map (
            O => \N__22582\,
            I => \N__22574\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__22577\,
            I => \N__22571\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__22574\,
            I => n2715
        );

    \I__2118\ : Odrv4
    port map (
            O => \N__22571\,
            I => n2715
        );

    \I__2117\ : CascadeMux
    port map (
            O => \N__22566\,
            I => \n2621_cascade_\
        );

    \I__2116\ : InMux
    port map (
            O => \N__22563\,
            I => \N__22560\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__22560\,
            I => \N__22557\
        );

    \I__2114\ : Span4Mux_v
    port map (
            O => \N__22557\,
            I => \N__22554\
        );

    \I__2113\ : Odrv4
    port map (
            O => \N__22554\,
            I => n2688
        );

    \I__2112\ : InMux
    port map (
            O => \N__22551\,
            I => \N__22548\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__22548\,
            I => \N__22545\
        );

    \I__2110\ : Span4Mux_v
    port map (
            O => \N__22545\,
            I => \N__22542\
        );

    \I__2109\ : Span4Mux_v
    port map (
            O => \N__22542\,
            I => \N__22539\
        );

    \I__2108\ : Odrv4
    port map (
            O => \N__22539\,
            I => n2696
        );

    \I__2107\ : InMux
    port map (
            O => \N__22536\,
            I => \N__22533\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__22533\,
            I => \N__22530\
        );

    \I__2105\ : Odrv12
    port map (
            O => \N__22530\,
            I => n2795
        );

    \I__2104\ : CascadeMux
    port map (
            O => \N__22527\,
            I => \n2728_cascade_\
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__22524\,
            I => \N__22521\
        );

    \I__2102\ : InMux
    port map (
            O => \N__22521\,
            I => \N__22518\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__22518\,
            I => \N__22515\
        );

    \I__2100\ : Odrv12
    port map (
            O => \N__22515\,
            I => n2691
        );

    \I__2099\ : CascadeMux
    port map (
            O => \N__22512\,
            I => \N__22509\
        );

    \I__2098\ : InMux
    port map (
            O => \N__22509\,
            I => \N__22506\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__22506\,
            I => \N__22503\
        );

    \I__2096\ : Span4Mux_s2_h
    port map (
            O => \N__22503\,
            I => \N__22499\
        );

    \I__2095\ : InMux
    port map (
            O => \N__22502\,
            I => \N__22496\
        );

    \I__2094\ : Odrv4
    port map (
            O => \N__22499\,
            I => n2723
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__22496\,
            I => n2723
        );

    \I__2092\ : InMux
    port map (
            O => \N__22491\,
            I => \N__22488\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__22488\,
            I => \N__22485\
        );

    \I__2090\ : Span4Mux_v
    port map (
            O => \N__22485\,
            I => \N__22482\
        );

    \I__2089\ : Odrv4
    port map (
            O => \N__22482\,
            I => n2790
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__22479\,
            I => \n2723_cascade_\
        );

    \I__2087\ : InMux
    port map (
            O => \N__22476\,
            I => \N__22473\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__22473\,
            I => \N__22470\
        );

    \I__2085\ : Odrv12
    port map (
            O => \N__22470\,
            I => n2693
        );

    \I__2084\ : InMux
    port map (
            O => \N__22467\,
            I => \N__22464\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__22464\,
            I => \N__22461\
        );

    \I__2082\ : Span4Mux_v
    port map (
            O => \N__22461\,
            I => \N__22458\
        );

    \I__2081\ : Span4Mux_v
    port map (
            O => \N__22458\,
            I => \N__22455\
        );

    \I__2080\ : Odrv4
    port map (
            O => \N__22455\,
            I => n2697
        );

    \I__2079\ : InMux
    port map (
            O => \N__22452\,
            I => \bfn_2_20_0_\
        );

    \I__2078\ : InMux
    port map (
            O => \N__22449\,
            I => n12810
        );

    \I__2077\ : InMux
    port map (
            O => \N__22446\,
            I => \N__22443\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__22443\,
            I => \N__22440\
        );

    \I__2075\ : Odrv12
    port map (
            O => \N__22440\,
            I => n2683
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__22437\,
            I => \N__22434\
        );

    \I__2073\ : InMux
    port map (
            O => \N__22434\,
            I => \N__22431\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__22431\,
            I => \N__22428\
        );

    \I__2071\ : Span4Mux_v
    port map (
            O => \N__22428\,
            I => \N__22425\
        );

    \I__2070\ : Odrv4
    port map (
            O => \N__22425\,
            I => n2677
        );

    \I__2069\ : InMux
    port map (
            O => \N__22422\,
            I => \N__22419\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__22419\,
            I => \N__22416\
        );

    \I__2067\ : Odrv12
    port map (
            O => \N__22416\,
            I => n2678
        );

    \I__2066\ : InMux
    port map (
            O => \N__22413\,
            I => \N__22410\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__22410\,
            I => \N__22407\
        );

    \I__2064\ : Odrv12
    port map (
            O => \N__22407\,
            I => n2797
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__22404\,
            I => \N__22401\
        );

    \I__2062\ : InMux
    port map (
            O => \N__22401\,
            I => \N__22398\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__22398\,
            I => \N__22395\
        );

    \I__2060\ : Sp12to4
    port map (
            O => \N__22395\,
            I => \N__22392\
        );

    \I__2059\ : Odrv12
    port map (
            O => \N__22392\,
            I => n2694
        );

    \I__2058\ : InMux
    port map (
            O => \N__22389\,
            I => \N__22386\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__22386\,
            I => \N__22383\
        );

    \I__2056\ : Span4Mux_v
    port map (
            O => \N__22383\,
            I => \N__22380\
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__22380\,
            I => n2793
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__22377\,
            I => \n2726_cascade_\
        );

    \I__2053\ : InMux
    port map (
            O => \N__22374\,
            I => n12800
        );

    \I__2052\ : InMux
    port map (
            O => \N__22371\,
            I => \bfn_2_19_0_\
        );

    \I__2051\ : InMux
    port map (
            O => \N__22368\,
            I => n12802
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__22365\,
            I => \N__22362\
        );

    \I__2049\ : InMux
    port map (
            O => \N__22362\,
            I => \N__22359\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__22359\,
            I => \N__22356\
        );

    \I__2047\ : Sp12to4
    port map (
            O => \N__22356\,
            I => \N__22353\
        );

    \I__2046\ : Odrv12
    port map (
            O => \N__22353\,
            I => n2783
        );

    \I__2045\ : InMux
    port map (
            O => \N__22350\,
            I => n12803
        );

    \I__2044\ : InMux
    port map (
            O => \N__22347\,
            I => n12804
        );

    \I__2043\ : InMux
    port map (
            O => \N__22344\,
            I => n12805
        );

    \I__2042\ : InMux
    port map (
            O => \N__22341\,
            I => n12806
        );

    \I__2041\ : InMux
    port map (
            O => \N__22338\,
            I => n12807
        );

    \I__2040\ : InMux
    port map (
            O => \N__22335\,
            I => n12808
        );

    \I__2039\ : InMux
    port map (
            O => \N__22332\,
            I => n12791
        );

    \I__2038\ : InMux
    port map (
            O => \N__22329\,
            I => n12792
        );

    \I__2037\ : InMux
    port map (
            O => \N__22326\,
            I => \bfn_2_18_0_\
        );

    \I__2036\ : InMux
    port map (
            O => \N__22323\,
            I => n12794
        );

    \I__2035\ : InMux
    port map (
            O => \N__22320\,
            I => n12795
        );

    \I__2034\ : InMux
    port map (
            O => \N__22317\,
            I => n12796
        );

    \I__2033\ : InMux
    port map (
            O => \N__22314\,
            I => n12797
        );

    \I__2032\ : InMux
    port map (
            O => \N__22311\,
            I => n12798
        );

    \I__2031\ : InMux
    port map (
            O => \N__22308\,
            I => n12799
        );

    \I__2030\ : InMux
    port map (
            O => \N__22305\,
            I => n12783
        );

    \I__2029\ : InMux
    port map (
            O => \N__22302\,
            I => n12784
        );

    \I__2028\ : InMux
    port map (
            O => \N__22299\,
            I => \bfn_2_16_0_\
        );

    \I__2027\ : InMux
    port map (
            O => \N__22296\,
            I => \N__22293\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__22293\,
            I => \N__22290\
        );

    \I__2025\ : Span4Mux_v
    port map (
            O => \N__22290\,
            I => \N__22287\
        );

    \I__2024\ : Span4Mux_v
    port map (
            O => \N__22287\,
            I => \N__22284\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__22284\,
            I => n2801
        );

    \I__2022\ : InMux
    port map (
            O => \N__22281\,
            I => \bfn_2_17_0_\
        );

    \I__2021\ : InMux
    port map (
            O => \N__22278\,
            I => n12786
        );

    \I__2020\ : InMux
    port map (
            O => \N__22275\,
            I => n12787
        );

    \I__2019\ : InMux
    port map (
            O => \N__22272\,
            I => n12788
        );

    \I__2018\ : InMux
    port map (
            O => \N__22269\,
            I => n12789
        );

    \I__2017\ : InMux
    port map (
            O => \N__22266\,
            I => n12790
        );

    \I__2016\ : InMux
    port map (
            O => \N__22263\,
            I => n12774
        );

    \I__2015\ : InMux
    port map (
            O => \N__22260\,
            I => n12775
        );

    \I__2014\ : InMux
    port map (
            O => \N__22257\,
            I => n12776
        );

    \I__2013\ : InMux
    port map (
            O => \N__22254\,
            I => \bfn_2_15_0_\
        );

    \I__2012\ : InMux
    port map (
            O => \N__22251\,
            I => n12778
        );

    \I__2011\ : InMux
    port map (
            O => \N__22248\,
            I => n12779
        );

    \I__2010\ : InMux
    port map (
            O => \N__22245\,
            I => \N__22242\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__22242\,
            I => \N__22239\
        );

    \I__2008\ : Sp12to4
    port map (
            O => \N__22239\,
            I => \N__22236\
        );

    \I__2007\ : Odrv12
    port map (
            O => \N__22236\,
            I => n2682
        );

    \I__2006\ : InMux
    port map (
            O => \N__22233\,
            I => n12780
        );

    \I__2005\ : InMux
    port map (
            O => \N__22230\,
            I => n12781
        );

    \I__2004\ : InMux
    port map (
            O => \N__22227\,
            I => n12782
        );

    \I__2003\ : InMux
    port map (
            O => \N__22224\,
            I => n12764
        );

    \I__2002\ : InMux
    port map (
            O => \N__22221\,
            I => n12765
        );

    \I__2001\ : InMux
    port map (
            O => \N__22218\,
            I => n12766
        );

    \I__2000\ : InMux
    port map (
            O => \N__22215\,
            I => n12767
        );

    \I__1999\ : InMux
    port map (
            O => \N__22212\,
            I => n12768
        );

    \I__1998\ : InMux
    port map (
            O => \N__22209\,
            I => \bfn_2_14_0_\
        );

    \I__1997\ : InMux
    port map (
            O => \N__22206\,
            I => n12770
        );

    \I__1996\ : InMux
    port map (
            O => \N__22203\,
            I => n12771
        );

    \I__1995\ : InMux
    port map (
            O => \N__22200\,
            I => n12772
        );

    \I__1994\ : InMux
    port map (
            O => \N__22197\,
            I => n12773
        );

    \I__1993\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22190\
        );

    \I__1992\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22187\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__22190\,
            I => \debounce.cnt_reg_5\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__22187\,
            I => \debounce.cnt_reg_5\
        );

    \I__1989\ : InMux
    port map (
            O => \N__22182\,
            I => \debounce.n13017\
        );

    \I__1988\ : InMux
    port map (
            O => \N__22179\,
            I => \N__22175\
        );

    \I__1987\ : InMux
    port map (
            O => \N__22178\,
            I => \N__22172\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__22175\,
            I => \debounce.cnt_reg_6\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__22172\,
            I => \debounce.cnt_reg_6\
        );

    \I__1984\ : InMux
    port map (
            O => \N__22167\,
            I => \debounce.n13018\
        );

    \I__1983\ : InMux
    port map (
            O => \N__22164\,
            I => \N__22160\
        );

    \I__1982\ : InMux
    port map (
            O => \N__22163\,
            I => \N__22157\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__22160\,
            I => \debounce.cnt_reg_7\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__22157\,
            I => \debounce.cnt_reg_7\
        );

    \I__1979\ : InMux
    port map (
            O => \N__22152\,
            I => \debounce.n13019\
        );

    \I__1978\ : InMux
    port map (
            O => \N__22149\,
            I => \N__22145\
        );

    \I__1977\ : InMux
    port map (
            O => \N__22148\,
            I => \N__22142\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__22145\,
            I => \N__22139\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__22142\,
            I => \debounce.cnt_reg_8\
        );

    \I__1974\ : Odrv4
    port map (
            O => \N__22139\,
            I => \debounce.cnt_reg_8\
        );

    \I__1973\ : InMux
    port map (
            O => \N__22134\,
            I => \bfn_1_32_0_\
        );

    \I__1972\ : InMux
    port map (
            O => \N__22131\,
            I => \debounce.n13021\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__22128\,
            I => \N__22125\
        );

    \I__1970\ : InMux
    port map (
            O => \N__22125\,
            I => \N__22121\
        );

    \I__1969\ : InMux
    port map (
            O => \N__22124\,
            I => \N__22118\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__22121\,
            I => \N__22115\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__22118\,
            I => \debounce.cnt_reg_9\
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__22115\,
            I => \debounce.cnt_reg_9\
        );

    \I__1965\ : SRMux
    port map (
            O => \N__22110\,
            I => \N__22107\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__22107\,
            I => \N__22103\
        );

    \I__1963\ : SRMux
    port map (
            O => \N__22106\,
            I => \N__22100\
        );

    \I__1962\ : Span4Mux_s1_v
    port map (
            O => \N__22103\,
            I => \N__22097\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__22100\,
            I => \N__22094\
        );

    \I__1960\ : Odrv4
    port map (
            O => \N__22097\,
            I => \debounce.cnt_next_9__N_424\
        );

    \I__1959\ : Odrv12
    port map (
            O => \N__22094\,
            I => \debounce.cnt_next_9__N_424\
        );

    \I__1958\ : InMux
    port map (
            O => \N__22089\,
            I => \bfn_2_13_0_\
        );

    \I__1957\ : InMux
    port map (
            O => \N__22086\,
            I => n12762
        );

    \I__1956\ : InMux
    port map (
            O => \N__22083\,
            I => n12763
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__22080\,
            I => \debounce.n16_cascade_\
        );

    \I__1954\ : InMux
    port map (
            O => \N__22077\,
            I => \N__22074\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__22074\,
            I => \debounce.n17\
        );

    \I__1952\ : InMux
    port map (
            O => \N__22071\,
            I => \N__22065\
        );

    \I__1951\ : InMux
    port map (
            O => \N__22070\,
            I => \N__22065\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__22065\,
            I => \reg_B_2\
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__22062\,
            I => \n14129_cascade_\
        );

    \I__1948\ : InMux
    port map (
            O => \N__22059\,
            I => \N__22055\
        );

    \I__1947\ : InMux
    port map (
            O => \N__22058\,
            I => \N__22052\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__22055\,
            I => \debounce.cnt_reg_0\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__22052\,
            I => \debounce.cnt_reg_0\
        );

    \I__1944\ : InMux
    port map (
            O => \N__22047\,
            I => \bfn_1_31_0_\
        );

    \I__1943\ : InMux
    port map (
            O => \N__22044\,
            I => \N__22040\
        );

    \I__1942\ : InMux
    port map (
            O => \N__22043\,
            I => \N__22037\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__22040\,
            I => \debounce.cnt_reg_1\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__22037\,
            I => \debounce.cnt_reg_1\
        );

    \I__1939\ : InMux
    port map (
            O => \N__22032\,
            I => \debounce.n13013\
        );

    \I__1938\ : CascadeMux
    port map (
            O => \N__22029\,
            I => \N__22025\
        );

    \I__1937\ : InMux
    port map (
            O => \N__22028\,
            I => \N__22022\
        );

    \I__1936\ : InMux
    port map (
            O => \N__22025\,
            I => \N__22019\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__22022\,
            I => \debounce.cnt_reg_2\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__22019\,
            I => \debounce.cnt_reg_2\
        );

    \I__1933\ : InMux
    port map (
            O => \N__22014\,
            I => \debounce.n13014\
        );

    \I__1932\ : InMux
    port map (
            O => \N__22011\,
            I => \N__22007\
        );

    \I__1931\ : InMux
    port map (
            O => \N__22010\,
            I => \N__22004\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__22007\,
            I => \debounce.cnt_reg_3\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__22004\,
            I => \debounce.cnt_reg_3\
        );

    \I__1928\ : InMux
    port map (
            O => \N__21999\,
            I => \debounce.n13015\
        );

    \I__1927\ : InMux
    port map (
            O => \N__21996\,
            I => \N__21992\
        );

    \I__1926\ : InMux
    port map (
            O => \N__21995\,
            I => \N__21989\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__21992\,
            I => \debounce.cnt_reg_4\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__21989\,
            I => \debounce.cnt_reg_4\
        );

    \I__1923\ : InMux
    port map (
            O => \N__21984\,
            I => \debounce.n13016\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__21981\,
            I => \n3120_cascade_\
        );

    \I__1921\ : CascadeMux
    port map (
            O => \N__21978\,
            I => \n3122_cascade_\
        );

    \I__1920\ : InMux
    port map (
            O => \N__21975\,
            I => \N__21972\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__21972\,
            I => n14146
        );

    \I__1918\ : InMux
    port map (
            O => \N__21969\,
            I => \N__21963\
        );

    \I__1917\ : InMux
    port map (
            O => \N__21968\,
            I => \N__21963\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__21963\,
            I => \debounce.reg_A_2\
        );

    \I__1915\ : CascadeMux
    port map (
            O => \N__21960\,
            I => \N__21956\
        );

    \I__1914\ : InMux
    port map (
            O => \N__21959\,
            I => \N__21951\
        );

    \I__1913\ : InMux
    port map (
            O => \N__21956\,
            I => \N__21951\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__21951\,
            I => \N__21948\
        );

    \I__1911\ : IoSpan4Mux
    port map (
            O => \N__21948\,
            I => \N__21945\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__21945\,
            I => \debounce.reg_A_1\
        );

    \I__1909\ : InMux
    port map (
            O => \N__21942\,
            I => \N__21938\
        );

    \I__1908\ : InMux
    port map (
            O => \N__21941\,
            I => \N__21935\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__21938\,
            I => \N__21932\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__21935\,
            I => \N__21929\
        );

    \I__1905\ : Span4Mux_h
    port map (
            O => \N__21932\,
            I => \N__21924\
        );

    \I__1904\ : Span4Mux_v
    port map (
            O => \N__21929\,
            I => \N__21924\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__21924\,
            I => \debounce.reg_A_0\
        );

    \I__1902\ : InMux
    port map (
            O => \N__21921\,
            I => \N__21917\
        );

    \I__1901\ : InMux
    port map (
            O => \N__21920\,
            I => \N__21914\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__21917\,
            I => \N__21911\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__21914\,
            I => \N__21908\
        );

    \I__1898\ : Odrv4
    port map (
            O => \N__21911\,
            I => \reg_B_0\
        );

    \I__1897\ : Odrv12
    port map (
            O => \N__21908\,
            I => \reg_B_0\
        );

    \I__1896\ : CascadeMux
    port map (
            O => \N__21903\,
            I => \debounce.n6_cascade_\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__21900\,
            I => \n3021_cascade_\
        );

    \I__1894\ : InMux
    port map (
            O => \N__21897\,
            I => \N__21894\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__21894\,
            I => n14728
        );

    \I__1892\ : CascadeMux
    port map (
            O => \N__21891\,
            I => \n14150_cascade_\
        );

    \I__1891\ : CascadeMux
    port map (
            O => \N__21888\,
            I => \n3128_cascade_\
        );

    \I__1890\ : InMux
    port map (
            O => \N__21885\,
            I => \N__21882\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__21882\,
            I => n14148
        );

    \I__1888\ : InMux
    port map (
            O => \N__21879\,
            I => \N__21876\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__21876\,
            I => \N__21873\
        );

    \I__1886\ : Span4Mux_v
    port map (
            O => \N__21873\,
            I => \N__21870\
        );

    \I__1885\ : Odrv4
    port map (
            O => \N__21870\,
            I => n2895
        );

    \I__1884\ : CascadeMux
    port map (
            O => \N__21867\,
            I => \n2927_cascade_\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__21864\,
            I => \n3024_cascade_\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__21861\,
            I => \n14730_cascade_\
        );

    \I__1881\ : InMux
    port map (
            O => \N__21858\,
            I => n12835
        );

    \I__1880\ : InMux
    port map (
            O => \N__21855\,
            I => n12836
        );

    \I__1879\ : InMux
    port map (
            O => \N__21852\,
            I => \N__21849\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__21849\,
            I => n2882
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__21846\,
            I => \N__21843\
        );

    \I__1876\ : InMux
    port map (
            O => \N__21843\,
            I => \N__21840\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__21840\,
            I => \N__21837\
        );

    \I__1874\ : Odrv12
    port map (
            O => \N__21837\,
            I => n2900
        );

    \I__1873\ : InMux
    port map (
            O => \N__21834\,
            I => \N__21831\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__21831\,
            I => n2876
        );

    \I__1871\ : CascadeMux
    port map (
            O => \N__21828\,
            I => \n2908_cascade_\
        );

    \I__1870\ : InMux
    port map (
            O => \N__21825\,
            I => \bfn_1_24_0_\
        );

    \I__1869\ : InMux
    port map (
            O => \N__21822\,
            I => n12827
        );

    \I__1868\ : InMux
    port map (
            O => \N__21819\,
            I => n12828
        );

    \I__1867\ : InMux
    port map (
            O => \N__21816\,
            I => n12829
        );

    \I__1866\ : InMux
    port map (
            O => \N__21813\,
            I => n12830
        );

    \I__1865\ : InMux
    port map (
            O => \N__21810\,
            I => n12831
        );

    \I__1864\ : InMux
    port map (
            O => \N__21807\,
            I => n12832
        );

    \I__1863\ : InMux
    port map (
            O => \N__21804\,
            I => n12833
        );

    \I__1862\ : InMux
    port map (
            O => \N__21801\,
            I => \bfn_1_25_0_\
        );

    \I__1861\ : InMux
    port map (
            O => \N__21798\,
            I => n12817
        );

    \I__1860\ : InMux
    port map (
            O => \N__21795\,
            I => \bfn_1_23_0_\
        );

    \I__1859\ : InMux
    port map (
            O => \N__21792\,
            I => n12819
        );

    \I__1858\ : InMux
    port map (
            O => \N__21789\,
            I => n12820
        );

    \I__1857\ : InMux
    port map (
            O => \N__21786\,
            I => n12821
        );

    \I__1856\ : InMux
    port map (
            O => \N__21783\,
            I => n12822
        );

    \I__1855\ : InMux
    port map (
            O => \N__21780\,
            I => n12823
        );

    \I__1854\ : InMux
    port map (
            O => \N__21777\,
            I => n12824
        );

    \I__1853\ : InMux
    port map (
            O => \N__21774\,
            I => n12825
        );

    \I__1852\ : InMux
    port map (
            O => \N__21771\,
            I => n12715
        );

    \I__1851\ : InMux
    port map (
            O => \N__21768\,
            I => n12716
        );

    \I__1850\ : InMux
    port map (
            O => \N__21765\,
            I => \bfn_1_22_0_\
        );

    \I__1849\ : InMux
    port map (
            O => \N__21762\,
            I => n12811
        );

    \I__1848\ : InMux
    port map (
            O => \N__21759\,
            I => n12812
        );

    \I__1847\ : InMux
    port map (
            O => \N__21756\,
            I => n12813
        );

    \I__1846\ : InMux
    port map (
            O => \N__21753\,
            I => n12814
        );

    \I__1845\ : InMux
    port map (
            O => \N__21750\,
            I => n12815
        );

    \I__1844\ : InMux
    port map (
            O => \N__21747\,
            I => n12816
        );

    \I__1843\ : InMux
    port map (
            O => \N__21744\,
            I => n12706
        );

    \I__1842\ : InMux
    port map (
            O => \N__21741\,
            I => n12707
        );

    \I__1841\ : InMux
    port map (
            O => \N__21738\,
            I => n12708
        );

    \I__1840\ : InMux
    port map (
            O => \N__21735\,
            I => n12709
        );

    \I__1839\ : InMux
    port map (
            O => \N__21732\,
            I => n12710
        );

    \I__1838\ : InMux
    port map (
            O => \N__21729\,
            I => \bfn_1_21_0_\
        );

    \I__1837\ : InMux
    port map (
            O => \N__21726\,
            I => n12712
        );

    \I__1836\ : InMux
    port map (
            O => \N__21723\,
            I => n12713
        );

    \I__1835\ : InMux
    port map (
            O => \N__21720\,
            I => n12714
        );

    \I__1834\ : InMux
    port map (
            O => \N__21717\,
            I => n12697
        );

    \I__1833\ : InMux
    port map (
            O => \N__21714\,
            I => n12698
        );

    \I__1832\ : InMux
    port map (
            O => \N__21711\,
            I => n12699
        );

    \I__1831\ : InMux
    port map (
            O => \N__21708\,
            I => n12700
        );

    \I__1830\ : InMux
    port map (
            O => \N__21705\,
            I => n12701
        );

    \I__1829\ : InMux
    port map (
            O => \N__21702\,
            I => n12702
        );

    \I__1828\ : InMux
    port map (
            O => \N__21699\,
            I => \bfn_1_20_0_\
        );

    \I__1827\ : InMux
    port map (
            O => \N__21696\,
            I => n12704
        );

    \I__1826\ : InMux
    port map (
            O => \N__21693\,
            I => n12705
        );

    \I__1825\ : InMux
    port map (
            O => \N__21690\,
            I => \bfn_1_19_0_\
        );

    \I__1824\ : InMux
    port map (
            O => \N__21687\,
            I => n12696
        );

    \I__1823\ : IoInMux
    port map (
            O => \N__21684\,
            I => \N__21681\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__21681\,
            I => \N__21678\
        );

    \I__1821\ : IoSpan4Mux
    port map (
            O => \N__21678\,
            I => \N__21675\
        );

    \I__1820\ : IoSpan4Mux
    port map (
            O => \N__21675\,
            I => \N__21672\
        );

    \I__1819\ : IoSpan4Mux
    port map (
            O => \N__21672\,
            I => \N__21669\
        );

    \I__1818\ : Odrv4
    port map (
            O => \N__21669\,
            I => \CLK_pad_gb_input\
        );

    \IN_MUX_bfv_7_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_29_0_\
        );

    \IN_MUX_bfv_7_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12928,
            carryinitout => \bfn_7_30_0_\
        );

    \IN_MUX_bfv_7_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12936,
            carryinitout => \bfn_7_31_0_\
        );

    \IN_MUX_bfv_7_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12944,
            carryinitout => \bfn_7_32_0_\
        );

    \IN_MUX_bfv_15_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_25_0_\
        );

    \IN_MUX_bfv_15_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12456,
            carryinitout => \bfn_15_26_0_\
        );

    \IN_MUX_bfv_15_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12464,
            carryinitout => \bfn_15_27_0_\
        );

    \IN_MUX_bfv_15_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12472,
            carryinitout => \bfn_15_28_0_\
        );

    \IN_MUX_bfv_11_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_26_0_\
        );

    \IN_MUX_bfv_11_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12433,
            carryinitout => \bfn_11_27_0_\
        );

    \IN_MUX_bfv_11_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12441,
            carryinitout => \bfn_11_28_0_\
        );

    \IN_MUX_bfv_16_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_25_0_\
        );

    \IN_MUX_bfv_16_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n13060,
            carryinitout => \bfn_16_26_0_\
        );

    \IN_MUX_bfv_16_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n13068,
            carryinitout => \bfn_16_27_0_\
        );

    \IN_MUX_bfv_10_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_18_0_\
        );

    \IN_MUX_bfv_10_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n13102\,
            carryinitout => \bfn_10_19_0_\
        );

    \IN_MUX_bfv_10_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n13110\,
            carryinitout => \bfn_10_20_0_\
        );

    \IN_MUX_bfv_10_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \quad_counter0.n13118\,
            carryinitout => \bfn_10_21_0_\
        );

    \IN_MUX_bfv_12_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_25_0_\
        );

    \IN_MUX_bfv_12_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12480,
            carryinitout => \bfn_12_26_0_\
        );

    \IN_MUX_bfv_12_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12488,
            carryinitout => \bfn_12_27_0_\
        );

    \IN_MUX_bfv_9_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_22_0_\
        );

    \IN_MUX_bfv_9_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12982,
            carryinitout => \bfn_9_23_0_\
        );

    \IN_MUX_bfv_9_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12990,
            carryinitout => \bfn_9_24_0_\
        );

    \IN_MUX_bfv_9_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12998,
            carryinitout => \bfn_9_25_0_\
        );

    \IN_MUX_bfv_16_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_17_0_\
        );

    \IN_MUX_bfv_16_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12559,
            carryinitout => \bfn_16_18_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12548,
            carryinitout => \bfn_14_21_0_\
        );

    \IN_MUX_bfv_16_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_21_0_\
        );

    \IN_MUX_bfv_16_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12538,
            carryinitout => \bfn_16_22_0_\
        );

    \IN_MUX_bfv_14_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_23_0_\
        );

    \IN_MUX_bfv_14_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12529,
            carryinitout => \bfn_14_24_0_\
        );

    \IN_MUX_bfv_16_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_23_0_\
        );

    \IN_MUX_bfv_16_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12521,
            carryinitout => \bfn_16_24_0_\
        );

    \IN_MUX_bfv_13_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_24_0_\
        );

    \IN_MUX_bfv_11_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_24_0_\
        );

    \IN_MUX_bfv_2_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_29_0_\
        );

    \IN_MUX_bfv_2_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12899,
            carryinitout => \bfn_2_30_0_\
        );

    \IN_MUX_bfv_2_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12907,
            carryinitout => \bfn_2_31_0_\
        );

    \IN_MUX_bfv_2_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12915,
            carryinitout => \bfn_2_32_0_\
        );

    \IN_MUX_bfv_3_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_28_0_\
        );

    \IN_MUX_bfv_3_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12871,
            carryinitout => \bfn_3_29_0_\
        );

    \IN_MUX_bfv_3_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12879,
            carryinitout => \bfn_3_30_0_\
        );

    \IN_MUX_bfv_3_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12887,
            carryinitout => \bfn_3_31_0_\
        );

    \IN_MUX_bfv_2_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_25_0_\
        );

    \IN_MUX_bfv_2_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12844,
            carryinitout => \bfn_2_26_0_\
        );

    \IN_MUX_bfv_2_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12852,
            carryinitout => \bfn_2_27_0_\
        );

    \IN_MUX_bfv_2_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12860,
            carryinitout => \bfn_2_28_0_\
        );

    \IN_MUX_bfv_1_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_22_0_\
        );

    \IN_MUX_bfv_1_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12818,
            carryinitout => \bfn_1_23_0_\
        );

    \IN_MUX_bfv_1_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12826,
            carryinitout => \bfn_1_24_0_\
        );

    \IN_MUX_bfv_1_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12834,
            carryinitout => \bfn_1_25_0_\
        );

    \IN_MUX_bfv_2_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_17_0_\
        );

    \IN_MUX_bfv_2_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12793,
            carryinitout => \bfn_2_18_0_\
        );

    \IN_MUX_bfv_2_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12801,
            carryinitout => \bfn_2_19_0_\
        );

    \IN_MUX_bfv_2_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12809,
            carryinitout => \bfn_2_20_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12769,
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12777,
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_2_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12785,
            carryinitout => \bfn_2_16_0_\
        );

    \IN_MUX_bfv_6_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_24_0_\
        );

    \IN_MUX_bfv_6_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12746,
            carryinitout => \bfn_6_25_0_\
        );

    \IN_MUX_bfv_6_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12754,
            carryinitout => \bfn_6_26_0_\
        );

    \IN_MUX_bfv_6_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_21_0_\
        );

    \IN_MUX_bfv_6_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12724,
            carryinitout => \bfn_6_22_0_\
        );

    \IN_MUX_bfv_6_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12732,
            carryinitout => \bfn_6_23_0_\
        );

    \IN_MUX_bfv_1_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_19_0_\
        );

    \IN_MUX_bfv_1_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12703,
            carryinitout => \bfn_1_20_0_\
        );

    \IN_MUX_bfv_1_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12711,
            carryinitout => \bfn_1_21_0_\
        );

    \IN_MUX_bfv_3_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_14_0_\
        );

    \IN_MUX_bfv_3_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12683,
            carryinitout => \bfn_3_15_0_\
        );

    \IN_MUX_bfv_3_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12691,
            carryinitout => \bfn_3_16_0_\
        );

    \IN_MUX_bfv_4_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_17_0_\
        );

    \IN_MUX_bfv_4_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12664,
            carryinitout => \bfn_4_18_0_\
        );

    \IN_MUX_bfv_4_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12672,
            carryinitout => \bfn_4_19_0_\
        );

    \IN_MUX_bfv_6_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_17_0_\
        );

    \IN_MUX_bfv_6_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12646,
            carryinitout => \bfn_6_18_0_\
        );

    \IN_MUX_bfv_6_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12654,
            carryinitout => \bfn_6_19_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_9_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12629,
            carryinitout => \bfn_9_17_0_\
        );

    \IN_MUX_bfv_9_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12637,
            carryinitout => \bfn_9_18_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12613,
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12621,
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_12_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12598,
            carryinitout => \bfn_12_21_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12584,
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_16_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_19_0_\
        );

    \IN_MUX_bfv_16_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12571,
            carryinitout => \bfn_16_20_0_\
        );

    \IN_MUX_bfv_9_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_29_0_\
        );

    \IN_MUX_bfv_1_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_31_0_\
        );

    \IN_MUX_bfv_1_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \debounce.n13020\,
            carryinitout => \bfn_1_32_0_\
        );

    \IN_MUX_bfv_10_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_29_0_\
        );

    \IN_MUX_bfv_10_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n13077,
            carryinitout => \bfn_10_30_0_\
        );

    \IN_MUX_bfv_10_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n13085,
            carryinitout => \bfn_10_31_0_\
        );

    \IN_MUX_bfv_10_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n13093,
            carryinitout => \bfn_10_32_0_\
        );

    \IN_MUX_bfv_7_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_25_0_\
        );

    \IN_MUX_bfv_7_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12959,
            carryinitout => \bfn_7_26_0_\
        );

    \IN_MUX_bfv_7_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n12967,
            carryinitout => \bfn_7_27_0_\
        );

    \IN_MUX_bfv_10_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_22_0_\
        );

    \IN_MUX_bfv_14_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_28_0_\
        );

    \IN_MUX_bfv_14_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWM.n13029\,
            carryinitout => \bfn_14_29_0_\
        );

    \IN_MUX_bfv_14_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWM.n13037\,
            carryinitout => \bfn_14_30_0_\
        );

    \IN_MUX_bfv_14_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PWM.n13045\,
            carryinitout => \bfn_14_31_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__21684\,
            GLOBALBUFFEROUTPUT => \CLK_N\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \i13072_1_lut_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35913\,
            lcout => n15802,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_2_lut_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38349\,
            in2 => \_gnd_net_\,
            in3 => \N__21690\,
            lcout => n2401,
            ltout => OPEN,
            carryin => \bfn_1_19_0_\,
            carryout => n12696,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_3_lut_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55031\,
            in2 => \N__29123\,
            in3 => \N__21687\,
            lcout => n2400,
            ltout => OPEN,
            carryin => n12696,
            carryout => n12697,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_4_lut_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28737\,
            in3 => \N__21717\,
            lcout => n2399,
            ltout => OPEN,
            carryin => n12697,
            carryout => n12698,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_5_lut_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55032\,
            in2 => \N__28637\,
            in3 => \N__21714\,
            lcout => n2398,
            ltout => OPEN,
            carryin => n12698,
            carryout => n12699,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_6_lut_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28832\,
            in3 => \N__21711\,
            lcout => n2397,
            ltout => OPEN,
            carryin => n12699,
            carryout => n12700,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_7_lut_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25904\,
            in3 => \N__21708\,
            lcout => n2396,
            ltout => OPEN,
            carryin => n12700,
            carryout => n12701,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_8_lut_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55418\,
            in2 => \N__25875\,
            in3 => \N__21705\,
            lcout => n2395,
            ltout => OPEN,
            carryin => n12701,
            carryout => n12702,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_9_lut_LC_1_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55033\,
            in2 => \N__25782\,
            in3 => \N__21702\,
            lcout => n2394,
            ltout => OPEN,
            carryin => n12702,
            carryout => n12703,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_10_lut_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55476\,
            in2 => \N__28863\,
            in3 => \N__21699\,
            lcout => n2393,
            ltout => OPEN,
            carryin => \bfn_1_20_0_\,
            carryout => n12704,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_11_lut_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55485\,
            in2 => \N__25653\,
            in3 => \N__21696\,
            lcout => n2392,
            ltout => OPEN,
            carryin => n12704,
            carryout => n12705,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_12_lut_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55477\,
            in2 => \N__23463\,
            in3 => \N__21693\,
            lcout => n2391,
            ltout => OPEN,
            carryin => n12705,
            carryout => n12706,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_13_lut_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55486\,
            in2 => \N__28922\,
            in3 => \N__21744\,
            lcout => n2390,
            ltout => OPEN,
            carryin => n12706,
            carryout => n12707,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_14_lut_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55478\,
            in2 => \N__28791\,
            in3 => \N__21741\,
            lcout => n2389,
            ltout => OPEN,
            carryin => n12707,
            carryout => n12708,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_15_lut_LC_1_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28688\,
            in2 => \N__55548\,
            in3 => \N__21738\,
            lcout => n2388,
            ltout => OPEN,
            carryin => n12708,
            carryout => n12709,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_16_lut_LC_1_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25623\,
            in2 => \N__55550\,
            in3 => \N__21735\,
            lcout => n2387,
            ltout => OPEN,
            carryin => n12709,
            carryout => n12710,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_17_lut_LC_1_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23439\,
            in2 => \N__55549\,
            in3 => \N__21732\,
            lcout => n2386,
            ltout => OPEN,
            carryin => n12710,
            carryout => n12711,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_18_lut_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28979\,
            in2 => \N__54721\,
            in3 => \N__21729\,
            lcout => n2385,
            ltout => OPEN,
            carryin => \bfn_1_21_0_\,
            carryout => n12712,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_19_lut_LC_1_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29024\,
            in2 => \N__54724\,
            in3 => \N__21726\,
            lcout => n2384,
            ltout => OPEN,
            carryin => n12712,
            carryout => n12713,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_20_lut_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25731\,
            in2 => \N__54722\,
            in3 => \N__21723\,
            lcout => n2383,
            ltout => OPEN,
            carryin => n12713,
            carryout => n12714,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_21_lut_LC_1_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30963\,
            in2 => \N__54725\,
            in3 => \N__21720\,
            lcout => n2382,
            ltout => OPEN,
            carryin => n12714,
            carryout => n12715,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_22_lut_LC_1_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25695\,
            in2 => \N__54723\,
            in3 => \N__21771\,
            lcout => n2381,
            ltout => OPEN,
            carryin => n12715,
            carryout => n12716,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1570_23_lut_LC_1_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__54324\,
            in1 => \N__35765\,
            in2 => \N__25812\,
            in3 => \N__21768\,
            lcout => n2412,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_2_lut_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33501\,
            in2 => \_gnd_net_\,
            in3 => \N__21765\,
            lcout => n2901,
            ltout => OPEN,
            carryin => \bfn_1_22_0_\,
            carryout => n12811,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_3_lut_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54708\,
            in2 => \N__26577\,
            in3 => \N__21762\,
            lcout => n2900,
            ltout => OPEN,
            carryin => n12811,
            carryout => n12812,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_4_lut_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29460\,
            in3 => \N__21759\,
            lcout => n2899,
            ltout => OPEN,
            carryin => n12812,
            carryout => n12813,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_5_lut_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54709\,
            in2 => \N__29649\,
            in3 => \N__21756\,
            lcout => n2898,
            ltout => OPEN,
            carryin => n12813,
            carryout => n12814,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_6_lut_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26544\,
            in3 => \N__21753\,
            lcout => n2897,
            ltout => OPEN,
            carryin => n12814,
            carryout => n12815,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_7_lut_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29884\,
            in3 => \N__21750\,
            lcout => n2896,
            ltout => OPEN,
            carryin => n12815,
            carryout => n12816,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_8_lut_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22757\,
            in2 => \N__55030\,
            in3 => \N__21747\,
            lcout => n2895,
            ltout => OPEN,
            carryin => n12816,
            carryout => n12817,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_9_lut_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54713\,
            in2 => \N__24584\,
            in3 => \N__21798\,
            lcout => n2894,
            ltout => OPEN,
            carryin => n12817,
            carryout => n12818,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_10_lut_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54283\,
            in2 => \N__29732\,
            in3 => \N__21795\,
            lcout => n2893,
            ltout => OPEN,
            carryin => \bfn_1_23_0_\,
            carryout => n12819,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_11_lut_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26740\,
            in2 => \N__54705\,
            in3 => \N__21792\,
            lcout => n2892,
            ltout => OPEN,
            carryin => n12819,
            carryout => n12820,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_12_lut_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54287\,
            in2 => \N__29336\,
            in3 => \N__21789\,
            lcout => n2891,
            ltout => OPEN,
            carryin => n12820,
            carryout => n12821,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_13_lut_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54292\,
            in2 => \N__24621\,
            in3 => \N__21786\,
            lcout => n2890,
            ltout => OPEN,
            carryin => n12821,
            carryout => n12822,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_14_lut_LC_1_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54288\,
            in2 => \N__24542\,
            in3 => \N__21783\,
            lcout => n2889,
            ltout => OPEN,
            carryin => n12822,
            carryout => n12823,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_15_lut_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54293\,
            in2 => \N__29831\,
            in3 => \N__21780\,
            lcout => n2888,
            ltout => OPEN,
            carryin => n12823,
            carryout => n12824,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_16_lut_LC_1_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24309\,
            in2 => \N__54707\,
            in3 => \N__21777\,
            lcout => n2887,
            ltout => OPEN,
            carryin => n12824,
            carryout => n12825,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_17_lut_LC_1_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26844\,
            in2 => \N__54706\,
            in3 => \N__21774\,
            lcout => n2886,
            ltout => OPEN,
            carryin => n12825,
            carryout => n12826,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_18_lut_LC_1_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26292\,
            in2 => \N__54240\,
            in3 => \N__21825\,
            lcout => n2885,
            ltout => OPEN,
            carryin => \bfn_1_24_0_\,
            carryout => n12827,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_19_lut_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27235\,
            in2 => \N__55275\,
            in3 => \N__21822\,
            lcout => n2884,
            ltout => OPEN,
            carryin => n12827,
            carryout => n12828,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_20_lut_LC_1_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26337\,
            in2 => \N__54241\,
            in3 => \N__21819\,
            lcout => n2883,
            ltout => OPEN,
            carryin => n12828,
            carryout => n12829,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_21_lut_LC_1_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53834\,
            in2 => \N__26504\,
            in3 => \N__21816\,
            lcout => n2882,
            ltout => OPEN,
            carryin => n12829,
            carryout => n12830,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_22_lut_LC_1_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29767\,
            in2 => \N__54242\,
            in3 => \N__21813\,
            lcout => n2881,
            ltout => OPEN,
            carryin => n12830,
            carryout => n12831,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_23_lut_LC_1_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26447\,
            in2 => \N__55276\,
            in3 => \N__21810\,
            lcout => n2880,
            ltout => OPEN,
            carryin => n12831,
            carryout => n12832,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_24_lut_LC_1_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26471\,
            in2 => \N__54243\,
            in3 => \N__21807\,
            lcout => n2879,
            ltout => OPEN,
            carryin => n12832,
            carryout => n12833,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_25_lut_LC_1_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26418\,
            in2 => \N__55277\,
            in3 => \N__21804\,
            lcout => n2878,
            ltout => OPEN,
            carryin => n12833,
            carryout => n12834,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_26_lut_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26901\,
            in2 => \N__54654\,
            in3 => \N__21801\,
            lcout => n2877,
            ltout => OPEN,
            carryin => \bfn_1_25_0_\,
            carryout => n12835,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_27_lut_LC_1_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26402\,
            in2 => \N__54655\,
            in3 => \N__21858\,
            lcout => n2876,
            ltout => OPEN,
            carryin => n12835,
            carryout => n12836,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1905_28_lut_LC_1_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__54236\,
            in1 => \N__34352\,
            in2 => \N__26367\,
            in3 => \N__21855\,
            lcout => n2907,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1914_3_lut_LC_1_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26500\,
            in2 => \N__34333\,
            in3 => \N__21852\,
            lcout => n2914,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1932_3_lut_LC_1_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__26572\,
            in1 => \_gnd_net_\,
            in2 => \N__21846\,
            in3 => \N__34316\,
            lcout => n2932,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1847_3_lut_LC_1_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36411\,
            in2 => \N__22365\,
            in3 => \N__22845\,
            lcout => n2815,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1778_3_lut_LC_1_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22245\,
            in2 => \N__29688\,
            in3 => \N__36295\,
            lcout => n2714,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.reg_out_i0_i0_LC_1_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46927\,
            in1 => \N__21921\,
            in2 => \_gnd_net_\,
            in3 => \N__38870\,
            lcout => h3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56199\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1908_3_lut_LC_1_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21834\,
            in2 => \N__34335\,
            in3 => \N__26403\,
            lcout => n2908,
            ltout => \n2908_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1975_3_lut_LC_1_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34513\,
            in1 => \_gnd_net_\,
            in2 => \N__21828\,
            in3 => \N__23028\,
            lcout => n3007,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1865_3_lut_LC_1_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22296\,
            in1 => \N__33539\,
            in2 => \_gnd_net_\,
            in3 => \N__36417\,
            lcout => n2833,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1927_3_lut_LC_1_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21879\,
            in2 => \N__22761\,
            in3 => \N__34328\,
            lcout => n2927,
            ltout => \n2927_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1994_3_lut_LC_1_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__22881\,
            in1 => \_gnd_net_\,
            in2 => \N__21867\,
            in3 => \N__34512\,
            lcout => n3026,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1993_3_lut_LC_1_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__22962\,
            in1 => \_gnd_net_\,
            in2 => \N__34509\,
            in3 => \N__26781\,
            lcout => n3025,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1990_3_lut_LC_1_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29301\,
            in2 => \N__22941\,
            in3 => \N__34483\,
            lcout => n3022,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1985_3_lut_LC_1_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__26817\,
            in1 => \N__23004\,
            in2 => \N__34511\,
            in3 => \_gnd_net_\,
            lcout => n3017,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1992_3_lut_LC_1_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22953\,
            in2 => \N__29715\,
            in3 => \N__34493\,
            lcout => n3024,
            ltout => \n3024_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_166_LC_1_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24736\,
            in1 => \N__24935\,
            in2 => \N__21864\,
            in3 => \N__24778\,
            lcout => OPEN,
            ltout => \n14730_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_168_LC_1_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24880\,
            in1 => \N__27278\,
            in2 => \N__21861\,
            in3 => \N__21897\,
            lcout => n14736,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1989_3_lut_LC_1_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22929\,
            in2 => \N__34510\,
            in3 => \N__26682\,
            lcout => n3021,
            ltout => \n3021_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_165_LC_1_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25006\,
            in2 => \N__21900\,
            in3 => \N__24830\,
            lcout => n14728,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_174_LC_1_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27968\,
            in1 => \N__32905\,
            in2 => \N__30811\,
            in3 => \N__27802\,
            lcout => OPEN,
            ltout => \n14150_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_176_LC_1_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30658\,
            in1 => \N__21885\,
            in2 => \N__21891\,
            in3 => \N__21975\,
            lcout => n14156,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1977_3_lut_LC_1_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27072\,
            in2 => \N__22974\,
            in3 => \N__34514\,
            lcout => n3009,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2062_3_lut_LC_1_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24804\,
            in2 => \N__30597\,
            in3 => \N__34710\,
            lcout => n3126,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2064_3_lut_LC_1_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__24843\,
            in1 => \_gnd_net_\,
            in2 => \N__34716\,
            in3 => \N__29958\,
            lcout => n3128,
            ltout => \n3128_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_175_LC_1_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27676\,
            in1 => \N__27751\,
            in2 => \N__21888\,
            in3 => \N__27735\,
            lcout => n14148,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.reg_B_i0_LC_1_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21942\,
            lcout => \reg_B_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56203\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2054_3_lut_LC_1_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30623\,
            in2 => \N__34708\,
            in3 => \N__24903\,
            lcout => n3118,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2060_3_lut_LC_1_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__24746\,
            in1 => \_gnd_net_\,
            in2 => \N__34709\,
            in3 => \N__24723\,
            lcout => n3124,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2056_3_lut_LC_1_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24951\,
            in2 => \N__24978\,
            in3 => \N__34681\,
            lcout => n3120,
            ltout => \n3120_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2123_3_lut_LC_1_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23085\,
            in2 => \N__21981\,
            in3 => \N__34911\,
            lcout => n3219,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2058_3_lut_LC_1_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30560\,
            in2 => \N__25035\,
            in3 => \N__34686\,
            lcout => n3122,
            ltout => \n3122_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_173_LC_1_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30883\,
            in1 => \N__23096\,
            in2 => \N__21978\,
            in3 => \N__27544\,
            lcout => n14146,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2059_3_lut_LC_1_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24707\,
            in2 => \N__24687\,
            in3 => \N__34682\,
            lcout => n3123,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.reg_B_i2_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21969\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \reg_B_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56207\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.reg_B_i1_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21959\,
            lcout => \reg_B_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56207\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.i2_4_lut_LC_1_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__21968\,
            in1 => \N__38885\,
            in2 => \N__21960\,
            in3 => \N__22070\,
            lcout => OPEN,
            ltout => \debounce.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.i3_4_lut_LC_1_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011011111111"
        )
    port map (
            in0 => \N__21941\,
            in1 => \N__21920\,
            in2 => \N__21903\,
            in3 => \N__38857\,
            lcout => \debounce.cnt_next_9__N_424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.i7_4_lut_LC_1_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__21995\,
            in1 => \N__22149\,
            in2 => \N__22128\,
            in3 => \N__22193\,
            lcout => \debounce.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.i6_4_lut_LC_1_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__22163\,
            in1 => \N__22058\,
            in2 => \N__22029\,
            in3 => \N__22043\,
            lcout => OPEN,
            ltout => \debounce.n16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.i9_4_lut_LC_1_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__22010\,
            in1 => \N__22178\,
            in2 => \N__22080\,
            in3 => \N__22077\,
            lcout => n14129,
            ltout => \n14129_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.reg_out_i0_i2_LC_1_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__22071\,
            in1 => \_gnd_net_\,
            in2 => \N__22062\,
            in3 => \N__46866\,
            lcout => h1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56207\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.cnt_reg_665__i0_LC_1_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22059\,
            in2 => \_gnd_net_\,
            in3 => \N__22047\,
            lcout => \debounce.cnt_reg_0\,
            ltout => OPEN,
            carryin => \bfn_1_31_0_\,
            carryout => \debounce.n13013\,
            clk => \N__56208\,
            ce => 'H',
            sr => \N__22106\
        );

    \debounce.cnt_reg_665__i1_LC_1_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22044\,
            in2 => \_gnd_net_\,
            in3 => \N__22032\,
            lcout => \debounce.cnt_reg_1\,
            ltout => OPEN,
            carryin => \debounce.n13013\,
            carryout => \debounce.n13014\,
            clk => \N__56208\,
            ce => 'H',
            sr => \N__22106\
        );

    \debounce.cnt_reg_665__i2_LC_1_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22028\,
            in2 => \_gnd_net_\,
            in3 => \N__22014\,
            lcout => \debounce.cnt_reg_2\,
            ltout => OPEN,
            carryin => \debounce.n13014\,
            carryout => \debounce.n13015\,
            clk => \N__56208\,
            ce => 'H',
            sr => \N__22106\
        );

    \debounce.cnt_reg_665__i3_LC_1_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22011\,
            in2 => \_gnd_net_\,
            in3 => \N__21999\,
            lcout => \debounce.cnt_reg_3\,
            ltout => OPEN,
            carryin => \debounce.n13015\,
            carryout => \debounce.n13016\,
            clk => \N__56208\,
            ce => 'H',
            sr => \N__22106\
        );

    \debounce.cnt_reg_665__i4_LC_1_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21996\,
            in2 => \_gnd_net_\,
            in3 => \N__21984\,
            lcout => \debounce.cnt_reg_4\,
            ltout => OPEN,
            carryin => \debounce.n13016\,
            carryout => \debounce.n13017\,
            clk => \N__56208\,
            ce => 'H',
            sr => \N__22106\
        );

    \debounce.cnt_reg_665__i5_LC_1_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22194\,
            in2 => \_gnd_net_\,
            in3 => \N__22182\,
            lcout => \debounce.cnt_reg_5\,
            ltout => OPEN,
            carryin => \debounce.n13017\,
            carryout => \debounce.n13018\,
            clk => \N__56208\,
            ce => 'H',
            sr => \N__22106\
        );

    \debounce.cnt_reg_665__i6_LC_1_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22179\,
            in2 => \_gnd_net_\,
            in3 => \N__22167\,
            lcout => \debounce.cnt_reg_6\,
            ltout => OPEN,
            carryin => \debounce.n13018\,
            carryout => \debounce.n13019\,
            clk => \N__56208\,
            ce => 'H',
            sr => \N__22106\
        );

    \debounce.cnt_reg_665__i7_LC_1_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22164\,
            in2 => \_gnd_net_\,
            in3 => \N__22152\,
            lcout => \debounce.cnt_reg_7\,
            ltout => OPEN,
            carryin => \debounce.n13019\,
            carryout => \debounce.n13020\,
            clk => \N__56208\,
            ce => 'H',
            sr => \N__22106\
        );

    \debounce.cnt_reg_665__i8_LC_1_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22148\,
            in2 => \_gnd_net_\,
            in3 => \N__22134\,
            lcout => \debounce.cnt_reg_8\,
            ltout => OPEN,
            carryin => \bfn_1_32_0_\,
            carryout => \debounce.n13021\,
            clk => \N__56210\,
            ce => 'H',
            sr => \N__22110\
        );

    \debounce.cnt_reg_665__i9_LC_1_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22124\,
            in2 => \_gnd_net_\,
            in3 => \N__22131\,
            lcout => \debounce.cnt_reg_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56210\,
            ce => 'H',
            sr => \N__22110\
        );

    \encoder0_position_31__I_0_add_1771_2_lut_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33582\,
            in2 => \_gnd_net_\,
            in3 => \N__22089\,
            lcout => n2701,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => n12762,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_3_lut_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26265\,
            in2 => \N__55563\,
            in3 => \N__22086\,
            lcout => n2700,
            ltout => OPEN,
            carryin => n12762,
            carryout => n12763,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_4_lut_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29259\,
            in3 => \N__22083\,
            lcout => n2699,
            ltout => OPEN,
            carryin => n12763,
            carryout => n12764,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_5_lut_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55436\,
            in2 => \N__29196\,
            in3 => \N__22224\,
            lcout => n2698,
            ltout => OPEN,
            carryin => n12764,
            carryout => n12765,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_6_lut_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29439\,
            in3 => \N__22221\,
            lcout => n2697,
            ltout => OPEN,
            carryin => n12765,
            carryout => n12766,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_7_lut_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29508\,
            in3 => \N__22218\,
            lcout => n2696,
            ltout => OPEN,
            carryin => n12766,
            carryout => n12767,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_8_lut_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55562\,
            in2 => \N__23589\,
            in3 => \N__22215\,
            lcout => n2695,
            ltout => OPEN,
            carryin => n12767,
            carryout => n12768,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_9_lut_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55437\,
            in2 => \N__29076\,
            in3 => \N__22212\,
            lcout => n2694,
            ltout => OPEN,
            carryin => n12768,
            carryout => n12769,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_10_lut_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55426\,
            in2 => \N__26037\,
            in3 => \N__22209\,
            lcout => n2693,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => n12770,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_11_lut_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55433\,
            in2 => \N__25971\,
            in3 => \N__22206\,
            lcout => n2692,
            ltout => OPEN,
            carryin => n12770,
            carryout => n12771,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_12_lut_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55427\,
            in2 => \N__33921\,
            in3 => \N__22203\,
            lcout => n2691,
            ltout => OPEN,
            carryin => n12771,
            carryout => n12772,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_13_lut_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24128\,
            in2 => \N__55535\,
            in3 => \N__22200\,
            lcout => n2690,
            ltout => OPEN,
            carryin => n12772,
            carryout => n12773,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_14_lut_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55431\,
            in2 => \N__23676\,
            in3 => \N__22197\,
            lcout => n2689,
            ltout => OPEN,
            carryin => n12773,
            carryout => n12774,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_15_lut_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55434\,
            in2 => \N__23880\,
            in3 => \N__22263\,
            lcout => n2688,
            ltout => OPEN,
            carryin => n12774,
            carryout => n12775,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_16_lut_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55432\,
            in2 => \N__29394\,
            in3 => \N__22260\,
            lcout => n2687,
            ltout => OPEN,
            carryin => n12775,
            carryout => n12776,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_17_lut_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55435\,
            in2 => \N__26148\,
            in3 => \N__22257\,
            lcout => n2686,
            ltout => OPEN,
            carryin => n12776,
            carryout => n12777,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_18_lut_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26235\,
            in2 => \N__55551\,
            in3 => \N__22254\,
            lcout => n2685,
            ltout => OPEN,
            carryin => \bfn_2_15_0_\,
            carryout => n12778,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_19_lut_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25997\,
            in2 => \N__55555\,
            in3 => \N__22251\,
            lcout => n2684,
            ltout => OPEN,
            carryin => n12778,
            carryout => n12779,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_20_lut_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32628\,
            in2 => \N__55552\,
            in3 => \N__22248\,
            lcout => n2683,
            ltout => OPEN,
            carryin => n12779,
            carryout => n12780,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_21_lut_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29684\,
            in2 => \N__55556\,
            in3 => \N__22233\,
            lcout => n2682,
            ltout => OPEN,
            carryin => n12780,
            carryout => n12781,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_22_lut_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26208\,
            in2 => \N__55553\,
            in3 => \N__22230\,
            lcout => n2681,
            ltout => OPEN,
            carryin => n12781,
            carryout => n12782,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_23_lut_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26175\,
            in2 => \N__55557\,
            in3 => \N__22227\,
            lcout => n2680,
            ltout => OPEN,
            carryin => n12782,
            carryout => n12783,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_24_lut_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29544\,
            in2 => \N__55554\,
            in3 => \N__22305\,
            lcout => n2679,
            ltout => OPEN,
            carryin => n12783,
            carryout => n12784,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_25_lut_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32559\,
            in2 => \N__55558\,
            in3 => \N__22302\,
            lcout => n2678,
            ltout => OPEN,
            carryin => n12784,
            carryout => n12785,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1771_26_lut_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54743\,
            in2 => \N__32736\,
            in3 => \N__22299\,
            lcout => n2677,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_2_lut_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33540\,
            in2 => \_gnd_net_\,
            in3 => \N__22281\,
            lcout => n2801,
            ltout => OPEN,
            carryin => \bfn_2_17_0_\,
            carryout => n12786,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_3_lut_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55493\,
            in2 => \N__26628\,
            in3 => \N__22278\,
            lcout => n2800,
            ltout => OPEN,
            carryin => n12786,
            carryout => n12787,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_4_lut_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24078\,
            in3 => \N__22275\,
            lcout => n2799,
            ltout => OPEN,
            carryin => n12787,
            carryout => n12788,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_5_lut_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55494\,
            in2 => \N__24369\,
            in3 => \N__22272\,
            lcout => n2798,
            ltout => OPEN,
            carryin => n12788,
            carryout => n12789,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_6_lut_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23838\,
            in3 => \N__22269\,
            lcout => n2797,
            ltout => OPEN,
            carryin => n12789,
            carryout => n12790,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_7_lut_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23916\,
            in2 => \_gnd_net_\,
            in3 => \N__22266\,
            lcout => n2796,
            ltout => OPEN,
            carryin => n12790,
            carryout => n12791,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_8_lut_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55496\,
            in2 => \N__23733\,
            in3 => \N__22332\,
            lcout => n2795,
            ltout => OPEN,
            carryin => n12791,
            carryout => n12792,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_9_lut_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55495\,
            in2 => \N__23562\,
            in3 => \N__22329\,
            lcout => n2794,
            ltout => OPEN,
            carryin => n12792,
            carryout => n12793,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_10_lut_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55349\,
            in2 => \N__23715\,
            in3 => \N__22326\,
            lcout => n2793,
            ltout => OPEN,
            carryin => \bfn_2_18_0_\,
            carryout => n12794,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_11_lut_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55355\,
            in2 => \N__22698\,
            in3 => \N__22323\,
            lcout => n2792,
            ltout => OPEN,
            carryin => n12794,
            carryout => n12795,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_12_lut_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55350\,
            in2 => \N__23637\,
            in3 => \N__22320\,
            lcout => n2791,
            ltout => OPEN,
            carryin => n12795,
            carryout => n12796,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_13_lut_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55356\,
            in2 => \N__22512\,
            in3 => \N__22317\,
            lcout => n2790,
            ltout => OPEN,
            carryin => n12796,
            carryout => n12797,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_14_lut_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55351\,
            in2 => \N__24102\,
            in3 => \N__22314\,
            lcout => n2789,
            ltout => OPEN,
            carryin => n12797,
            carryout => n12798,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_15_lut_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55357\,
            in2 => \N__23756\,
            in3 => \N__22311\,
            lcout => n2788,
            ltout => OPEN,
            carryin => n12798,
            carryout => n12799,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_16_lut_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24227\,
            in2 => \N__55492\,
            in3 => \N__22308\,
            lcout => n2787,
            ltout => OPEN,
            carryin => n12799,
            carryout => n12800,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_17_lut_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23990\,
            in2 => \N__55491\,
            in3 => \N__22374\,
            lcout => n2786,
            ltout => OPEN,
            carryin => n12800,
            carryout => n12801,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_18_lut_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24165\,
            in2 => \N__55526\,
            in3 => \N__22371\,
            lcout => n2785,
            ltout => OPEN,
            carryin => \bfn_2_19_0_\,
            carryout => n12802,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_19_lut_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23952\,
            in2 => \N__55530\,
            in3 => \N__22368\,
            lcout => n2784,
            ltout => OPEN,
            carryin => n12802,
            carryout => n12803,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_20_lut_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22844\,
            in2 => \N__55527\,
            in3 => \N__22350\,
            lcout => n2783,
            ltout => OPEN,
            carryin => n12803,
            carryout => n12804,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_21_lut_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22582\,
            in2 => \N__55531\,
            in3 => \N__22347\,
            lcout => n2782,
            ltout => OPEN,
            carryin => n12804,
            carryout => n12805,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_22_lut_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24279\,
            in2 => \N__55528\,
            in3 => \N__22344\,
            lcout => n2781,
            ltout => OPEN,
            carryin => n12805,
            carryout => n12806,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_23_lut_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24417\,
            in2 => \N__55532\,
            in3 => \N__22341\,
            lcout => n2780,
            ltout => OPEN,
            carryin => n12806,
            carryout => n12807,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_24_lut_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26106\,
            in2 => \N__55529\,
            in3 => \N__22338\,
            lcout => n2779,
            ltout => OPEN,
            carryin => n12807,
            carryout => n12808,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_25_lut_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24039\,
            in2 => \N__55533\,
            in3 => \N__22335\,
            lcout => n2778,
            ltout => OPEN,
            carryin => n12808,
            carryout => n12809,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_26_lut_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24463\,
            in2 => \N__55547\,
            in3 => \N__22452\,
            lcout => n2777,
            ltout => OPEN,
            carryin => \bfn_2_20_0_\,
            carryout => n12810,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1838_27_lut_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__53967\,
            in1 => \N__22799\,
            in2 => \N__36491\,
            in3 => \N__22449\,
            lcout => n2808,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1779_3_lut_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32624\,
            in2 => \N__36293\,
            in3 => \N__22446\,
            lcout => n2715,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1773_3_lut_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32732\,
            in2 => \N__22437\,
            in3 => \N__36275\,
            lcout => n2709,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1774_3_lut_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__32555\,
            in1 => \_gnd_net_\,
            in2 => \N__36294\,
            in3 => \N__22422\,
            lcout => n2710,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13045_1_lut_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35744\,
            lcout => n15775,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1861_3_lut_LC_2_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22413\,
            in2 => \N__36453\,
            in3 => \N__23831\,
            lcout => n2829,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1790_3_lut_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29069\,
            in2 => \N__22404\,
            in3 => \N__36262\,
            lcout => n2726,
            ltout => \n2726_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1857_3_lut_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__36422\,
            in1 => \N__22389\,
            in2 => \N__22377\,
            in3 => \_gnd_net_\,
            lcout => n2825,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1717_3_lut_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__34086\,
            in1 => \_gnd_net_\,
            in2 => \N__32484\,
            in3 => \N__36095\,
            lcout => n2621,
            ltout => \n2621_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1784_3_lut_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__36266\,
            in1 => \_gnd_net_\,
            in2 => \N__22566\,
            in3 => \N__22563\,
            lcout => n2720,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1792_3_lut_LC_2_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29501\,
            in2 => \N__36292\,
            in3 => \N__22551\,
            lcout => n2728,
            ltout => \n2728_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1859_3_lut_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22536\,
            in2 => \N__22527\,
            in3 => \N__36418\,
            lcout => n2827,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_54_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22502\,
            in1 => \N__23551\,
            in2 => \N__22690\,
            in3 => \N__24220\,
            lcout => n14346,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1787_3_lut_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33917\,
            in2 => \N__22524\,
            in3 => \N__36234\,
            lcout => n2723,
            ltout => \n2723_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1854_3_lut_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22491\,
            in2 => \N__22479\,
            in3 => \N__36423\,
            lcout => n2822,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1789_3_lut_LC_2_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22476\,
            in2 => \N__26033\,
            in3 => \N__36235\,
            lcout => n2725,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1793_3_lut_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29434\,
            in2 => \N__36279\,
            in3 => \N__22467\,
            lcout => n2729,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1777_3_lut_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26207\,
            in2 => \N__22665\,
            in3 => \N__36239\,
            lcout => n2713,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1858_3_lut_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23552\,
            in2 => \N__22650\,
            in3 => \N__36424\,
            lcout => n2826,
            ltout => \n2826_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_61_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22756\,
            in1 => \N__24577\,
            in2 => \N__22635\,
            in3 => \N__24535\,
            lcout => n14688,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_59_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23886\,
            in1 => \N__22583\,
            in2 => \N__22843\,
            in3 => \N__22605\,
            lcout => OPEN,
            ltout => \n14362_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_60_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24278\,
            in1 => \N__26098\,
            in2 => \N__22632\,
            in3 => \N__24415\,
            lcout => n14368,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1853_3_lut_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24092\,
            in2 => \N__36445\,
            in3 => \N__22629\,
            lcout => n2821,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_56_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__24091\,
            in1 => \_gnd_net_\,
            in2 => \N__22617\,
            in3 => \N__23983\,
            lcout => OPEN,
            ltout => \n14350_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_57_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23694\,
            in1 => \N__24157\,
            in2 => \N__22608\,
            in3 => \N__23945\,
            lcout => n14356,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1846_3_lut_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22599\,
            in2 => \N__22587\,
            in3 => \N__36408\,
            lcout => n2814,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1849_3_lut_LC_2_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24158\,
            in2 => \N__36446\,
            in3 => \N__22872\,
            lcout => n2817,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1780_3_lut_LC_2_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22860\,
            in2 => \N__25998\,
            in3 => \N__36258\,
            lcout => n2716,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1775_3_lut_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__29540\,
            in1 => \_gnd_net_\,
            in2 => \N__22818\,
            in3 => \N__36245\,
            lcout => n2711,
            ltout => \n2711_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12595_4_lut_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22800\,
            in1 => \N__24467\,
            in2 => \N__22785\,
            in3 => \N__22782\,
            lcout => n2742,
            ltout => \n2742_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1860_3_lut_LC_2_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22776\,
            in2 => \N__22764\,
            in3 => \N__23915\,
            lcout => n2828,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12592_1_lut_LC_2_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36437\,
            lcout => n15322,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1852_3_lut_LC_2_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23757\,
            in2 => \N__36457\,
            in3 => \N__22731\,
            lcout => n2820,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1783_3_lut_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29387\,
            in2 => \N__36280\,
            in3 => \N__22719\,
            lcout => n2719,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1856_3_lut_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22707\,
            in2 => \N__36456\,
            in3 => \N__22694\,
            lcout => n2824,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1855_3_lut_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__22911\,
            in1 => \_gnd_net_\,
            in2 => \N__23636\,
            in3 => \N__36438\,
            lcout => n2823,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_2_lut_LC_2_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35178\,
            in2 => \_gnd_net_\,
            in3 => \N__22902\,
            lcout => n3001,
            ltout => OPEN,
            carryin => \bfn_2_25_0_\,
            carryout => n12837,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_3_lut_LC_2_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30222\,
            in2 => \N__55083\,
            in3 => \N__22899\,
            lcout => n3000,
            ltout => OPEN,
            carryin => n12837,
            carryout => n12838,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_4_lut_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30130\,
            in2 => \_gnd_net_\,
            in3 => \N__22896\,
            lcout => n2999,
            ltout => OPEN,
            carryin => n12838,
            carryout => n12839,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_5_lut_LC_2_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30007\,
            in2 => \N__55084\,
            in3 => \N__22893\,
            lcout => n2998,
            ltout => OPEN,
            carryin => n12839,
            carryout => n12840,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_6_lut_LC_2_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29598\,
            in3 => \N__22890\,
            lcout => n2997,
            ltout => OPEN,
            carryin => n12840,
            carryout => n12841,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_7_lut_LC_2_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27167\,
            in3 => \N__22887\,
            lcout => n2996,
            ltout => OPEN,
            carryin => n12841,
            carryout => n12842,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_8_lut_LC_2_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29856\,
            in2 => \N__55066\,
            in3 => \N__22884\,
            lcout => n2995,
            ltout => OPEN,
            carryin => n12842,
            carryout => n12843,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_9_lut_LC_2_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26795\,
            in2 => \N__55085\,
            in3 => \N__22875\,
            lcout => n2994,
            ltout => OPEN,
            carryin => n12843,
            carryout => n12844,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_10_lut_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26774\,
            in2 => \N__55062\,
            in3 => \N__22956\,
            lcout => n2993,
            ltout => OPEN,
            carryin => \bfn_2_26_0_\,
            carryout => n12845,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_11_lut_LC_2_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29708\,
            in2 => \N__55080\,
            in3 => \N__22947\,
            lcout => n2992,
            ltout => OPEN,
            carryin => n12845,
            carryout => n12846,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_12_lut_LC_2_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29562\,
            in2 => \N__55063\,
            in3 => \N__22944\,
            lcout => n2991,
            ltout => OPEN,
            carryin => n12846,
            carryout => n12847,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_13_lut_LC_2_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54813\,
            in2 => \N__29300\,
            in3 => \N__22932\,
            lcout => n2990,
            ltout => OPEN,
            carryin => n12847,
            carryout => n12848,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_14_lut_LC_2_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26675\,
            in2 => \N__55064\,
            in3 => \N__22923\,
            lcout => n2989,
            ltout => OPEN,
            carryin => n12848,
            carryout => n12849,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_15_lut_LC_2_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26699\,
            in2 => \N__55081\,
            in3 => \N__22920\,
            lcout => n2988,
            ltout => OPEN,
            carryin => n12849,
            carryout => n12850,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_16_lut_LC_2_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30179\,
            in2 => \N__55065\,
            in3 => \N__22917\,
            lcout => n2987,
            ltout => OPEN,
            carryin => n12850,
            carryout => n12851,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_17_lut_LC_2_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26654\,
            in2 => \N__55082\,
            in3 => \N__22914\,
            lcout => n2986,
            ltout => OPEN,
            carryin => n12851,
            carryout => n12852,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_18_lut_LC_2_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26813\,
            in2 => \N__55058\,
            in3 => \N__22998\,
            lcout => n2985,
            ltout => OPEN,
            carryin => \bfn_2_27_0_\,
            carryout => n12853,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_19_lut_LC_2_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30368\,
            in2 => \N__55076\,
            in3 => \N__22995\,
            lcout => n2984,
            ltout => OPEN,
            carryin => n12853,
            carryout => n12854,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_20_lut_LC_2_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27204\,
            in2 => \N__55059\,
            in3 => \N__22992\,
            lcout => n2983,
            ltout => OPEN,
            carryin => n12854,
            carryout => n12855,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_21_lut_LC_2_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27123\,
            in2 => \N__55077\,
            in3 => \N__22989\,
            lcout => n2982,
            ltout => OPEN,
            carryin => n12855,
            carryout => n12856,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_22_lut_LC_2_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27093\,
            in2 => \N__55060\,
            in3 => \N__22986\,
            lcout => n2981,
            ltout => OPEN,
            carryin => n12856,
            carryout => n12857,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_23_lut_LC_2_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30294\,
            in2 => \N__55078\,
            in3 => \N__22983\,
            lcout => n2980,
            ltout => OPEN,
            carryin => n12857,
            carryout => n12858,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_24_lut_LC_2_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27042\,
            in2 => \N__55061\,
            in3 => \N__22980\,
            lcout => n2979,
            ltout => OPEN,
            carryin => n12858,
            carryout => n12859,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_25_lut_LC_2_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26937\,
            in2 => \N__55079\,
            in3 => \N__22977\,
            lcout => n2978,
            ltout => OPEN,
            carryin => n12859,
            carryout => n12860,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_26_lut_LC_2_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27071\,
            in2 => \N__55057\,
            in3 => \N__22965\,
            lcout => n2977,
            ltout => OPEN,
            carryin => \bfn_2_28_0_\,
            carryout => n12861,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_27_lut_LC_2_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54792\,
            in2 => \N__26979\,
            in3 => \N__23031\,
            lcout => n2976,
            ltout => OPEN,
            carryin => n12861,
            carryout => n12862,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_28_lut_LC_2_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54793\,
            in2 => \N__27030\,
            in3 => \N__23019\,
            lcout => n2975,
            ltout => OPEN,
            carryin => n12862,
            carryout => n12863,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1972_29_lut_LC_2_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__54794\,
            in1 => \N__27002\,
            in2 => \N__34532\,
            in3 => \N__23016\,
            lcout => n3006,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2061_3_lut_LC_2_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24788\,
            in2 => \N__24762\,
            in3 => \N__34649\,
            lcout => n3125,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2055_3_lut_LC_2_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24912\,
            in2 => \N__34695\,
            in3 => \N__24934\,
            lcout => n3119,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2057_3_lut_LC_2_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25010\,
            in2 => \N__24990\,
            in3 => \N__34653\,
            lcout => n3121,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2052_3_lut_LC_2_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24864\,
            in2 => \N__34696\,
            in3 => \N__24884\,
            lcout => n3116,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_2_lut_LC_2_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34170\,
            in2 => \_gnd_net_\,
            in3 => \N__23013\,
            lcout => n3201,
            ltout => OPEN,
            carryin => \bfn_2_29_0_\,
            carryout => n12892,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_3_lut_LC_2_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54572\,
            in2 => \N__30432\,
            in3 => \N__23010\,
            lcout => n3200,
            ltout => OPEN,
            carryin => n12892,
            carryout => n12893,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_4_lut_LC_2_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30510\,
            in3 => \N__23007\,
            lcout => n3199,
            ltout => OPEN,
            carryin => n12893,
            carryout => n12894,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_5_lut_LC_2_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54573\,
            in2 => \N__30396\,
            in3 => \N__23058\,
            lcout => n3198,
            ltout => OPEN,
            carryin => n12894,
            carryout => n12895,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_6_lut_LC_2_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32957\,
            in2 => \_gnd_net_\,
            in3 => \N__23055\,
            lcout => n3197,
            ltout => OPEN,
            carryin => n12895,
            carryout => n12896,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_7_lut_LC_2_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30492\,
            in3 => \N__23052\,
            lcout => n3196,
            ltout => OPEN,
            carryin => n12896,
            carryout => n12897,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_8_lut_LC_2_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54582\,
            in2 => \N__28007\,
            in3 => \N__23049\,
            lcout => n3195,
            ltout => OPEN,
            carryin => n12897,
            carryout => n12898,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_9_lut_LC_2_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27733\,
            in2 => \N__54879\,
            in3 => \N__23046\,
            lcout => n3194,
            ltout => OPEN,
            carryin => n12898,
            carryout => n12899,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_10_lut_LC_2_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54556\,
            in2 => \N__32916\,
            in3 => \N__23043\,
            lcout => n3193,
            ltout => OPEN,
            carryin => \bfn_2_30_0_\,
            carryout => n12900,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_11_lut_LC_2_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54564\,
            in2 => \N__27764\,
            in3 => \N__23040\,
            lcout => n3192,
            ltout => OPEN,
            carryin => n12900,
            carryout => n12901,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_12_lut_LC_2_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54557\,
            in2 => \N__30812\,
            in3 => \N__23037\,
            lcout => n3191,
            ltout => OPEN,
            carryin => n12901,
            carryout => n12902,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_13_lut_LC_2_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54565\,
            in2 => \N__27551\,
            in3 => \N__23034\,
            lcout => n3190,
            ltout => OPEN,
            carryin => n12902,
            carryout => n12903,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_14_lut_LC_2_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30692\,
            in2 => \N__54877\,
            in3 => \N__23103\,
            lcout => n3189,
            ltout => OPEN,
            carryin => n12903,
            carryout => n12904,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_15_lut_LC_2_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27809\,
            in2 => \N__54875\,
            in3 => \N__23100\,
            lcout => n3188,
            ltout => OPEN,
            carryin => n12904,
            carryout => n12905,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_16_lut_LC_2_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23097\,
            in2 => \N__54878\,
            in3 => \N__23079\,
            lcout => n3187,
            ltout => OPEN,
            carryin => n12905,
            carryout => n12906,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_17_lut_LC_2_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27683\,
            in2 => \N__54876\,
            in3 => \N__23076\,
            lcout => n3186,
            ltout => OPEN,
            carryin => n12906,
            carryout => n12907,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_18_lut_LC_2_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30890\,
            in2 => \N__54871\,
            in3 => \N__23073\,
            lcout => n3185,
            ltout => OPEN,
            carryin => \bfn_2_31_0_\,
            carryout => n12908,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_19_lut_LC_2_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27969\,
            in2 => \N__54726\,
            in3 => \N__23070\,
            lcout => n3184,
            ltout => OPEN,
            carryin => n12908,
            carryout => n12909,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_20_lut_LC_2_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30665\,
            in2 => \N__54872\,
            in3 => \N__23067\,
            lcout => n3183,
            ltout => OPEN,
            carryin => n12909,
            carryout => n12910,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_21_lut_LC_2_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30038\,
            in2 => \N__54727\,
            in3 => \N__23064\,
            lcout => n3182,
            ltout => OPEN,
            carryin => n12910,
            carryout => n12911,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_22_lut_LC_2_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27914\,
            in2 => \N__54873\,
            in3 => \N__23061\,
            lcout => n3181,
            ltout => OPEN,
            carryin => n12911,
            carryout => n12912,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_23_lut_LC_2_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27882\,
            in2 => \N__54728\,
            in3 => \N__23130\,
            lcout => n3180,
            ltout => OPEN,
            carryin => n12912,
            carryout => n12913,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_24_lut_LC_2_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30738\,
            in2 => \N__54874\,
            in3 => \N__23127\,
            lcout => n3179,
            ltout => OPEN,
            carryin => n12913,
            carryout => n12914,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_25_lut_LC_2_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31064\,
            in2 => \N__54729\,
            in3 => \N__23124\,
            lcout => n3178,
            ltout => OPEN,
            carryin => n12914,
            carryout => n12915,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_26_lut_LC_2_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31028\,
            in2 => \N__54325\,
            in3 => \N__23121\,
            lcout => n3177,
            ltout => OPEN,
            carryin => \bfn_2_32_0_\,
            carryout => n12916,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_27_lut_LC_2_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30852\,
            in2 => \N__54328\,
            in3 => \N__23118\,
            lcout => n3176,
            ltout => OPEN,
            carryin => n12916,
            carryout => n12917,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_28_lut_LC_2_32_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27843\,
            in2 => \N__54326\,
            in3 => \N__23115\,
            lcout => n3175,
            ltout => OPEN,
            carryin => n12917,
            carryout => n12918,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_29_lut_LC_2_32_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28076\,
            in2 => \N__54329\,
            in3 => \N__23112\,
            lcout => n3174,
            ltout => OPEN,
            carryin => n12918,
            carryout => n12919,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_30_lut_LC_2_32_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28058\,
            in2 => \N__54327\,
            in3 => \N__23109\,
            lcout => n3173,
            ltout => OPEN,
            carryin => n12919,
            carryout => n12920,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2106_31_lut_LC_2_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__53935\,
            in1 => \N__28040\,
            in2 => \N__34940\,
            in3 => \N__23106\,
            lcout => n3204,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_2_lut_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38206\,
            in2 => \_gnd_net_\,
            in3 => \N__23157\,
            lcout => n2301,
            ltout => OPEN,
            carryin => \bfn_3_14_0_\,
            carryout => n12676,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_3_lut_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55543\,
            in2 => \N__23238\,
            in3 => \N__23154\,
            lcout => n2300,
            ltout => OPEN,
            carryin => n12676,
            carryout => n12677,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_4_lut_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25235\,
            in3 => \N__23151\,
            lcout => n2299,
            ltout => OPEN,
            carryin => n12677,
            carryout => n12678,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_5_lut_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55544\,
            in2 => \N__25208\,
            in3 => \N__23148\,
            lcout => n2298,
            ltout => OPEN,
            carryin => n12678,
            carryout => n12679,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_6_lut_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28386\,
            in3 => \N__23145\,
            lcout => n2297,
            ltout => OPEN,
            carryin => n12679,
            carryout => n12680,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_7_lut_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25152\,
            in3 => \N__23142\,
            lcout => n2296,
            ltout => OPEN,
            carryin => n12680,
            carryout => n12681,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_8_lut_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55546\,
            in2 => \N__25400\,
            in3 => \N__23139\,
            lcout => n2295,
            ltout => OPEN,
            carryin => n12681,
            carryout => n12682,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_9_lut_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55545\,
            in2 => \N__28254\,
            in3 => \N__23136\,
            lcout => n2294,
            ltout => OPEN,
            carryin => n12682,
            carryout => n12683,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_10_lut_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55540\,
            in2 => \N__25376\,
            in3 => \N__23133\,
            lcout => n2293,
            ltout => OPEN,
            carryin => \bfn_3_15_0_\,
            carryout => n12684,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_11_lut_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55419\,
            in2 => \N__25349\,
            in3 => \N__23184\,
            lcout => n2292,
            ltout => OPEN,
            carryin => n12684,
            carryout => n12685,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_12_lut_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55541\,
            in2 => \N__28305\,
            in3 => \N__23181\,
            lcout => n2291,
            ltout => OPEN,
            carryin => n12685,
            carryout => n12686,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_13_lut_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55420\,
            in2 => \N__28341\,
            in3 => \N__23178\,
            lcout => n2290,
            ltout => OPEN,
            carryin => n12686,
            carryout => n12687,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_14_lut_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55542\,
            in2 => \N__23310\,
            in3 => \N__23175\,
            lcout => n2289,
            ltout => OPEN,
            carryin => n12687,
            carryout => n12688,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_15_lut_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55421\,
            in2 => \N__25178\,
            in3 => \N__23172\,
            lcout => n2288,
            ltout => OPEN,
            carryin => n12688,
            carryout => n12689,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_16_lut_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25494\,
            in2 => \N__55534\,
            in3 => \N__23169\,
            lcout => n2287,
            ltout => OPEN,
            carryin => n12689,
            carryout => n12690,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_17_lut_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55425\,
            in2 => \N__23349\,
            in3 => \N__23166\,
            lcout => n2286,
            ltout => OPEN,
            carryin => n12690,
            carryout => n12691,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_18_lut_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54732\,
            in2 => \N__25539\,
            in3 => \N__23163\,
            lcout => n2285,
            ltout => OPEN,
            carryin => \bfn_3_16_0_\,
            carryout => n12692,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_19_lut_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54736\,
            in2 => \N__28539\,
            in3 => \N__23160\,
            lcout => n2284,
            ltout => OPEN,
            carryin => n12692,
            carryout => n12693,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_20_lut_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30992\,
            in2 => \N__55035\,
            in3 => \N__23247\,
            lcout => n2283,
            ltout => OPEN,
            carryin => n12693,
            carryout => n12694,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_21_lut_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28488\,
            in2 => \N__55034\,
            in3 => \N__23244\,
            lcout => n2282,
            ltout => OPEN,
            carryin => n12694,
            carryout => n12695,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1503_22_lut_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__25578\,
            in1 => \N__35612\,
            in2 => \N__55036\,
            in3 => \N__23241\,
            lcout => n2313,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10000_4_lut_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__25201\,
            in1 => \N__38210\,
            in2 => \N__23234\,
            in3 => \N__25231\,
            lcout => n11977,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1457_3_lut_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33633\,
            in1 => \N__25317\,
            in2 => \_gnd_net_\,
            in3 => \N__35447\,
            lcout => n2233,
            ltout => \n2233_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1524_3_lut_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23217\,
            in2 => \N__23208\,
            in3 => \N__35574\,
            lcout => n2332,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1523_3_lut_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__25236\,
            in1 => \N__23205\,
            in2 => \N__35595\,
            in3 => \_gnd_net_\,
            lcout => n2331,
            ltout => \n2331_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9994_4_lut_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__38345\,
            in1 => \N__29104\,
            in2 => \N__23196\,
            in3 => \N__28720\,
            lcout => n11971,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1525_3_lut_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__23193\,
            in1 => \N__38211\,
            in2 => \N__35594\,
            in3 => \_gnd_net_\,
            lcout => n2333,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_38_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28336\,
            in1 => \N__23303\,
            in2 => \N__25177\,
            in3 => \N__25323\,
            lcout => n14594,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13018_1_lut_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35596\,
            in3 => \_gnd_net_\,
            lcout => n15748,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1446_3_lut_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25440\,
            in2 => \N__31200\,
            in3 => \N__35436\,
            lcout => n2222,
            ltout => \n2222_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1513_3_lut_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__35538\,
            in1 => \_gnd_net_\,
            in2 => \N__23292\,
            in3 => \N__23289\,
            lcout => n2321,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1515_3_lut_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23280\,
            in2 => \N__28304\,
            in3 => \N__35537\,
            lcout => n2323,
            ltout => \n2323_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_42_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28849\,
            in1 => \N__25636\,
            in2 => \N__23271\,
            in3 => \N__28774\,
            lcout => n14382,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1443_3_lut_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25416\,
            in2 => \N__33114\,
            in3 => \N__35437\,
            lcout => n2219,
            ltout => \n2219_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1510_3_lut_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__35539\,
            in1 => \_gnd_net_\,
            in2 => \N__23268\,
            in3 => \N__23265\,
            lcout => n2318,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1514_3_lut_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23256\,
            in2 => \N__28340\,
            in3 => \N__35533\,
            lcout => n2322,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1517_3_lut_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25377\,
            in2 => \N__35573\,
            in3 => \N__23406\,
            lcout => n2325,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1522_3_lut_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__23397\,
            in1 => \_gnd_net_\,
            in2 => \N__35588\,
            in3 => \N__25212\,
            lcout => n2330,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1519_rep_17_3_lut_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23388\,
            in2 => \N__25404\,
            in3 => \N__35554\,
            lcout => n2327,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1520_3_lut_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__25151\,
            in1 => \_gnd_net_\,
            in2 => \N__35587\,
            in3 => \N__23379\,
            lcout => n2328,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_39_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25150\,
            in2 => \_gnd_net_\,
            in3 => \N__28384\,
            lcout => OPEN,
            ltout => \n14808_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_40_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__25486\,
            in1 => \N__23370\,
            in2 => \N__23361\,
            in3 => \N__23358\,
            lcout => OPEN,
            ltout => \n14598_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_41_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25529\,
            in1 => \N__23342\,
            in2 => \N__23331\,
            in3 => \N__28531\,
            lcout => OPEN,
            ltout => \n14604_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13021_4_lut_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30985\,
            in1 => \N__28484\,
            in2 => \N__23328\,
            in3 => \N__25574\,
            lcout => n2247,
            ltout => \n2247_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1521_3_lut_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28385\,
            in2 => \N__23325\,
            in3 => \N__23322\,
            lcout => n2329,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1512_3_lut_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23523\,
            in2 => \N__25185\,
            in3 => \N__35561\,
            lcout => n2320,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12484_3_lut_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23514\,
            in2 => \N__23462\,
            in3 => \N__35716\,
            lcout => n2423,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1511_3_lut_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23505\,
            in1 => \N__25490\,
            in2 => \_gnd_net_\,
            in3 => \N__35562\,
            lcout => n2319,
            ltout => \n2319_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1578_3_lut_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23496\,
            in2 => \N__23487\,
            in3 => \N__35717\,
            lcout => n2418,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_46_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__25894\,
            in1 => \N__23484\,
            in2 => \N__28831\,
            in3 => \N__23412\,
            lcout => n14392,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12483_3_lut_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__23475\,
            in1 => \N__25353\,
            in2 => \N__35589\,
            in3 => \_gnd_net_\,
            lcout => n2324,
            ltout => \n2324_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_43_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25864\,
            in1 => \N__25774\,
            in2 => \N__23442\,
            in3 => \N__28681\,
            lcout => OPEN,
            ltout => \n14384_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_45_LC_3_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25618\,
            in1 => \N__23435\,
            in2 => \N__23424\,
            in3 => \N__23421\,
            lcout => n14390,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1718_3_lut_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__32499\,
            in1 => \_gnd_net_\,
            in2 => \N__36102\,
            in3 => \N__32513\,
            lcout => n2622,
            ltout => \n2622_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1785_3_lut_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23772\,
            in2 => \N__23760\,
            in3 => \N__36268\,
            lcout => n2721,
            ltout => \n2721_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_55_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23726\,
            in1 => \N__23708\,
            in2 => \N__23697\,
            in3 => \N__23620\,
            lcout => n14348,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1719_3_lut_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32070\,
            in2 => \N__32090\,
            in3 => \N__36094\,
            lcout => n2623,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1575_3_lut_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__23685\,
            in1 => \_gnd_net_\,
            in2 => \N__35745\,
            in3 => \N__25727\,
            lcout => n2415,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1724_3_lut_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__32244\,
            in1 => \_gnd_net_\,
            in2 => \N__32217\,
            in3 => \N__36090\,
            lcout => n2628,
            ltout => \n2628_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_32_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26017\,
            in1 => \N__23666\,
            in2 => \N__23655\,
            in3 => \N__33907\,
            lcout => n14668,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1788_3_lut_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36267\,
            in2 => \N__25964\,
            in3 => \N__23652\,
            lcout => n2724,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1791_3_lut_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23604\,
            in2 => \N__23582\,
            in3 => \N__36224\,
            lcout => n2727,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1796_3_lut_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23538\,
            in2 => \N__36276\,
            in3 => \N__26261\,
            lcout => n2732,
            ltout => \n2732_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9980_3_lut_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26614\,
            in2 => \N__23919\,
            in3 => \N__33523\,
            lcout => OPEN,
            ltout => \n11957_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_58_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__23905\,
            in1 => \N__23827\,
            in2 => \N__23889\,
            in3 => \N__24352\,
            lcout => n13808,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_50_LC_3_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29383\,
            in1 => \N__23870\,
            in2 => \N__26231\,
            in3 => \N__23859\,
            lcout => n14674,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1794_3_lut_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29195\,
            in2 => \N__36277\,
            in3 => \N__23853\,
            lcout => n2730,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1795_3_lut_LC_3_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__23811\,
            in1 => \_gnd_net_\,
            in2 => \N__36278\,
            in3 => \N__29252\,
            lcout => n2731,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1797_3_lut_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33577\,
            in1 => \N__23796\,
            in2 => \_gnd_net_\,
            in3 => \N__36240\,
            lcout => n2733,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_28_LC_3_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__26134\,
            in1 => \N__24124\,
            in2 => \N__26244\,
            in3 => \N__25827\,
            lcout => OPEN,
            ltout => \n14650_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_31_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29683\,
            in1 => \N__32617\,
            in2 => \N__23778\,
            in3 => \N__25932\,
            lcout => OPEN,
            ltout => \n14654_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_34_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26164\,
            in1 => \N__26191\,
            in2 => \N__23775\,
            in3 => \N__29533\,
            lcout => OPEN,
            ltout => \n14660_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12565_4_lut_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32548\,
            in1 => \N__32722\,
            in2 => \N__24189\,
            in3 => \N__24186\,
            lcout => n2643,
            ltout => \n2643_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1782_3_lut_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__26135\,
            in1 => \_gnd_net_\,
            in2 => \N__24180\,
            in3 => \N__24177\,
            lcout => n2718,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1786_3_lut_LC_3_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24144\,
            in2 => \N__24129\,
            in3 => \N__36241\,
            lcout => n2722,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1863_3_lut_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24074\,
            in2 => \N__24054\,
            in3 => \N__36427\,
            lcout => n2831,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1842_3_lut_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__24035\,
            in1 => \_gnd_net_\,
            in2 => \N__36455\,
            in3 => \N__24021\,
            lcout => n2810,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1850_3_lut_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24003\,
            in2 => \N__23991\,
            in3 => \N__36429\,
            lcout => n2818,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1781_3_lut_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__26230\,
            in1 => \_gnd_net_\,
            in2 => \N__36281\,
            in3 => \N__23967\,
            lcout => n2717,
            ltout => \n2717_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1848_3_lut_LC_3_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23934\,
            in2 => \N__23922\,
            in3 => \N__36430\,
            lcout => n2816,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1844_3_lut_LC_3_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24416\,
            in2 => \N__36454\,
            in3 => \N__24393\,
            lcout => n2812,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1862_3_lut_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24381\,
            in2 => \N__24368\,
            in3 => \N__36428\,
            lcout => n2830,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1776_3_lut_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26168\,
            in2 => \N__36282\,
            in3 => \N__24336\,
            lcout => n2712,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1919_3_lut_LC_3_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__24308\,
            in1 => \N__24321\,
            in2 => \N__34323\,
            in3 => \_gnd_net_\,
            lcout => n2919,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_62_LC_3_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24616\,
            in1 => \N__29329\,
            in2 => \N__26750\,
            in3 => \N__29827\,
            lcout => OPEN,
            ltout => \n14690_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_63_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24307\,
            in1 => \N__26833\,
            in2 => \N__24294\,
            in3 => \N__24291\,
            lcout => OPEN,
            ltout => \n14696_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_65_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27239\,
            in1 => \N__26281\,
            in2 => \N__24282\,
            in3 => \N__26514\,
            lcout => n14702,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1845_3_lut_LC_3_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24277\,
            in2 => \N__24246\,
            in3 => \N__36410\,
            lcout => n2813,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1851_3_lut_LC_3_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24231\,
            in2 => \N__24204\,
            in3 => \N__36409\,
            lcout => n2819,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1922_3_lut_LC_3_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__24617\,
            in1 => \_gnd_net_\,
            in2 => \N__24603\,
            in3 => \N__34293\,
            lcout => n2922,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1926_3_lut_LC_3_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24588\,
            in2 => \N__24561\,
            in3 => \N__34277\,
            lcout => n2926,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1921_3_lut_LC_3_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24546\,
            in2 => \N__24519\,
            in3 => \N__34278\,
            lcout => n2921,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1982_3_lut_LC_3_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27118\,
            in2 => \N__24504\,
            in3 => \N__34461\,
            lcout => n3014,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1986_3_lut_LC_3_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26655\,
            in2 => \N__24495\,
            in3 => \N__34460\,
            lcout => n3018,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i16_1_lut_LC_3_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46500\,
            lcout => n10_adj_582,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1911_3_lut_LC_3_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26472\,
            in2 => \N__34320\,
            in3 => \N__24486\,
            lcout => n2911,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1841_3_lut_LC_3_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24471\,
            in2 => \N__24444\,
            in3 => \N__36458\,
            lcout => n2809,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1996_3_lut_LC_3_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24426\,
            in2 => \N__27168\,
            in3 => \N__34453\,
            lcout => n3028,
            ltout => \n3028_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2063_3_lut_LC_3_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__24813\,
            in1 => \_gnd_net_\,
            in2 => \N__24672\,
            in3 => \N__34603\,
            lcout => n3127,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1988_3_lut_LC_3_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26700\,
            in2 => \N__24669\,
            in3 => \N__34454\,
            lcout => n3020,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1912_3_lut_LC_3_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24660\,
            in2 => \N__26448\,
            in3 => \N__34332\,
            lcout => n2912,
            ltout => \n2912_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1979_3_lut_LC_3_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__24648\,
            in1 => \_gnd_net_\,
            in2 => \N__24642\,
            in3 => \N__34459\,
            lcout => n3011,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12654_1_lut_LC_3_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34502\,
            in3 => \_gnd_net_\,
            lcout => n15384,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1983_3_lut_LC_3_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27200\,
            in2 => \N__24639\,
            in3 => \N__34458\,
            lcout => n3015,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_2_lut_LC_3_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41570\,
            in2 => \_gnd_net_\,
            in3 => \N__24630\,
            lcout => n3101,
            ltout => OPEN,
            carryin => \bfn_3_28_0_\,
            carryout => n12864,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_3_lut_LC_3_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54443\,
            in2 => \N__30099\,
            in3 => \N__24627\,
            lcout => n3100,
            ltout => OPEN,
            carryin => n12864,
            carryout => n12865,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_4_lut_LC_3_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30078\,
            in3 => \N__24624\,
            lcout => n3099,
            ltout => OPEN,
            carryin => n12865,
            carryout => n12866,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_5_lut_LC_3_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54444\,
            in2 => \N__29931\,
            in3 => \N__24849\,
            lcout => n3098,
            ltout => OPEN,
            carryin => n12866,
            carryout => n12867,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_6_lut_LC_3_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29979\,
            in3 => \N__24846\,
            lcout => n3097,
            ltout => OPEN,
            carryin => n12867,
            carryout => n12868,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_7_lut_LC_3_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29954\,
            in3 => \N__24834\,
            lcout => n3096,
            ltout => OPEN,
            carryin => n12868,
            carryout => n12869,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_8_lut_LC_3_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54446\,
            in2 => \N__24831\,
            in3 => \N__24807\,
            lcout => n3095,
            ltout => OPEN,
            carryin => n12869,
            carryout => n12870,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_9_lut_LC_3_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54445\,
            in2 => \N__30587\,
            in3 => \N__24795\,
            lcout => n3094,
            ltout => OPEN,
            carryin => n12870,
            carryout => n12871,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_10_lut_LC_3_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54574\,
            in2 => \N__24792\,
            in3 => \N__24753\,
            lcout => n3093,
            ltout => OPEN,
            carryin => \bfn_3_29_0_\,
            carryout => n12872,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_11_lut_LC_3_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54578\,
            in2 => \N__24750\,
            in3 => \N__24714\,
            lcout => n3092,
            ltout => OPEN,
            carryin => n12872,
            carryout => n12873,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_12_lut_LC_3_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54575\,
            in2 => \N__24711\,
            in3 => \N__24675\,
            lcout => n3091,
            ltout => OPEN,
            carryin => n12873,
            carryout => n12874,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_13_lut_LC_3_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54579\,
            in2 => \N__30561\,
            in3 => \N__25020\,
            lcout => n3090,
            ltout => OPEN,
            carryin => n12874,
            carryout => n12875,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_14_lut_LC_3_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54576\,
            in2 => \N__25017\,
            in3 => \N__24981\,
            lcout => n3089,
            ltout => OPEN,
            carryin => n12875,
            carryout => n12876,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_15_lut_LC_3_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54580\,
            in2 => \N__24977\,
            in3 => \N__24942\,
            lcout => n3088,
            ltout => OPEN,
            carryin => n12876,
            carryout => n12877,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_16_lut_LC_3_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54577\,
            in2 => \N__24939\,
            in3 => \N__24906\,
            lcout => n3087,
            ltout => OPEN,
            carryin => n12877,
            carryout => n12878,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_17_lut_LC_3_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54581\,
            in2 => \N__30624\,
            in3 => \N__24894\,
            lcout => n3086,
            ltout => OPEN,
            carryin => n12878,
            carryout => n12879,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_18_lut_LC_3_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27282\,
            in2 => \N__54864\,
            in3 => \N__24891\,
            lcout => n3085,
            ltout => OPEN,
            carryin => \bfn_3_30_0_\,
            carryout => n12880,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_19_lut_LC_3_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24888\,
            in2 => \N__54868\,
            in3 => \N__24855\,
            lcout => n3084,
            ltout => OPEN,
            carryin => n12880,
            carryout => n12881,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_20_lut_LC_3_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30323\,
            in2 => \N__54865\,
            in3 => \N__24852\,
            lcout => n3083,
            ltout => OPEN,
            carryin => n12881,
            carryout => n12882,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_21_lut_LC_3_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27494\,
            in2 => \N__54869\,
            in3 => \N__25062\,
            lcout => n3082,
            ltout => OPEN,
            carryin => n12882,
            carryout => n12883,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_22_lut_LC_3_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27462\,
            in2 => \N__54866\,
            in3 => \N__25059\,
            lcout => n3081,
            ltout => OPEN,
            carryin => n12883,
            carryout => n12884,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_23_lut_LC_3_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27587\,
            in2 => \N__54870\,
            in3 => \N__25056\,
            lcout => n3080,
            ltout => OPEN,
            carryin => n12884,
            carryout => n12885,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_24_lut_LC_3_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30251\,
            in2 => \N__54867\,
            in3 => \N__25053\,
            lcout => n3079,
            ltout => OPEN,
            carryin => n12885,
            carryout => n12886,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_25_lut_LC_3_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54534\,
            in2 => \N__27431\,
            in3 => \N__25050\,
            lcout => n3078,
            ltout => OPEN,
            carryin => n12886,
            carryout => n12887,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_26_lut_LC_3_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28208\,
            in2 => \N__54860\,
            in3 => \N__25047\,
            lcout => n3077,
            ltout => OPEN,
            carryin => \bfn_3_31_0_\,
            carryout => n12888,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_27_lut_LC_3_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27404\,
            in2 => \N__54862\,
            in3 => \N__25044\,
            lcout => n3076,
            ltout => OPEN,
            carryin => n12888,
            carryout => n12889,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_28_lut_LC_3_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27347\,
            in2 => \N__54861\,
            in3 => \N__25041\,
            lcout => n3075,
            ltout => OPEN,
            carryin => n12889,
            carryout => n12890,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_29_lut_LC_3_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27323\,
            in2 => \N__54863\,
            in3 => \N__25038\,
            lcout => n3074,
            ltout => OPEN,
            carryin => n12890,
            carryout => n12891,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2039_30_lut_LC_3_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__54515\,
            in1 => \N__34739\,
            in2 => \N__27369\,
            in3 => \N__25128\,
            lcout => n3105,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2043_3_lut_LC_3_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__27348\,
            in1 => \_gnd_net_\,
            in2 => \N__25125\,
            in3 => \N__34664\,
            lcout => n3107,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2050_3_lut_LC_3_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25116\,
            in2 => \N__34697\,
            in3 => \N__27498\,
            lcout => n3114,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2042_3_lut_LC_3_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27324\,
            in2 => \N__25110\,
            in3 => \N__34665\,
            lcout => n3106,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2109_3_lut_LC_3_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28059\,
            in2 => \N__34906\,
            in3 => \N__25101\,
            lcout => n3205,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12721_1_lut_LC_3_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34858\,
            lcout => n15451,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2110_3_lut_LC_3_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25095\,
            in2 => \N__34907\,
            in3 => \N__28077\,
            lcout => n3206,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2047_3_lut_LC_3_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25089\,
            in2 => \N__30258\,
            in3 => \N__34698\,
            lcout => n3111,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2046_3_lut_LC_3_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27432\,
            in2 => \N__25080\,
            in3 => \N__34699\,
            lcout => n3110,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2044_3_lut_LC_3_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25068\,
            in2 => \N__34714\,
            in3 => \N__27405\,
            lcout => n3108,
            ltout => \n3108_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2111_3_lut_LC_3_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25245\,
            in2 => \N__25239\,
            in3 => \N__34862\,
            lcout => n3207,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1456_3_lut_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25308\,
            in2 => \N__35446\,
            in3 => \N__33677\,
            lcout => n2232,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1455_3_lut_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25296\,
            in2 => \N__35445\,
            in3 => \N__33705\,
            lcout => n2231,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_33_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__28097\,
            in1 => \N__28150\,
            in2 => \N__25271\,
            in3 => \N__33645\,
            lcout => n13787,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1450_3_lut_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__25467\,
            in1 => \_gnd_net_\,
            in2 => \N__28128\,
            in3 => \N__35419\,
            lcout => n2226,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1445_3_lut_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28455\,
            in2 => \N__35444\,
            in3 => \N__25431\,
            lcout => n2221,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1449_rep_20_3_lut_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25458\,
            in2 => \N__28611\,
            in3 => \N__35418\,
            lcout => n2225,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1453_3_lut_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25281\,
            in2 => \N__35443\,
            in3 => \N__28151\,
            lcout => n2229,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1385_3_lut_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33777\,
            in2 => \N__31170\,
            in3 => \N__35298\,
            lcout => n2129,
            ltout => \n2129_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1452_3_lut_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__35420\,
            in1 => \_gnd_net_\,
            in2 => \N__25407\,
            in3 => \N__25254\,
            lcout => n2228,
            ltout => \n2228_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_37_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25369\,
            in1 => \N__25342\,
            in2 => \N__25326\,
            in3 => \N__28356\,
            lcout => n14588,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_2_lut_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33632\,
            in2 => \_gnd_net_\,
            in3 => \N__25311\,
            lcout => n2201,
            ltout => OPEN,
            carryin => \bfn_4_17_0_\,
            carryout => n12657,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_3_lut_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55453\,
            in2 => \N__33678\,
            in3 => \N__25299\,
            lcout => n2200,
            ltout => OPEN,
            carryin => n12657,
            carryout => n12658,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_4_lut_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33704\,
            in3 => \N__25287\,
            lcout => n2199,
            ltout => OPEN,
            carryin => n12658,
            carryout => n12659,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_5_lut_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55454\,
            in2 => \N__28101\,
            in3 => \N__25284\,
            lcout => n2198,
            ltout => OPEN,
            carryin => n12659,
            carryout => n12660,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_6_lut_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28155\,
            in3 => \N__25275\,
            lcout => n2197,
            ltout => OPEN,
            carryin => n12660,
            carryout => n12661,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_7_lut_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25272\,
            in3 => \N__25248\,
            lcout => n2196,
            ltout => OPEN,
            carryin => n12661,
            carryout => n12662,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_8_lut_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54351\,
            in2 => \N__28224\,
            in3 => \N__25470\,
            lcout => n2195,
            ltout => OPEN,
            carryin => n12662,
            carryout => n12663,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_9_lut_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55455\,
            in2 => \N__28127\,
            in3 => \N__25461\,
            lcout => n2194,
            ltout => OPEN,
            carryin => n12663,
            carryout => n12664,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_10_lut_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55444\,
            in2 => \N__28607\,
            in3 => \N__25449\,
            lcout => n2193,
            ltout => OPEN,
            carryin => \bfn_4_18_0_\,
            carryout => n12665,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_11_lut_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54346\,
            in2 => \N__28574\,
            in3 => \N__25446\,
            lcout => n2192,
            ltout => OPEN,
            carryin => n12665,
            carryout => n12666,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_12_lut_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55445\,
            in2 => \N__28425\,
            in3 => \N__25443\,
            lcout => n2191,
            ltout => OPEN,
            carryin => n12666,
            carryout => n12667,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_13_lut_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54347\,
            in2 => \N__31199\,
            in3 => \N__25434\,
            lcout => n2190,
            ltout => OPEN,
            carryin => n12667,
            carryout => n12668,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_14_lut_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55446\,
            in2 => \N__28451\,
            in3 => \N__25422\,
            lcout => n2189,
            ltout => OPEN,
            carryin => n12668,
            carryout => n12669,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_15_lut_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31313\,
            in2 => \N__55538\,
            in3 => \N__25419\,
            lcout => n2188,
            ltout => OPEN,
            carryin => n12669,
            carryout => n12670,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_16_lut_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33110\,
            in2 => \N__54731\,
            in3 => \N__25410\,
            lcout => n2187,
            ltout => OPEN,
            carryin => n12670,
            carryout => n12671,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_17_lut_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33227\,
            in2 => \N__55539\,
            in3 => \N__25593\,
            lcout => n2186,
            ltout => OPEN,
            carryin => n12671,
            carryout => n12672,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_18_lut_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28891\,
            in2 => \N__55536\,
            in3 => \N__25590\,
            lcout => n2185,
            ltout => OPEN,
            carryin => \bfn_4_19_0_\,
            carryout => n12673,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_19_lut_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31355\,
            in2 => \N__54730\,
            in3 => \N__25587\,
            lcout => n2184,
            ltout => OPEN,
            carryin => n12673,
            carryout => n12674,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_20_lut_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28499\,
            in2 => \N__55537\,
            in3 => \N__25584\,
            lcout => n2183,
            ltout => OPEN,
            carryin => n12674,
            carryout => n12675,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1436_21_lut_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__54345\,
            in1 => \N__35462\,
            in2 => \N__31224\,
            in3 => \N__25581\,
            lcout => n2214,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1518_3_lut_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__28246\,
            in1 => \_gnd_net_\,
            in2 => \N__25563\,
            in3 => \N__35540\,
            lcout => n2326,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1442_3_lut_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33228\,
            in2 => \N__25548\,
            in3 => \N__35417\,
            lcout => n2218,
            ltout => \n2218_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1509_3_lut_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__25518\,
            in1 => \_gnd_net_\,
            in2 => \N__25506\,
            in3 => \N__35541\,
            lcout => n2317,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1444_3_lut_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31314\,
            in2 => \N__25503\,
            in3 => \N__35416\,
            lcout => n2220,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_47_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25723\,
            in1 => \N__28972\,
            in2 => \N__29017\,
            in3 => \N__25818\,
            lcout => OPEN,
            ltout => \n14398_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13048_4_lut_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25805\,
            in1 => \N__30952\,
            in2 => \N__25785\,
            in3 => \N__25688\,
            lcout => n2346,
            ltout => \n2346_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12485_3_lut_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__25778\,
            in1 => \_gnd_net_\,
            in2 => \N__25758\,
            in3 => \N__25755\,
            lcout => n2426,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1508_3_lut_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25743\,
            in2 => \N__28535\,
            in3 => \N__35566\,
            lcout => n2316,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1506_3_lut_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25707\,
            in2 => \N__35590\,
            in3 => \N__28483\,
            lcout => n2314,
            ltout => \n2314_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1573_3_lut_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__35708\,
            in1 => \_gnd_net_\,
            in2 => \N__25677\,
            in3 => \N__25674\,
            lcout => n2413,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1584_3_lut_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25662\,
            in2 => \N__25652\,
            in3 => \N__35704\,
            lcout => n2424,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1579_3_lut_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25622\,
            in2 => \N__35740\,
            in3 => \N__25602\,
            lcout => n2419,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1574_3_lut_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__25926\,
            in1 => \_gnd_net_\,
            in2 => \N__35742\,
            in3 => \N__30962\,
            lcout => n2414,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1588_3_lut_LC_4_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25917\,
            in2 => \N__25905\,
            in3 => \N__35709\,
            lcout => n2428,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1587_3_lut_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25874\,
            in2 => \N__35741\,
            in3 => \N__25848\,
            lcout => n2427,
            ltout => \n2427_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_48_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33968\,
            in1 => \N__31798\,
            in2 => \N__25836\,
            in3 => \N__31420\,
            lcout => OPEN,
            ltout => \n14620_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_49_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31498\,
            in2 => \N__25833\,
            in3 => \N__34102\,
            lcout => n14622,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1654_3_lut_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31464\,
            in2 => \N__31449\,
            in3 => \N__35911\,
            lcout => n2526,
            ltout => \n2526_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1721_3_lut_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32109\,
            in2 => \N__25830\,
            in3 => \N__36097\,
            lcout => n2625,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29438\,
            in3 => \N__29500\,
            lcout => n14816,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1647_3_lut_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31710\,
            in2 => \N__31728\,
            in3 => \N__35862\,
            lcout => n2519,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1652_3_lut_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31404\,
            in2 => \N__35898\,
            in3 => \N__31430\,
            lcout => n2524,
            ltout => \n2524_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_154_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32189\,
            in2 => \N__26055\,
            in3 => \N__32120\,
            lcout => OPEN,
            ltout => \n14574_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_159_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32404\,
            in1 => \N__26046\,
            in2 => \N__26052\,
            in3 => \N__32661\,
            lcout => n14117,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1651_3_lut_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__31808\,
            in1 => \_gnd_net_\,
            in2 => \N__31785\,
            in3 => \N__35861\,
            lcout => n2523,
            ltout => \n2523_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_156_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32156\,
            in2 => \N__26049\,
            in3 => \N__32446\,
            lcout => n14576,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1655_3_lut_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31502\,
            in2 => \N__31482\,
            in3 => \N__35860\,
            lcout => n2527,
            ltout => \n2527_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1722_3_lut_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32145\,
            in2 => \N__26040\,
            in3 => \N__36068\,
            lcout => n2626,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1713_3_lut_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33840\,
            in2 => \N__32370\,
            in3 => \N__36048\,
            lcout => n2617,
            ltout => \n2617_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_29_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25963\,
            in2 => \N__25935\,
            in3 => \N__29059\,
            lcout => n14812,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1729_3_lut_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35145\,
            in1 => \N__31881\,
            in2 => \_gnd_net_\,
            in3 => \N__36044\,
            lcout => n2633,
            ltout => \n2633_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10082_4_lut_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__29182\,
            in1 => \N__33581\,
            in2 => \N__26247\,
            in3 => \N__29239\,
            lcout => n12059,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1714_3_lut_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32408\,
            in2 => \N__32388\,
            in3 => \N__36049\,
            lcout => n2618,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1710_3_lut_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__32858\,
            in1 => \_gnd_net_\,
            in2 => \N__36086\,
            in3 => \N__32844\,
            lcout => n2614,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1709_3_lut_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32822\,
            in2 => \N__32802\,
            in3 => \N__36050\,
            lcout => n2613,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1715_3_lut_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__32450\,
            in1 => \_gnd_net_\,
            in2 => \N__36085\,
            in3 => \N__32430\,
            lcout => n2619,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1929_3_lut_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26118\,
            in2 => \N__26540\,
            in3 => \N__34301\,
            lcout => n2929,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1843_3_lut_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26102\,
            in2 => \N__26082\,
            in3 => \N__36426\,
            lcout => n2811,
            ltout => \n2811_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1910_3_lut_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26067\,
            in2 => \N__26058\,
            in3 => \N__34302\,
            lcout => n2910,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1864_3_lut_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26618\,
            in2 => \N__26598\,
            in3 => \N__36425\,
            lcout => n2832,
            ltout => \n2832_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9976_3_lut_LC_4_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33496\,
            in2 => \N__26580\,
            in3 => \N__26573\,
            lcout => OPEN,
            ltout => \n11953_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_64_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__29635\,
            in1 => \N__26533\,
            in2 => \N__26517\,
            in3 => \N__29888\,
            lcout => n13857,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_66_LC_4_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29774\,
            in1 => \N__26332\,
            in2 => \N__26508\,
            in3 => \N__26478\,
            lcout => OPEN,
            ltout => \n14708_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_67_LC_4_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26464\,
            in1 => \N__26434\,
            in2 => \N__26421\,
            in3 => \N__26414\,
            lcout => OPEN,
            ltout => \n14714_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12626_4_lut_LC_4_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26395\,
            in1 => \N__26893\,
            in2 => \N__26370\,
            in3 => \N__26366\,
            lcout => n2841,
            ltout => \n2841_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1915_3_lut_LC_4_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__26333\,
            in1 => \_gnd_net_\,
            in2 => \N__26319\,
            in3 => \N__26316\,
            lcout => n2915,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1917_3_lut_LC_4_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26304\,
            in2 => \N__26291\,
            in3 => \N__34297\,
            lcout => n2917,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2049_3_lut_LC_4_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26913\,
            in2 => \N__27461\,
            in3 => \N__34659\,
            lcout => n3113,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1909_3_lut_LC_4_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__26894\,
            in1 => \_gnd_net_\,
            in2 => \N__34324\,
            in3 => \N__26880\,
            lcout => n2909,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1976_3_lut_LC_4_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__26971\,
            in1 => \_gnd_net_\,
            in2 => \N__26871\,
            in3 => \N__34479\,
            lcout => n3008,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1918_3_lut_LC_4_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__34290\,
            in1 => \N__26856\,
            in2 => \N__26843\,
            in3 => \_gnd_net_\,
            lcout => n2918,
            ltout => \n2918_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_155_LC_4_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26796\,
            in1 => \N__26773\,
            in2 => \N__26757\,
            in3 => \N__29277\,
            lcout => n14216,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1924_3_lut_LC_4_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__34292\,
            in1 => \N__26754\,
            in2 => \N__26715\,
            in3 => \_gnd_net_\,
            lcout => n2924,
            ltout => \n2924_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_69_LC_4_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26698\,
            in1 => \N__26674\,
            in2 => \N__26658\,
            in3 => \N__26653\,
            lcout => OPEN,
            ltout => \n14212_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_161_LC_4_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27196\,
            in1 => \N__30355\,
            in2 => \N__26637\,
            in3 => \N__26634\,
            lcout => n14222,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12622_1_lut_LC_4_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34289\,
            lcout => n15352,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1916_3_lut_LC_4_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34291\,
            in1 => \N__27243\,
            in2 => \_gnd_net_\,
            in3 => \N__27216\,
            lcout => n2916,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1981_3_lut_LC_4_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27092\,
            in2 => \N__27180\,
            in3 => \N__34474\,
            lcout => n3013,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_162_LC_4_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__29590\,
            in1 => \N__30198\,
            in2 => \N__27166\,
            in3 => \N__27129\,
            lcout => OPEN,
            ltout => \n14224_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_163_LC_4_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30286\,
            in1 => \N__27119\,
            in2 => \N__27096\,
            in3 => \N__27091\,
            lcout => OPEN,
            ltout => \n14230_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_164_LC_4_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27064\,
            in1 => \N__26935\,
            in2 => \N__27045\,
            in3 => \N__27041\,
            lcout => OPEN,
            ltout => \n14236_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12658_4_lut_LC_4_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27026\,
            in1 => \N__27003\,
            in2 => \N__26982\,
            in3 => \N__26972\,
            lcout => n2940,
            ltout => \n2940_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1997_3_lut_LC_4_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__29591\,
            in1 => \_gnd_net_\,
            in2 => \N__26952\,
            in3 => \N__26949\,
            lcout => n3029,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1978_3_lut_LC_4_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26936\,
            in1 => \N__34475\,
            in2 => \_gnd_net_\,
            in3 => \N__26922\,
            lcout => n3010,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1995_3_lut_LC_4_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__34473\,
            in1 => \_gnd_net_\,
            in2 => \N__27528\,
            in3 => \N__29852\,
            lcout => n3027,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2000_3_lut_LC_4_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30221\,
            in2 => \N__27513\,
            in3 => \N__34462\,
            lcout => n3032,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_170_LC_4_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27487\,
            in1 => \N__30310\,
            in2 => \N__30528\,
            in3 => \N__27474\,
            lcout => OPEN,
            ltout => \n14742_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_171_LC_4_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30238\,
            in1 => \N__27457\,
            in2 => \N__27435\,
            in3 => \N__27574\,
            lcout => OPEN,
            ltout => \n14748_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_172_LC_4_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27418\,
            in1 => \N__27394\,
            in2 => \N__27372\,
            in3 => \N__28196\,
            lcout => OPEN,
            ltout => \n14754_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12691_4_lut_LC_4_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27365\,
            in1 => \N__27341\,
            in2 => \N__27327\,
            in3 => \N__27311\,
            lcout => n3039,
            ltout => \n3039_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2067_3_lut_LC_4_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27291\,
            in2 => \N__27285\,
            in3 => \N__30077\,
            lcout => n3131,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2053_3_lut_LC_4_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27277\,
            in2 => \N__27252\,
            in3 => \N__34604\,
            lcout => n3117,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2066_3_lut_LC_4_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__34612\,
            in1 => \N__29927\,
            in2 => \N__27633\,
            in3 => \_gnd_net_\,
            lcout => n3130,
            ltout => \n3130_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_177_LC_4_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__30484\,
            in1 => \N__30385\,
            in2 => \N__27624\,
            in3 => \N__27600\,
            lcout => n13831,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2069_3_lut_LC_4_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__27621\,
            in1 => \_gnd_net_\,
            in2 => \N__34657\,
            in3 => \N__41571\,
            lcout => n3133,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2065_3_lut_LC_4_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27615\,
            in2 => \N__29978\,
            in3 => \N__34611\,
            lcout => n3129,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2068_3_lut_LC_4_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30095\,
            in2 => \N__34658\,
            in3 => \N__27609\,
            lcout => n3132,
            ltout => \n3132_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9968_3_lut_LC_4_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34166\,
            in2 => \N__27603\,
            in3 => \N__30421\,
            lcout => n11945,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2048_3_lut_LC_4_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__34613\,
            in1 => \N__27594\,
            in2 => \N__27588\,
            in3 => \_gnd_net_\,
            lcout => n3112,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2195_3_lut_LC_4_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37152\,
            in2 => \N__37172\,
            in3 => \N__35041\,
            lcout => OPEN,
            ltout => \n23_adj_715_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_89_LC_4_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__35045\,
            in1 => \N__36999\,
            in2 => \N__27558\,
            in3 => \N__37019\,
            lcout => n14260,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2126_3_lut_LC_4_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27555\,
            in2 => \N__27825\,
            in3 => \N__34824\,
            lcout => n3222,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2124_3_lut_LC_4_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27813\,
            in2 => \N__34881\,
            in3 => \N__27786\,
            lcout => n3220,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2128_3_lut_LC_4_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27777\,
            in2 => \N__27768\,
            in3 => \N__34823\,
            lcout => n3224,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_90_LC_4_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101100"
        )
    port map (
            in0 => \N__36677\,
            in1 => \N__36663\,
            in2 => \N__35087\,
            in3 => \N__30756\,
            lcout => n14264,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2130_3_lut_LC_4_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27734\,
            in2 => \N__27705\,
            in3 => \N__34825\,
            lcout => n3226,
            ltout => \n3226_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_121_LC_4_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36712\,
            in1 => \N__37165\,
            in2 => \N__27690\,
            in3 => \N__37090\,
            lcout => n14768,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2122_3_lut_LC_4_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27687\,
            in2 => \N__27663\,
            in3 => \N__34876\,
            lcout => n3218,
            ltout => \n3218_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_128_LC_4_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37015\,
            in2 => \N__27648\,
            in3 => \N__36976\,
            lcout => n14798,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2116_3_lut_LC_4_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27881\,
            in2 => \N__27645\,
            in3 => \N__34880\,
            lcout => n3212,
            ltout => \n3212_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_131_LC_4_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37432\,
            in1 => \N__37550\,
            in2 => \N__28086\,
            in3 => \N__28083\,
            lcout => n14804,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12725_4_lut_LC_4_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28075\,
            in1 => \N__28057\,
            in2 => \N__28041\,
            in3 => \N__27831\,
            lcout => n3138,
            ltout => \n3138_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2131_3_lut_LC_4_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28026\,
            in2 => \N__28014\,
            in3 => \N__28011\,
            lcout => n3227,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2117_3_lut_LC_4_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27915\,
            in2 => \N__27990\,
            in3 => \N__34875\,
            lcout => n3213,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2120_3_lut_LC_4_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__27978\,
            in1 => \N__27967\,
            in2 => \N__34910\,
            in3 => \_gnd_net_\,
            lcout => n3216,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2051_3_lut_LC_4_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30324\,
            in2 => \N__27939\,
            in3 => \N__34704\,
            lcout => n3115,
            ltout => \n3115_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_178_LC_4_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27924\,
            in1 => \N__27913\,
            in2 => \N__27897\,
            in3 => \N__27894\,
            lcout => OPEN,
            ltout => \n14162_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_179_LC_4_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30737\,
            in1 => \N__27877\,
            in2 => \N__27849\,
            in3 => \N__31063\,
            lcout => OPEN,
            ltout => \n14168_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_180_LC_4_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30847\,
            in1 => \N__31027\,
            in2 => \N__27846\,
            in3 => \N__27842\,
            lcout => n14174,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2045_3_lut_LC_4_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28209\,
            in2 => \N__28185\,
            in3 => \N__34703\,
            lcout => n3109,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_95_LC_4_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30867\,
            in1 => \N__28176\,
            in2 => \N__28167\,
            in3 => \N__33000\,
            lcout => n14282,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1386_3_lut_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30912\,
            in2 => \N__35302\,
            in3 => \N__33345\,
            lcout => n2130,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_30_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28581\,
            in1 => \N__33103\,
            in2 => \N__31312\,
            in3 => \N__28107\,
            lcout => OPEN,
            ltout => \n14324_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_35_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28895\,
            in1 => \N__33220\,
            in2 => \N__28137\,
            in3 => \N__28134\,
            lcout => n14330,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1383_3_lut_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31143\,
            in2 => \N__35303\,
            in3 => \N__33447\,
            lcout => n2127,
            ltout => \n2127_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28450\,
            in2 => \N__28110\,
            in3 => \N__28573\,
            lcout => n14318,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1387_3_lut_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33369\,
            in2 => \N__30924\,
            in3 => \N__35292\,
            lcout => n2131,
            ltout => \n2131_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1454_3_lut_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__28395\,
            in1 => \_gnd_net_\,
            in2 => \N__28389\,
            in3 => \N__35399\,
            lcout => n2230,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_36_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28247\,
            in3 => \N__28288\,
            lcout => n14584,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1447_3_lut_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28421\,
            in2 => \N__28350\,
            in3 => \N__35379\,
            lcout => n2223,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1382_3_lut_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33393\,
            in2 => \N__31134\,
            in3 => \N__35258\,
            lcout => n2126,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1448_3_lut_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__28311\,
            in1 => \_gnd_net_\,
            in2 => \N__28575\,
            in3 => \N__35378\,
            lcout => n2224,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1372_3_lut_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__33180\,
            in1 => \_gnd_net_\,
            in2 => \N__31239\,
            in3 => \N__35262\,
            lcout => n2116,
            ltout => \n2116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12995_4_lut_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31356\,
            in1 => \N__28272\,
            in2 => \N__28266\,
            in3 => \N__31217\,
            lcout => n2148,
            ltout => \n2148_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1451_3_lut_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28223\,
            in2 => \N__28263\,
            in3 => \N__28260\,
            lcout => n2227,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1384_3_lut_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31152\,
            in2 => \N__35288\,
            in3 => \N__33810\,
            lcout => n2128,
            ltout => \n2128_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28420\,
            in1 => \N__28600\,
            in2 => \N__28584\,
            in3 => \N__31181\,
            lcout => n14316,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1381_3_lut_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__31122\,
            in1 => \_gnd_net_\,
            in2 => \N__35280\,
            in3 => \N__33420\,
            lcout => n2125,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1441_3_lut_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28548\,
            in2 => \N__28896\,
            in3 => \N__35409\,
            lcout => n2217,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1439_3_lut_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__28506\,
            in1 => \N__28500\,
            in2 => \N__35441\,
            in3 => \_gnd_net_\,
            lcout => n2215,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12992_1_lut_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35408\,
            lcout => n15722,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1440_3_lut_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__28461\,
            in1 => \_gnd_net_\,
            in2 => \N__35442\,
            in3 => \N__31345\,
            lcout => n2216,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1378_3_lut_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31101\,
            in2 => \N__33270\,
            in3 => \N__35244\,
            lcout => n2122,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1380_3_lut_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31113\,
            in2 => \N__35281\,
            in3 => \N__33465\,
            lcout => n2124,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1593_3_lut_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__28407\,
            in1 => \_gnd_net_\,
            in2 => \N__35738\,
            in3 => \N__38344\,
            lcout => n2433,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1582_3_lut_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28932\,
            in2 => \N__28923\,
            in3 => \N__35702\,
            lcout => n2422,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1374_3_lut_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31254\,
            in2 => \N__41272\,
            in3 => \N__35279\,
            lcout => n2118,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1585_3_lut_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28872\,
            in2 => \N__28859\,
            in3 => \N__35695\,
            lcout => n2425,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1589_3_lut_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__28833\,
            in1 => \_gnd_net_\,
            in2 => \N__35739\,
            in3 => \N__28803\,
            lcout => n2429,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1581_3_lut_LC_5_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28790\,
            in2 => \N__28761\,
            in3 => \N__35703\,
            lcout => n2421,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1591_3_lut_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28749\,
            in2 => \N__35743\,
            in3 => \N__28736\,
            lcout => n2431,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1580_3_lut_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28704\,
            in2 => \N__28692\,
            in3 => \N__35723\,
            lcout => n2420,
            ltout => \n2420_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_81_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31753\,
            in1 => \N__34030\,
            in2 => \N__28659\,
            in3 => \N__28656\,
            lcout => n14628,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1590_3_lut_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28650\,
            in2 => \N__28638\,
            in3 => \N__35722\,
            lcout => n2430,
            ltout => \n2430_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_82_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__31531\,
            in1 => \N__31606\,
            in2 => \N__29139\,
            in3 => \N__29085\,
            lcout => n13828,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1592_3_lut_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29136\,
            in2 => \N__29124\,
            in3 => \N__35718\,
            lcout => n2432,
            ltout => \n2432_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9990_3_lut_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__33605\,
            in1 => \_gnd_net_\,
            in2 => \N__29088\,
            in3 => \N__31909\,
            lcout => n11967,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1656_3_lut_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31515\,
            in2 => \N__31542\,
            in3 => \N__35867\,
            lcout => n2528,
            ltout => \n2528_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1723_3_lut_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__32178\,
            in1 => \_gnd_net_\,
            in2 => \N__29079\,
            in3 => \N__36057\,
            lcout => n2627,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1576_3_lut_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29040\,
            in2 => \N__29028\,
            in3 => \N__35746\,
            lcout => n2416,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_149_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32695\,
            in1 => \N__28992\,
            in2 => \N__33871\,
            in3 => \N__28986\,
            lcout => n14634,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1577_3_lut_LC_5_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28980\,
            in2 => \N__28947\,
            in3 => \N__35747\,
            lcout => n2417,
            ltout => \n2417_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1644_3_lut_LC_5_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__35868\,
            in1 => \_gnd_net_\,
            in2 => \N__29163\,
            in3 => \N__31680\,
            lcout => n2516,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1659_3_lut_LC_5_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31623\,
            in2 => \N__31641\,
            in3 => \N__35866\,
            lcout => n2531,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_160_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__29145\,
            in1 => \N__32330\,
            in2 => \N__29268\,
            in3 => \N__34134\,
            lcout => n14188,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1642_3_lut_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__32053\,
            in1 => \N__32031\,
            in2 => \N__35897\,
            in3 => \_gnd_net_\,
            lcout => n2514,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1648_3_lut_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31737\,
            in2 => \N__31764\,
            in3 => \N__35855\,
            lcout => n2520,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_150_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31666\,
            in1 => \N__31691\,
            in2 => \N__32055\,
            in3 => \N__29160\,
            lcout => OPEN,
            ltout => \n14640_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13075_4_lut_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31972\,
            in1 => \N__32008\,
            in2 => \N__29154\,
            in3 => \N__31940\,
            lcout => n2445,
            ltout => \n2445_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1657_3_lut_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__31554\,
            in1 => \_gnd_net_\,
            in2 => \N__29151\,
            in3 => \N__31572\,
            lcout => n2529,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1658_3_lut_LC_5_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31611\,
            in2 => \N__31587\,
            in3 => \N__35856\,
            lcout => n2530,
            ltout => \n2530_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_158_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29148\,
            in3 => \N__32233\,
            lcout => n14646,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1661_3_lut_LC_5_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31278\,
            in1 => \N__33609\,
            in2 => \_gnd_net_\,
            in3 => \N__35870\,
            lcout => n2533,
            ltout => \n2533_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10086_4_lut_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__31834\,
            in1 => \N__35141\,
            in2 => \N__29271\,
            in3 => \N__32305\,
            lcout => n12063,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1728_3_lut_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31865\,
            in2 => \N__31851\,
            in3 => \N__36011\,
            lcout => n2632,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1640_3_lut_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31953\,
            in2 => \N__35899\,
            in3 => \N__31980\,
            lcout => n2512,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1643_3_lut_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31671\,
            in2 => \N__31650\,
            in3 => \N__35874\,
            lcout => n2515,
            ltout => \n2515_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_27_LC_5_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29220\,
            in1 => \N__32818\,
            in2 => \N__29214\,
            in3 => \N__29211\,
            lcout => OPEN,
            ltout => \n14194_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13103_4_lut_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32780\,
            in1 => \N__32579\,
            in2 => \N__29202\,
            in3 => \N__32750\,
            lcout => n2544,
            ltout => \n2544_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1727_3_lut_LC_5_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__31835\,
            in1 => \_gnd_net_\,
            in2 => \N__29199\,
            in3 => \N__31821\,
            lcout => n2631,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1641_3_lut_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31992\,
            in2 => \N__32022\,
            in3 => \N__35896\,
            lcout => n2513,
            ltout => \n2513_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1708_3_lut_LC_5_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__36031\,
            in1 => \_gnd_net_\,
            in2 => \N__29547\,
            in3 => \N__32769\,
            lcout => n2612,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1725_3_lut_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32253\,
            in2 => \N__32274\,
            in3 => \N__36023\,
            lcout => n2629,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13100_1_lut_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36070\,
            in3 => \_gnd_net_\,
            lcout => n15830,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1931_3_lut_LC_5_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29472\,
            in2 => \N__34321\,
            in3 => \N__29453\,
            lcout => n2931,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1726_3_lut_LC_5_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__32283\,
            in1 => \_gnd_net_\,
            in2 => \N__36069\,
            in3 => \N__32306\,
            lcout => n2630,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1716_3_lut_LC_5_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32466\,
            in2 => \N__34014\,
            in3 => \N__36030\,
            lcout => n2620,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1933_3_lut_LC_5_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33500\,
            in1 => \N__29352\,
            in2 => \_gnd_net_\,
            in3 => \N__34282\,
            lcout => n2933,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1923_3_lut_LC_5_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29340\,
            in2 => \N__34315\,
            in3 => \N__29313\,
            lcout => n2923,
            ltout => \n2923_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_68_LC_5_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29848\,
            in1 => \N__29701\,
            in2 => \N__29280\,
            in3 => \N__30172\,
            lcout => n14214,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1928_3_lut_LC_5_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29907\,
            in2 => \N__29895\,
            in3 => \N__34263\,
            lcout => n2928,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1920_3_lut_LC_5_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29832\,
            in2 => \N__34314\,
            in3 => \N__29805\,
            lcout => n2920,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12688_1_lut_LC_5_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34660\,
            lcout => n15418,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1913_3_lut_LC_5_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__34271\,
            in1 => \N__29793\,
            in2 => \N__29781\,
            in3 => \_gnd_net_\,
            lcout => n2913,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1925_3_lut_LC_5_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29751\,
            in2 => \N__29739\,
            in3 => \N__34267\,
            lcout => n2925,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1711_3_lut_LC_5_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32319\,
            in2 => \N__36100\,
            in3 => \N__32349\,
            lcout => n2615,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1930_3_lut_LC_5_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29648\,
            in2 => \N__29616\,
            in3 => \N__34322\,
            lcout => n2930,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1991_3_lut_LC_5_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29574\,
            in2 => \N__34504\,
            in3 => \N__29561\,
            lcout => n3023,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1980_3_lut_LC_5_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30290\,
            in2 => \N__30270\,
            in3 => \N__34472\,
            lcout => n3012,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10076_4_lut_LC_5_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__35177\,
            in1 => \N__30220\,
            in2 => \N__30008\,
            in3 => \N__30140\,
            lcout => n12053,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1987_3_lut_LC_5_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30192\,
            in2 => \N__30180\,
            in3 => \N__34468\,
            lcout => n3019,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1999_3_lut_LC_5_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30156\,
            in2 => \N__30144\,
            in3 => \N__34466\,
            lcout => n3031,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2001_3_lut_LC_5_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__30111\,
            in1 => \N__35176\,
            in2 => \N__34503\,
            in3 => \_gnd_net_\,
            lcout => n3033,
            ltout => \n3033_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9970_3_lut_LC_5_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41563\,
            in2 => \N__30081\,
            in3 => \N__30073\,
            lcout => n11947,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2118_3_lut_LC_5_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30057\,
            in2 => \N__30045\,
            in3 => \N__34889\,
            lcout => n3214,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1998_3_lut_LC_5_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30021\,
            in2 => \N__30009\,
            in3 => \N__34467\,
            lcout => n3030,
            ltout => \n3030_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_167_LC_5_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__29947\,
            in1 => \N__29926\,
            in2 => \N__30633\,
            in3 => \N__30630\,
            lcout => OPEN,
            ltout => \n13871_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_169_LC_5_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30608\,
            in1 => \N__30580\,
            in2 => \N__30564\,
            in3 => \N__30544\,
            lcout => n14078,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2135_3_lut_LC_5_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30519\,
            in2 => \N__34915\,
            in3 => \N__30506\,
            lcout => n3231,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2132_3_lut_LC_5_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30488\,
            in2 => \N__30468\,
            in3 => \N__34890\,
            lcout => n3228,
            ltout => \n3228_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_125_LC_5_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37129\,
            in2 => \N__30453\,
            in3 => \N__30450\,
            lcout => n14770,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2136_3_lut_LC_5_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30444\,
            in2 => \N__30431\,
            in3 => \N__34891\,
            lcout => n3232,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2134_3_lut_LC_5_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30405\,
            in2 => \N__34916\,
            in3 => \N__30389\,
            lcout => n3230,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1984_3_lut_LC_5_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30369\,
            in2 => \N__30339\,
            in3 => \N__34505\,
            lcout => n3016,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_129_LC_5_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37048\,
            in1 => \N__37598\,
            in2 => \N__37211\,
            in3 => \N__32868\,
            lcout => n14025,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2127_3_lut_LC_5_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30816\,
            in2 => \N__30786\,
            in3 => \N__34835\,
            lcout => n3223,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12759_4_lut_LC_5_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__37639\,
            in1 => \N__30774\,
            in2 => \N__30768\,
            in3 => \N__32973\,
            lcout => n3237,
            ltout => \n3237_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2200_3_lut_LC_5_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36774\,
            in2 => \N__30759\,
            in3 => \N__36801\,
            lcout => n13_adj_713,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2115_3_lut_LC_5_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__30750\,
            in1 => \_gnd_net_\,
            in2 => \N__34888\,
            in3 => \N__30730\,
            lcout => n3211,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_126_LC_5_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37399\,
            in1 => \N__37366\,
            in2 => \N__37472\,
            in3 => \N__30711\,
            lcout => OPEN,
            ltout => \n14776_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_127_LC_5_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37273\,
            in1 => \N__37333\,
            in2 => \N__30705\,
            in3 => \N__37247\,
            lcout => n14782,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2125_3_lut_LC_5_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30702\,
            in2 => \N__30681\,
            in3 => \N__34839\,
            lcout => n3221,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2119_3_lut_LC_5_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30669\,
            in2 => \N__30645\,
            in3 => \N__34866\,
            lcout => n3215,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2121_3_lut_LC_5_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__30903\,
            in1 => \_gnd_net_\,
            in2 => \N__34908\,
            in3 => \N__30894\,
            lcout => n3217,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2193_3_lut_LC_5_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37094\,
            in2 => \N__35088\,
            in3 => \N__37074\,
            lcout => OPEN,
            ltout => \n27_adj_716_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_87_LC_5_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__37471\,
            in1 => \N__37449\,
            in2 => \N__30870\,
            in3 => \N__35050\,
            lcout => n14266,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_91_LC_5_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001010"
        )
    port map (
            in0 => \N__36738\,
            in1 => \N__36758\,
            in2 => \N__35090\,
            in3 => \N__30861\,
            lcout => n14268,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2189_3_lut_LC_5_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36932\,
            in2 => \N__36918\,
            in3 => \N__35049\,
            lcout => n35_adj_719,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2198_3_lut_LC_5_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36696\,
            in2 => \N__35089\,
            in3 => \N__36716\,
            lcout => OPEN,
            ltout => \n17_adj_714_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_93_LC_5_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__37416\,
            in1 => \N__37436\,
            in2 => \N__30855\,
            in3 => \N__35057\,
            lcout => n14272,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2112_3_lut_LC_5_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30851\,
            in2 => \N__30831\,
            in3 => \N__34874\,
            lcout => n3208,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2190_3_lut_LC_5_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36986\,
            in2 => \N__36954\,
            in3 => \N__35091\,
            lcout => OPEN,
            ltout => \n33_adj_718_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_94_LC_5_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__35092\,
            in1 => \N__37113\,
            in2 => \N__30819\,
            in3 => \N__37139\,
            lcout => OPEN,
            ltout => \n14262_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_97_LC_5_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31089\,
            in1 => \N__31083\,
            in2 => \N__31077\,
            in3 => \N__31074\,
            lcout => n14284,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2114_3_lut_LC_5_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31068\,
            in2 => \N__31047\,
            in3 => \N__34870\,
            lcout => n3210,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2113_3_lut_LC_5_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31032\,
            in2 => \N__34909\,
            in3 => \N__31011\,
            lcout => n3209,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1507_3_lut_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31002\,
            in2 => \N__30993\,
            in3 => \N__35597\,
            lcout => n2315,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_2_lut_LC_6_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38087\,
            in2 => \_gnd_net_\,
            in3 => \N__30930\,
            lcout => n2101,
            ltout => OPEN,
            carryin => \bfn_6_17_0_\,
            carryout => n12639,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_3_lut_LC_6_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55346\,
            in2 => \N__33732\,
            in3 => \N__30927\,
            lcout => n2100,
            ltout => OPEN,
            carryin => n12639,
            carryout => n12640,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_4_lut_LC_6_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33368\,
            in3 => \N__30915\,
            lcout => n2099,
            ltout => OPEN,
            carryin => n12640,
            carryout => n12641,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_5_lut_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55347\,
            in2 => \N__33341\,
            in3 => \N__30906\,
            lcout => n2098,
            ltout => OPEN,
            carryin => n12641,
            carryout => n12642,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_6_lut_LC_6_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33776\,
            in3 => \N__31155\,
            lcout => n2097,
            ltout => OPEN,
            carryin => n12642,
            carryout => n12643,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_7_lut_LC_6_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33806\,
            in3 => \N__31146\,
            lcout => n2096,
            ltout => OPEN,
            carryin => n12643,
            carryout => n12644,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_8_lut_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55045\,
            in2 => \N__33443\,
            in3 => \N__31137\,
            lcout => n2095,
            ltout => OPEN,
            carryin => n12644,
            carryout => n12645,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_9_lut_LC_6_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55348\,
            in2 => \N__33392\,
            in3 => \N__31125\,
            lcout => n2094,
            ltout => OPEN,
            carryin => n12645,
            carryout => n12646,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_10_lut_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55157\,
            in2 => \N__33419\,
            in3 => \N__31116\,
            lcout => n2093,
            ltout => OPEN,
            carryin => \bfn_6_18_0_\,
            carryout => n12647,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_11_lut_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55160\,
            in2 => \N__33464\,
            in3 => \N__31107\,
            lcout => n2092,
            ltout => OPEN,
            carryin => n12647,
            carryout => n12648,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_12_lut_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33287\,
            in2 => \N__55345\,
            in3 => \N__31104\,
            lcout => n2091,
            ltout => OPEN,
            carryin => n12648,
            carryout => n12649,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_13_lut_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55164\,
            in2 => \N__33269\,
            in3 => \N__31095\,
            lcout => n2090,
            ltout => OPEN,
            carryin => n12649,
            carryout => n12650,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_14_lut_LC_6_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55158\,
            in2 => \N__33314\,
            in3 => \N__31092\,
            lcout => n2089,
            ltout => OPEN,
            carryin => n12650,
            carryout => n12651,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_15_lut_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55165\,
            in2 => \N__33141\,
            in3 => \N__31260\,
            lcout => n2088,
            ltout => OPEN,
            carryin => n12651,
            carryout => n12652,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_16_lut_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55159\,
            in2 => \N__33084\,
            in3 => \N__31257\,
            lcout => n2087,
            ltout => OPEN,
            carryin => n12652,
            carryout => n12653,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_17_lut_LC_6_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55166\,
            in2 => \N__41274\,
            in3 => \N__31245\,
            lcout => n2086,
            ltout => OPEN,
            carryin => n12653,
            carryout => n12654,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_18_lut_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31377\,
            in2 => \N__55490\,
            in3 => \N__31242\,
            lcout => n2085,
            ltout => OPEN,
            carryin => \bfn_6_19_0_\,
            carryout => n12655,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_19_lut_LC_6_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33176\,
            in2 => \N__55240\,
            in3 => \N__31230\,
            lcout => n2084,
            ltout => OPEN,
            carryin => n12655,
            carryout => n12656,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1369_20_lut_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__55344\,
            in1 => \N__35315\,
            in2 => \N__37929\,
            in3 => \N__31227\,
            lcout => n2115,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1379_3_lut_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31206\,
            in2 => \N__33291\,
            in3 => \N__35257\,
            lcout => n2123,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_148_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33140\,
            in1 => \N__33083\,
            in2 => \N__41273\,
            in3 => \N__33750\,
            lcout => OPEN,
            ltout => \n14558_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12970_4_lut_LC_6_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31376\,
            in1 => \N__33175\,
            in2 => \N__31392\,
            in3 => \N__37925\,
            lcout => n2049,
            ltout => \n2049_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1389_3_lut_LC_6_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__31389\,
            in1 => \_gnd_net_\,
            in2 => \N__31380\,
            in3 => \N__38088\,
            lcout => n2133,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1311_3_lut_LC_6_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38064\,
            in2 => \N__41132\,
            in3 => \N__41359\,
            lcout => n2023,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12967_1_lut_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35277\,
            lcout => n15697,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1306_3_lut_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38142\,
            in2 => \N__37986\,
            in3 => \N__41374\,
            lcout => n2018,
            ltout => \n2018_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1373_3_lut_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__35278\,
            in1 => \N__31365\,
            in2 => \N__31359\,
            in3 => \_gnd_net_\,
            lcout => n2117,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1377_3_lut_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31323\,
            in2 => \N__33315\,
            in3 => \N__35276\,
            lcout => n2121,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_2_lut_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33601\,
            in2 => \_gnd_net_\,
            in3 => \N__31266\,
            lcout => n2501,
            ltout => OPEN,
            carryin => \bfn_6_21_0_\,
            carryout => n12717,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_3_lut_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54787\,
            in2 => \N__31916\,
            in3 => \N__31263\,
            lcout => n2500,
            ltout => OPEN,
            carryin => n12717,
            carryout => n12718,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_4_lut_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31640\,
            in3 => \N__31614\,
            lcout => n2499,
            ltout => OPEN,
            carryin => n12718,
            carryout => n12719,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_5_lut_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54788\,
            in2 => \N__31610\,
            in3 => \N__31575\,
            lcout => n2498,
            ltout => OPEN,
            carryin => n12719,
            carryout => n12720,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_6_lut_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31571\,
            in3 => \N__31545\,
            lcout => n2497,
            ltout => OPEN,
            carryin => n12720,
            carryout => n12721,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_7_lut_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31538\,
            in3 => \N__31509\,
            lcout => n2496,
            ltout => OPEN,
            carryin => n12721,
            carryout => n12722,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_8_lut_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54763\,
            in2 => \N__31506\,
            in3 => \N__31467\,
            lcout => n2495,
            ltout => OPEN,
            carryin => n12722,
            carryout => n12723,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_9_lut_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31463\,
            in2 => \N__55041\,
            in3 => \N__31437\,
            lcout => n2494,
            ltout => OPEN,
            carryin => n12723,
            carryout => n12724,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_10_lut_LC_6_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54756\,
            in2 => \N__33984\,
            in3 => \N__31434\,
            lcout => n2493,
            ltout => OPEN,
            carryin => \bfn_6_22_0_\,
            carryout => n12725,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_11_lut_LC_6_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54784\,
            in2 => \N__31431\,
            in3 => \N__31395\,
            lcout => n2492,
            ltout => OPEN,
            carryin => n12725,
            carryout => n12726,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_12_lut_LC_6_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54757\,
            in2 => \N__31812\,
            in3 => \N__31773\,
            lcout => n2491,
            ltout => OPEN,
            carryin => n12726,
            carryout => n12727,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_13_lut_LC_6_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54785\,
            in2 => \N__34119\,
            in3 => \N__31770\,
            lcout => n2490,
            ltout => OPEN,
            carryin => n12727,
            carryout => n12728,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_14_lut_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54758\,
            in2 => \N__34043\,
            in3 => \N__31767\,
            lcout => n2489,
            ltout => OPEN,
            carryin => n12728,
            carryout => n12729,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_15_lut_LC_6_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31760\,
            in2 => \N__55040\,
            in3 => \N__31731\,
            lcout => n2488,
            ltout => OPEN,
            carryin => n12729,
            carryout => n12730,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_16_lut_LC_6_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54762\,
            in2 => \N__31727\,
            in3 => \N__31701\,
            lcout => n2487,
            ltout => OPEN,
            carryin => n12730,
            carryout => n12731,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_17_lut_LC_6_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54786\,
            in2 => \N__33878\,
            in3 => \N__31698\,
            lcout => n2486,
            ltout => OPEN,
            carryin => n12731,
            carryout => n12732,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_18_lut_LC_6_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54746\,
            in2 => \N__32702\,
            in3 => \N__31695\,
            lcout => n2485,
            ltout => OPEN,
            carryin => \bfn_6_23_0_\,
            carryout => n12733,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_19_lut_LC_6_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31692\,
            in2 => \N__55037\,
            in3 => \N__31674\,
            lcout => n2484,
            ltout => OPEN,
            carryin => n12733,
            carryout => n12734,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_20_lut_LC_6_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31667\,
            in2 => \N__55055\,
            in3 => \N__32058\,
            lcout => n2483,
            ltout => OPEN,
            carryin => n12734,
            carryout => n12735,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_21_lut_LC_6_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32054\,
            in2 => \N__55038\,
            in3 => \N__32025\,
            lcout => n2482,
            ltout => OPEN,
            carryin => n12735,
            carryout => n12736,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_22_lut_LC_6_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32015\,
            in2 => \N__55056\,
            in3 => \N__31983\,
            lcout => n2481,
            ltout => OPEN,
            carryin => n12736,
            carryout => n12737,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_23_lut_LC_6_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31979\,
            in2 => \N__55039\,
            in3 => \N__31947\,
            lcout => n2480,
            ltout => OPEN,
            carryin => n12737,
            carryout => n12738,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1637_24_lut_LC_6_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__54783\,
            in1 => \N__31944\,
            in2 => \N__35948\,
            in3 => \N__31923\,
            lcout => n2511,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1660_3_lut_LC_6_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31920\,
            in2 => \N__31893\,
            in3 => \N__35869\,
            lcout => n2532,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_2_lut_LC_6_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35137\,
            in2 => \_gnd_net_\,
            in3 => \N__31869\,
            lcout => n2601,
            ltout => OPEN,
            carryin => \bfn_6_24_0_\,
            carryout => n12739,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_3_lut_LC_6_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53816\,
            in2 => \N__31866\,
            in3 => \N__31842\,
            lcout => n2600,
            ltout => OPEN,
            carryin => n12739,
            carryout => n12740,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_4_lut_LC_6_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31839\,
            in3 => \N__31815\,
            lcout => n2599,
            ltout => OPEN,
            carryin => n12740,
            carryout => n12741,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_5_lut_LC_6_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53817\,
            in2 => \N__32310\,
            in3 => \N__32277\,
            lcout => n2598,
            ltout => OPEN,
            carryin => n12741,
            carryout => n12742,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_6_lut_LC_6_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32270\,
            in3 => \N__32247\,
            lcout => n2597,
            ltout => OPEN,
            carryin => n12742,
            carryout => n12743,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_7_lut_LC_6_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32240\,
            in3 => \N__32202\,
            lcout => n2596,
            ltout => OPEN,
            carryin => n12743,
            carryout => n12744,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_8_lut_LC_6_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53819\,
            in2 => \N__32199\,
            in3 => \N__32169\,
            lcout => n2595,
            ltout => OPEN,
            carryin => n12744,
            carryout => n12745,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_9_lut_LC_6_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53818\,
            in2 => \N__32166\,
            in3 => \N__32133\,
            lcout => n2594,
            ltout => OPEN,
            carryin => n12745,
            carryout => n12746,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_10_lut_LC_6_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54506\,
            in2 => \N__32130\,
            in3 => \N__32097\,
            lcout => n2593,
            ltout => OPEN,
            carryin => \bfn_6_25_0_\,
            carryout => n12747,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_11_lut_LC_6_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54417\,
            in2 => \N__33951\,
            in3 => \N__32094\,
            lcout => n2592,
            ltout => OPEN,
            carryin => n12747,
            carryout => n12748,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_12_lut_LC_6_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32091\,
            in2 => \N__54776\,
            in3 => \N__32523\,
            lcout => n2591,
            ltout => OPEN,
            carryin => n12748,
            carryout => n12749,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_13_lut_LC_6_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54421\,
            in2 => \N__32520\,
            in3 => \N__32487\,
            lcout => n2590,
            ltout => OPEN,
            carryin => n12749,
            carryout => n12750,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_14_lut_LC_6_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54507\,
            in2 => \N__34082\,
            in3 => \N__32469\,
            lcout => n2589,
            ltout => OPEN,
            carryin => n12750,
            carryout => n12751,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_15_lut_LC_6_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54422\,
            in2 => \N__34010\,
            in3 => \N__32457\,
            lcout => n2588,
            ltout => OPEN,
            carryin => n12751,
            carryout => n12752,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_16_lut_LC_6_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54508\,
            in2 => \N__32454\,
            in3 => \N__32418\,
            lcout => n2587,
            ltout => OPEN,
            carryin => n12752,
            carryout => n12753,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_17_lut_LC_6_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54423\,
            in2 => \N__32415\,
            in3 => \N__32373\,
            lcout => n2586,
            ltout => OPEN,
            carryin => n12753,
            carryout => n12754,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_18_lut_LC_6_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33839\,
            in2 => \N__54744\,
            in3 => \N__32355\,
            lcout => n2585,
            ltout => OPEN,
            carryin => \bfn_6_26_0_\,
            carryout => n12755,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_19_lut_LC_6_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54373\,
            in2 => \N__32657\,
            in3 => \N__32352\,
            lcout => n2584,
            ltout => OPEN,
            carryin => n12755,
            carryout => n12756,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_20_lut_LC_6_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54379\,
            in2 => \N__32348\,
            in3 => \N__32313\,
            lcout => n2583,
            ltout => OPEN,
            carryin => n12756,
            carryout => n12757,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_21_lut_LC_6_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54374\,
            in2 => \N__32862\,
            in3 => \N__32832\,
            lcout => n2582,
            ltout => OPEN,
            carryin => n12757,
            carryout => n12758,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_22_lut_LC_6_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54380\,
            in2 => \N__32829\,
            in3 => \N__32787\,
            lcout => n2581,
            ltout => OPEN,
            carryin => n12758,
            carryout => n12759,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_23_lut_LC_6_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54375\,
            in2 => \N__32784\,
            in3 => \N__32763\,
            lcout => n2580,
            ltout => OPEN,
            carryin => n12759,
            carryout => n12760,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_24_lut_LC_6_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32591\,
            in2 => \N__54745\,
            in3 => \N__32760\,
            lcout => n2579,
            ltout => OPEN,
            carryin => n12760,
            carryout => n12761,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1704_25_lut_LC_6_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__54381\,
            in1 => \N__36113\,
            in2 => \N__32757\,
            in3 => \N__32739\,
            lcout => n2610,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1645_3_lut_LC_6_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32703\,
            in2 => \N__32673\,
            in3 => \N__35900\,
            lcout => n2517,
            ltout => \n2517_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1712_3_lut_LC_6_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32637\,
            in2 => \N__32631\,
            in3 => \N__36098\,
            lcout => n2616,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1707_3_lut_LC_6_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__32592\,
            in1 => \_gnd_net_\,
            in2 => \N__32568\,
            in3 => \N__36099\,
            lcout => n2611,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12755_1_lut_LC_6_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35099\,
            lcout => n15485,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2133_3_lut_LC_6_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32961\,
            in2 => \N__32943\,
            in3 => \N__34917\,
            lcout => n3229,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2129_3_lut_LC_6_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32928\,
            in2 => \N__34923\,
            in3 => \N__32915\,
            lcout => n3225,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12562_1_lut_LC_6_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36297\,
            lcout => n15292,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i8_1_lut_LC_6_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36135\,
            lcout => n18_adj_558,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2137_3_lut_LC_6_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32889\,
            in1 => \N__34165\,
            in2 => \_gnd_net_\,
            in3 => \N__34918\,
            lcout => n3233,
            ltout => \n3233_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9966_3_lut_LC_6_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__36592\,
            in1 => \_gnd_net_\,
            in2 => \N__32874\,
            in3 => \N__36895\,
            lcout => OPEN,
            ltout => \n11943_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_120_LC_6_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__36793\,
            in1 => \N__36832\,
            in2 => \N__32871\,
            in3 => \N__36865\,
            lcout => n13875,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2192_3_lut_LC_6_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37032\,
            in2 => \N__37058\,
            in3 => \N__35035\,
            lcout => OPEN,
            ltout => \n29_adj_717_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_88_LC_6_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__35036\,
            in1 => \N__37207\,
            in2 => \N__33003\,
            in3 => \N__37185\,
            lcout => n14270,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9964_4_lut_LC_6_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__32985\,
            in1 => \N__36540\,
            in2 => \N__36558\,
            in3 => \N__35038\,
            lcout => OPEN,
            ltout => \n11941_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10062_4_lut_LC_6_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__35039\,
            in1 => \N__36879\,
            in2 => \N__32988\,
            in3 => \N__36899\,
            lcout => n12039,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9902_4_lut_LC_6_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111100"
        )
    port map (
            in0 => \N__36594\,
            in1 => \N__36618\,
            in2 => \N__36570\,
            in3 => \N__35037\,
            lcout => n11878,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12763_4_lut_LC_6_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100111"
        )
    port map (
            in0 => \N__35040\,
            in1 => \N__37554\,
            in2 => \N__37521\,
            in3 => \N__33060\,
            lcout => n12051,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_130_LC_6_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37753\,
            in1 => \N__37672\,
            in2 => \N__37716\,
            in3 => \N__32979\,
            lcout => n14788,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_113_LC_6_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111000"
        )
    port map (
            in0 => \N__37754\,
            in1 => \N__35076\,
            in2 => \N__37731\,
            in3 => \N__33009\,
            lcout => OPEN,
            ltout => \n14300_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_114_LC_6_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__35077\,
            in1 => \N__37714\,
            in2 => \N__32967\,
            in3 => \N__37689\,
            lcout => OPEN,
            ltout => \n14302_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_115_LC_6_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__37673\,
            in1 => \N__37653\,
            in2 => \N__32964\,
            in3 => \N__35078\,
            lcout => OPEN,
            ltout => \n14304_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_116_LC_6_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__35079\,
            in1 => \N__37611\,
            in2 => \N__33066\,
            in3 => \N__37641\,
            lcout => OPEN,
            ltout => \n14306_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_117_LC_6_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__37599\,
            in1 => \N__37566\,
            in2 => \N__33063\,
            in3 => \N__35080\,
            lcout => n14308,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16_4_lut_LC_6_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__36813\,
            in1 => \N__36866\,
            in2 => \N__35095\,
            in3 => \N__36833\,
            lcout => n5_adj_704,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_103_LC_6_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__33162\,
            in1 => \N__33054\,
            in2 => \N__33048\,
            in3 => \N__33024\,
            lcout => OPEN,
            ltout => \n14292_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_104_LC_6_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__37307\,
            in1 => \N__37290\,
            in2 => \N__33036\,
            in3 => \N__35068\,
            lcout => n14294,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_98_LC_6_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001010"
        )
    port map (
            in0 => \N__37383\,
            in1 => \N__37403\,
            in2 => \N__35093\,
            in3 => \N__33033\,
            lcout => OPEN,
            ltout => \n14286_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_102_LC_6_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__37374\,
            in1 => \N__37350\,
            in2 => \N__33027\,
            in3 => \N__35067\,
            lcout => n14288,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_109_LC_6_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001010"
        )
    port map (
            in0 => \N__37257\,
            in1 => \N__37277\,
            in2 => \N__35094\,
            in3 => \N__33018\,
            lcout => OPEN,
            ltout => \n14296_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_111_LC_6_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__37224\,
            in1 => \N__37246\,
            in2 => \N__33012\,
            in3 => \N__35072\,
            lcout => n14298,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i2184_3_lut_LC_6_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37341\,
            in2 => \N__37320\,
            in3 => \N__35066\,
            lcout => n45_adj_720,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.a_new_i0_LC_6_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33156\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \quad_counter0.a_new_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1318_3_lut_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37866\,
            in2 => \N__39354\,
            in3 => \N__41370\,
            lcout => n2030,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1242_3_lut_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__41007\,
            in1 => \_gnd_net_\,
            in2 => \N__43035\,
            in3 => \N__41515\,
            lcout => n1922,
            ltout => \n1922_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1309_3_lut_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38016\,
            in2 => \N__33144\,
            in3 => \N__41357\,
            lcout => n2021,
            ltout => \n2021_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1376_3_lut_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__33123\,
            in1 => \_gnd_net_\,
            in2 => \N__33117\,
            in3 => \N__35296\,
            lcout => n2120,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1317_3_lut_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39123\,
            in2 => \N__37854\,
            in3 => \N__41356\,
            lcout => n2029,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10008_4_lut_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001000"
        )
    port map (
            in0 => \N__38118\,
            in1 => \N__39536\,
            in2 => \N__39321\,
            in3 => \N__39353\,
            lcout => n11985,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1308_3_lut_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37911\,
            in2 => \N__38004\,
            in3 => \N__41358\,
            lcout => n2020,
            ltout => \n2020_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1375_3_lut_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33237\,
            in2 => \N__33231\,
            in3 => \N__35297\,
            lcout => n2119,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1316_3_lut_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39285\,
            in2 => \N__37836\,
            in3 => \N__41332\,
            lcout => n2028,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12944_1_lut_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41367\,
            in3 => \_gnd_net_\,
            lcout => n15674,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1315_3_lut_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39246\,
            in2 => \N__37818\,
            in3 => \N__41333\,
            lcout => n2027,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_142_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38027\,
            in1 => \N__37906\,
            in2 => \N__39555\,
            in3 => \N__41103\,
            lcout => OPEN,
            ltout => \n14446_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_144_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__38169\,
            in1 => \N__41420\,
            in2 => \N__33195\,
            in3 => \N__33192\,
            lcout => OPEN,
            ltout => \n14450_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12947_4_lut_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__38138\,
            in1 => \N__41636\,
            in2 => \N__33186\,
            in3 => \N__38159\,
            lcout => n1950,
            ltout => \n1950_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1305_3_lut_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__38160\,
            in1 => \_gnd_net_\,
            in2 => \N__33183\,
            in3 => \N__37968\,
            lcout => n2017,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1319_3_lut_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__37881\,
            in1 => \_gnd_net_\,
            in2 => \N__41366\,
            in3 => \N__39540\,
            lcout => n2031,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1314_3_lut_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37800\,
            in2 => \N__41745\,
            in3 => \N__41340\,
            lcout => n2026,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1312_3_lut_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39612\,
            in2 => \N__41368\,
            in3 => \N__37770\,
            lcout => n2024,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1313_3_lut_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37785\,
            in2 => \N__41703\,
            in3 => \N__41342\,
            lcout => n2025,
            ltout => \n2025_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_145_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33436\,
            in1 => \N__33412\,
            in2 => \N__33396\,
            in3 => \N__33385\,
            lcout => n14544,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1321_3_lut_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38117\,
            in1 => \N__37506\,
            in2 => \_gnd_net_\,
            in3 => \N__41341\,
            lcout => n2033,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1310_3_lut_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39582\,
            in2 => \N__41369\,
            in3 => \N__38049\,
            lcout => n2022,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1320_3_lut_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39320\,
            in2 => \N__37491\,
            in3 => \N__41343\,
            lcout => n2032,
            ltout => \n2032_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10004_4_lut_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__38080\,
            in1 => \N__33334\,
            in2 => \N__33318\,
            in3 => \N__33721\,
            lcout => n11981,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12922_1_lut_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41519\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n15652,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_146_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33307\,
            in1 => \N__33286\,
            in2 => \N__33268\,
            in3 => \N__33243\,
            lcout => OPEN,
            ltout => \n14550_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_147_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__33816\,
            in1 => \N__33805\,
            in2 => \N__33780\,
            in3 => \N__33775\,
            lcout => n14552,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1388_3_lut_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33744\,
            in2 => \N__33731\,
            in3 => \N__35243\,
            lcout => n2132,
            ltout => \n2132_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9933_3_lut_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33620\,
            in2 => \N__33681\,
            in3 => \N__33661\,
            lcout => n11909,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i13_3_lut_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38364\,
            in1 => \N__49591\,
            in2 => \_gnd_net_\,
            in3 => \N__39972\,
            lcout => n307,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i10_3_lut_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38415\,
            in1 => \N__49592\,
            in2 => \_gnd_net_\,
            in3 => \N__39699\,
            lcout => n310,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i8_3_lut_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49593\,
            in1 => \N__38469\,
            in2 => \_gnd_net_\,
            in3 => \N__39765\,
            lcout => n312,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i7_3_lut_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38490\,
            in1 => \N__49623\,
            in2 => \_gnd_net_\,
            in3 => \N__39384\,
            lcout => n313,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i6_3_lut_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49624\,
            in1 => \N__38511\,
            in2 => \_gnd_net_\,
            in3 => \N__39414\,
            lcout => n314,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i3_3_lut_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38262\,
            in1 => \N__49625\,
            in2 => \_gnd_net_\,
            in3 => \N__39477\,
            lcout => n317,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i2_3_lut_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49626\,
            in1 => \N__38286\,
            in2 => \_gnd_net_\,
            in3 => \N__45804\,
            lcout => n318,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_157_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33944\,
            in1 => \N__33997\,
            in2 => \N__34075\,
            in3 => \N__33832\,
            lcout => n14184,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i1_3_lut_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49621\,
            in1 => \N__38301\,
            in2 => \_gnd_net_\,
            in3 => \N__39513\,
            lcout => n319,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1650_3_lut_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35903\,
            in1 => \N__34125\,
            in2 => \_gnd_net_\,
            in3 => \N__34118\,
            lcout => n2522,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1649_3_lut_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34053\,
            in2 => \N__34047\,
            in3 => \N__35902\,
            lcout => n2521,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12486_3_lut_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33983\,
            in2 => \N__35912\,
            in3 => \N__33957\,
            lcout => n2525,
            ltout => \n2525_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1720_3_lut_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33933\,
            in2 => \N__33924\,
            in3 => \N__36096\,
            lcout => n2624,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1646_3_lut_LC_7_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__35904\,
            in1 => \N__33885\,
            in2 => \N__33879\,
            in3 => \_gnd_net_\,
            lcout => n2518,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i5_3_lut_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49605\,
            in1 => \N__38226\,
            in2 => \_gnd_net_\,
            in3 => \N__39447\,
            lcout => n315,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i9_3_lut_LC_7_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38442\,
            in1 => \N__49604\,
            in2 => \_gnd_net_\,
            in3 => \N__39735\,
            lcout => n311,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i0_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__36627\,
            in1 => \N__40111\,
            in2 => \N__36648\,
            in3 => \N__35118\,
            lcout => encoder0_position_scaled_0,
            ltout => OPEN,
            carryin => \bfn_7_25_0_\,
            carryout => n12952,
            clk => \N__56209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i1_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__35115\,
            in1 => \N__35103\,
            in2 => \N__40169\,
            in3 => \N__34950\,
            lcout => encoder0_position_scaled_1,
            ltout => OPEN,
            carryin => n12952,
            carryout => n12953,
            clk => \N__56209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i2_LC_7_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__34947\,
            in1 => \N__34922\,
            in2 => \N__40173\,
            in3 => \N__34743\,
            lcout => encoder0_position_scaled_2,
            ltout => OPEN,
            carryin => n12953,
            carryout => n12954,
            clk => \N__56209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i3_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__34740\,
            in1 => \N__34715\,
            in2 => \N__40170\,
            in3 => \N__34542\,
            lcout => encoder0_position_scaled_3,
            ltout => OPEN,
            carryin => n12954,
            carryout => n12955,
            clk => \N__56209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i4_LC_7_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__34539\,
            in1 => \N__34515\,
            in2 => \N__40174\,
            in3 => \N__34359\,
            lcout => encoder0_position_scaled_4,
            ltout => OPEN,
            carryin => n12955,
            carryout => n12956,
            clk => \N__56209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i5_LC_7_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__34356\,
            in1 => \N__34334\,
            in2 => \N__40171\,
            in3 => \N__34173\,
            lcout => encoder0_position_scaled_5,
            ltout => OPEN,
            carryin => n12956,
            carryout => n12957,
            clk => \N__56209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i6_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__36492\,
            in1 => \N__36465\,
            in2 => \N__40175\,
            in3 => \N__36312\,
            lcout => encoder0_position_scaled_6,
            ltout => OPEN,
            carryin => n12957,
            carryout => n12958,
            clk => \N__56209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i7_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__36309\,
            in1 => \N__36296\,
            in2 => \N__40172\,
            in3 => \N__36123\,
            lcout => encoder0_position_scaled_7,
            ltout => OPEN,
            carryin => n12958,
            carryout => n12959,
            clk => \N__56209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i8_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__36120\,
            in1 => \N__36101\,
            in2 => \N__40220\,
            in3 => \N__35952\,
            lcout => encoder0_position_scaled_8,
            ltout => OPEN,
            carryin => \bfn_7_26_0_\,
            carryout => n12960,
            clk => \N__56211\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i9_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__35949\,
            in1 => \N__35901\,
            in2 => \N__40224\,
            in3 => \N__35781\,
            lcout => encoder0_position_scaled_9,
            ltout => OPEN,
            carryin => n12960,
            carryout => n12961,
            clk => \N__56211\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i10_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__35778\,
            in1 => \N__35754\,
            in2 => \N__40221\,
            in3 => \N__35628\,
            lcout => encoder0_position_scaled_10,
            ltout => OPEN,
            carryin => n12961,
            carryout => n12962,
            clk => \N__56211\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i11_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__35625\,
            in1 => \N__35601\,
            in2 => \N__40225\,
            in3 => \N__35475\,
            lcout => encoder0_position_scaled_11,
            ltout => OPEN,
            carryin => n12962,
            carryout => n12963,
            clk => \N__56211\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i12_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__35472\,
            in1 => \N__35451\,
            in2 => \N__40222\,
            in3 => \N__35328\,
            lcout => encoder0_position_scaled_12,
            ltout => OPEN,
            carryin => n12963,
            carryout => n12964,
            clk => \N__56211\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i13_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__35325\,
            in1 => \N__35304\,
            in2 => \N__40226\,
            in3 => \N__35181\,
            lcout => encoder0_position_scaled_13,
            ltout => OPEN,
            carryin => n12964,
            carryout => n12965,
            clk => \N__56211\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i14_LC_7_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__37952\,
            in1 => \N__41382\,
            in2 => \N__40223\,
            in3 => \N__36531\,
            lcout => encoder0_position_scaled_14,
            ltout => OPEN,
            carryin => n12965,
            carryout => n12966,
            clk => \N__56211\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i15_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__36528\,
            in1 => \N__41523\,
            in2 => \N__40227\,
            in3 => \N__36516\,
            lcout => encoder0_position_scaled_15,
            ltout => OPEN,
            carryin => n12966,
            carryout => n12967,
            clk => \N__56211\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i16_LC_7_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__45399\,
            in1 => \N__45510\,
            in2 => \N__40228\,
            in3 => \N__36513\,
            lcout => encoder0_position_scaled_16,
            ltout => OPEN,
            carryin => \bfn_7_27_0_\,
            carryout => n12968,
            clk => \N__56214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i17_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__45180\,
            in1 => \N__45621\,
            in2 => \N__40232\,
            in3 => \N__36510\,
            lcout => encoder0_position_scaled_17,
            ltout => OPEN,
            carryin => n12968,
            carryout => n12969,
            clk => \N__56214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i18_LC_7_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__52479\,
            in1 => \N__48900\,
            in2 => \N__40229\,
            in3 => \N__36507\,
            lcout => encoder0_position_scaled_18,
            ltout => OPEN,
            carryin => n12969,
            carryout => n12970,
            clk => \N__56214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i19_LC_7_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__51753\,
            in1 => \N__40206\,
            in2 => \N__49014\,
            in3 => \N__36504\,
            lcout => encoder0_position_scaled_19,
            ltout => OPEN,
            carryin => n12970,
            carryout => n12971,
            clk => \N__56214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i20_LC_7_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__47502\,
            in1 => \N__52359\,
            in2 => \N__40230\,
            in3 => \N__36501\,
            lcout => encoder0_position_scaled_20,
            ltout => OPEN,
            carryin => n12971,
            carryout => n12972,
            clk => \N__56214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i21_LC_7_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__52632\,
            in1 => \N__40210\,
            in2 => \N__53193\,
            in3 => \N__36498\,
            lcout => encoder0_position_scaled_21,
            ltout => OPEN,
            carryin => n12972,
            carryout => n12973,
            clk => \N__56214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i22_LC_7_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__47745\,
            in1 => \N__49953\,
            in2 => \N__40231\,
            in3 => \N__36495\,
            lcout => encoder0_position_scaled_22,
            ltout => OPEN,
            carryin => n12973,
            carryout => n12974,
            clk => \N__56214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_scaled_i23_LC_7_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__38673\,
            in1 => \N__49881\,
            in2 => \N__40233\,
            in3 => \N__36651\,
            lcout => encoder0_position_scaled_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i15_1_lut_LC_7_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44121\,
            lcout => n11_adj_583,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12760_1_lut_LC_7_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36641\,
            lcout => n15490,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i10_1_lut_LC_7_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44270\,
            lcout => n16_adj_588,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i12_1_lut_LC_7_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44202\,
            lcout => n14_adj_586,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i9_1_lut_LC_7_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44310\,
            lcout => n17_adj_589,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_2_LC_7_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36617\,
            in2 => \N__54369\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_29_0_\,
            carryout => n12921,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_3_lut_LC_7_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36593\,
            in2 => \_gnd_net_\,
            in3 => \N__36561\,
            lcout => n3301,
            ltout => OPEN,
            carryin => n12921,
            carryout => n12922,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_4_lut_LC_7_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54074\,
            in2 => \N__36557\,
            in3 => \N__36534\,
            lcout => n3300,
            ltout => OPEN,
            carryin => n12922,
            carryout => n12923,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_5_lut_LC_7_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36903\,
            in3 => \N__36873\,
            lcout => n3299,
            ltout => OPEN,
            carryin => n12923,
            carryout => n12924,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_6_lut_LC_7_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54075\,
            in2 => \N__36870\,
            in3 => \N__36846\,
            lcout => n3298,
            ltout => OPEN,
            carryin => n12924,
            carryout => n12925,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_7_lut_LC_7_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__36843\,
            in1 => \_gnd_net_\,
            in2 => \N__36837\,
            in3 => \N__36804\,
            lcout => n15079,
            ltout => OPEN,
            carryin => n12925,
            carryout => n12926,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_8_lut_LC_7_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36800\,
            in3 => \N__36762\,
            lcout => n3296,
            ltout => OPEN,
            carryin => n12926,
            carryout => n12927,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_9_lut_LC_7_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53982\,
            in2 => \N__36759\,
            in3 => \N__36726\,
            lcout => n3295,
            ltout => OPEN,
            carryin => n12927,
            carryout => n12928,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_10_lut_LC_7_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53975\,
            in2 => \N__36723\,
            in3 => \N__36684\,
            lcout => n3294,
            ltout => OPEN,
            carryin => \bfn_7_30_0_\,
            carryout => n12929,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_11_lut_LC_7_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54021\,
            in2 => \N__36681\,
            in3 => \N__36654\,
            lcout => n3293,
            ltout => OPEN,
            carryin => n12929,
            carryout => n12930,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_12_lut_LC_7_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53976\,
            in2 => \N__37212\,
            in3 => \N__37179\,
            lcout => n3292,
            ltout => OPEN,
            carryin => n12930,
            carryout => n12931,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_13_lut_LC_7_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54022\,
            in2 => \N__37176\,
            in3 => \N__37143\,
            lcout => n3291,
            ltout => OPEN,
            carryin => n12931,
            carryout => n12932,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_14_lut_LC_7_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53977\,
            in2 => \N__37140\,
            in3 => \N__37101\,
            lcout => n3290,
            ltout => OPEN,
            carryin => n12932,
            carryout => n12933,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_15_lut_LC_7_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54023\,
            in2 => \N__37098\,
            in3 => \N__37062\,
            lcout => n3289,
            ltout => OPEN,
            carryin => n12933,
            carryout => n12934,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_16_lut_LC_7_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53978\,
            in2 => \N__37059\,
            in3 => \N__37026\,
            lcout => n3288,
            ltout => OPEN,
            carryin => n12934,
            carryout => n12935,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_17_lut_LC_7_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54024\,
            in2 => \N__37023\,
            in3 => \N__36990\,
            lcout => n3287,
            ltout => OPEN,
            carryin => n12935,
            carryout => n12936,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_18_lut_LC_7_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53968\,
            in2 => \N__36987\,
            in3 => \N__36939\,
            lcout => n3286,
            ltout => OPEN,
            carryin => \bfn_7_31_0_\,
            carryout => n12937,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_19_lut_LC_7_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54010\,
            in2 => \N__36936\,
            in3 => \N__36906\,
            lcout => n3285,
            ltout => OPEN,
            carryin => n12937,
            carryout => n12938,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_20_lut_LC_7_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37473\,
            in2 => \N__54414\,
            in3 => \N__37440\,
            lcout => n3284,
            ltout => OPEN,
            carryin => n12938,
            carryout => n12939,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_21_lut_LC_7_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37437\,
            in2 => \N__54367\,
            in3 => \N__37407\,
            lcout => n3283,
            ltout => OPEN,
            carryin => n12939,
            carryout => n12940,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_22_lut_LC_7_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37404\,
            in2 => \N__54415\,
            in3 => \N__37377\,
            lcout => n3282,
            ltout => OPEN,
            carryin => n12940,
            carryout => n12941,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_23_lut_LC_7_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37373\,
            in2 => \N__54368\,
            in3 => \N__37344\,
            lcout => n3281,
            ltout => OPEN,
            carryin => n12941,
            carryout => n12942,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_24_lut_LC_7_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37340\,
            in2 => \N__54416\,
            in3 => \N__37311\,
            lcout => n3280,
            ltout => OPEN,
            carryin => n12942,
            carryout => n12943,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_25_lut_LC_7_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54020\,
            in2 => \N__37308\,
            in3 => \N__37284\,
            lcout => n3279,
            ltout => OPEN,
            carryin => n12943,
            carryout => n12944,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_26_lut_LC_7_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37281\,
            in2 => \N__53646\,
            in3 => \N__37251\,
            lcout => n3278,
            ltout => OPEN,
            carryin => \bfn_7_32_0_\,
            carryout => n12945,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_27_lut_LC_7_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37248\,
            in2 => \N__53917\,
            in3 => \N__37215\,
            lcout => n3277,
            ltout => OPEN,
            carryin => n12945,
            carryout => n12946,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_28_lut_LC_7_32_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37755\,
            in2 => \N__53647\,
            in3 => \N__37719\,
            lcout => n3276,
            ltout => OPEN,
            carryin => n12946,
            carryout => n12947,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_29_lut_LC_7_32_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37715\,
            in2 => \N__53918\,
            in3 => \N__37680\,
            lcout => n3275,
            ltout => OPEN,
            carryin => n12947,
            carryout => n12948,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_30_lut_LC_7_32_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37677\,
            in2 => \N__53648\,
            in3 => \N__37644\,
            lcout => n3274,
            ltout => OPEN,
            carryin => n12948,
            carryout => n12949,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_31_lut_LC_7_32_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37640\,
            in2 => \N__53919\,
            in3 => \N__37602\,
            lcout => n3273,
            ltout => OPEN,
            carryin => n12949,
            carryout => n12950,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_32_lut_LC_7_32_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37594\,
            in2 => \N__53649\,
            in3 => \N__37557\,
            lcout => n3272,
            ltout => OPEN,
            carryin => n12950,
            carryout => n12951,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_2173_33_lut_LC_7_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__53659\,
            in1 => \N__37549\,
            in2 => \_gnd_net_\,
            in3 => \N__37524\,
            lcout => n3271,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_2_lut_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38107\,
            in2 => \_gnd_net_\,
            in3 => \N__37494\,
            lcout => n2001,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => n12622,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_3_lut_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55209\,
            in2 => \N__39313\,
            in3 => \N__37476\,
            lcout => n2000,
            ltout => OPEN,
            carryin => n12622,
            carryout => n12623,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_4_lut_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39535\,
            in3 => \N__37869\,
            lcout => n1999,
            ltout => OPEN,
            carryin => n12623,
            carryout => n12624,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_5_lut_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55210\,
            in2 => \N__39349\,
            in3 => \N__37857\,
            lcout => n1998,
            ltout => OPEN,
            carryin => n12624,
            carryout => n12625,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_6_lut_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39118\,
            in3 => \N__37839\,
            lcout => n1997,
            ltout => OPEN,
            carryin => n12625,
            carryout => n12626,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_7_lut_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39281\,
            in3 => \N__37821\,
            lcout => n1996,
            ltout => OPEN,
            carryin => n12626,
            carryout => n12627,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_8_lut_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55218\,
            in2 => \N__39242\,
            in3 => \N__37803\,
            lcout => n1995,
            ltout => OPEN,
            carryin => n12627,
            carryout => n12628,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_9_lut_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55211\,
            in2 => \N__41744\,
            in3 => \N__37788\,
            lcout => n1994,
            ltout => OPEN,
            carryin => n12628,
            carryout => n12629,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_10_lut_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55203\,
            in2 => \N__41702\,
            in3 => \N__37773\,
            lcout => n1993,
            ltout => OPEN,
            carryin => \bfn_9_17_0_\,
            carryout => n12630,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_11_lut_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55212\,
            in2 => \N__39608\,
            in3 => \N__37758\,
            lcout => n1992,
            ltout => OPEN,
            carryin => n12630,
            carryout => n12631,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_12_lut_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55204\,
            in2 => \N__41133\,
            in3 => \N__38052\,
            lcout => n1991,
            ltout => OPEN,
            carryin => n12631,
            carryout => n12632,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_13_lut_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55213\,
            in2 => \N__39578\,
            in3 => \N__38037\,
            lcout => n1990,
            ltout => OPEN,
            carryin => n12632,
            carryout => n12633,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_14_lut_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55205\,
            in2 => \N__38034\,
            in3 => \N__38007\,
            lcout => n1989,
            ltout => OPEN,
            carryin => n12633,
            carryout => n12634,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_15_lut_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55214\,
            in2 => \N__37907\,
            in3 => \N__37992\,
            lcout => n1988,
            ltout => OPEN,
            carryin => n12634,
            carryout => n12635,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_16_lut_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41421\,
            in2 => \N__55393\,
            in3 => \N__37989\,
            lcout => n1987,
            ltout => OPEN,
            carryin => n12635,
            carryout => n12636,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_17_lut_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38137\,
            in2 => \N__55392\,
            in3 => \N__37971\,
            lcout => n1986,
            ltout => OPEN,
            carryin => n12636,
            carryout => n12637,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_18_lut_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38158\,
            in2 => \N__55340\,
            in3 => \N__37956\,
            lcout => n1985,
            ltout => OPEN,
            carryin => \bfn_9_18_0_\,
            carryout => n12638,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1302_19_lut_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__41637\,
            in1 => \N__55151\,
            in2 => \N__37953\,
            in3 => \N__37932\,
            lcout => n2016,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1241_3_lut_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41091\,
            in2 => \N__41193\,
            in3 => \N__41495\,
            lcout => n1921,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_143_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39122\,
            in3 => \N__39280\,
            lcout => n14530,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1238_3_lut_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41229\,
            in2 => \N__41160\,
            in3 => \N__41497\,
            lcout => n1918,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1239_3_lut_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43194\,
            in2 => \N__41175\,
            in3 => \N__41496\,
            lcout => n1919,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39469\,
            lcout => n31_adj_649,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39403\,
            lcout => n28_adj_646,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i15_3_lut_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49589\,
            in1 => \N__38598\,
            in2 => \_gnd_net_\,
            in3 => \N__39632\,
            lcout => n305,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39506\,
            in3 => \_gnd_net_\,
            lcout => n33_adj_651,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i14_3_lut_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38625\,
            in1 => \N__49590\,
            in2 => \_gnd_net_\,
            in3 => \N__39928\,
            lcout => n306,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i16_3_lut_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__39827\,
            in1 => \_gnd_net_\,
            in2 => \N__49580\,
            in3 => \N__38574\,
            lcout => n304,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i20_3_lut_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38538\,
            in1 => \N__49513\,
            in2 => \_gnd_net_\,
            in3 => \N__39799\,
            lcout => n300,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39631\,
            lcout => n19_adj_637,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39826\,
            lcout => n18_adj_636,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39664\,
            lcout => n23_adj_641,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39727\,
            in3 => \_gnd_net_\,
            lcout => n25_adj_643,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i12_3_lut_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49517\,
            in1 => \N__38376\,
            in2 => \_gnd_net_\,
            in3 => \N__40000\,
            lcout => n308,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39691\,
            lcout => n24_adj_642,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39760\,
            lcout => n26_adj_644,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39801\,
            in3 => \_gnd_net_\,
            lcout => n14_adj_632,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41596\,
            lcout => n30_adj_648,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39380\,
            lcout => n27_adj_645,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i11_3_lut_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38388\,
            in1 => \N__49538\,
            in2 => \_gnd_net_\,
            in3 => \N__39671\,
            lcout => n309,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41949\,
            lcout => n4_adj_622,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39440\,
            lcout => n29_adj_647,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_2_lut_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38313\,
            in3 => \N__38289\,
            lcout => n33,
            ltout => OPEN,
            carryin => \bfn_9_22_0_\,
            carryout => n12975,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_3_lut_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45771\,
            in3 => \N__38277\,
            lcout => n32,
            ltout => OPEN,
            carryin => n12975,
            carryout => n12976,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_4_lut_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38274\,
            in3 => \N__38250\,
            lcout => n31,
            ltout => OPEN,
            carryin => n12976,
            carryout => n12977,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_5_lut_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38247\,
            in3 => \N__38238\,
            lcout => n30,
            ltout => OPEN,
            carryin => n12977,
            carryout => n12978,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_6_lut_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38235\,
            in3 => \N__38214\,
            lcout => n29,
            ltout => OPEN,
            carryin => n12978,
            carryout => n12979,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_7_lut_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38523\,
            in3 => \N__38502\,
            lcout => n28,
            ltout => OPEN,
            carryin => n12979,
            carryout => n12980,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_8_lut_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38499\,
            in3 => \N__38481\,
            lcout => n27,
            ltout => OPEN,
            carryin => n12980,
            carryout => n12981,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_9_lut_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38478\,
            in3 => \N__38457\,
            lcout => n26,
            ltout => OPEN,
            carryin => n12981,
            carryout => n12982,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_10_lut_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38454\,
            in3 => \N__38430\,
            lcout => n25,
            ltout => OPEN,
            carryin => \bfn_9_23_0_\,
            carryout => n12983,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_11_lut_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38427\,
            in3 => \N__38403\,
            lcout => n24,
            ltout => OPEN,
            carryin => n12983,
            carryout => n12984,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_12_lut_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38400\,
            in3 => \N__38379\,
            lcout => n23,
            ltout => OPEN,
            carryin => n12984,
            carryout => n12985,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_13_lut_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39981\,
            in3 => \N__38367\,
            lcout => n22,
            ltout => OPEN,
            carryin => n12985,
            carryout => n12986,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_14_lut_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39939\,
            in3 => \N__38352\,
            lcout => n21,
            ltout => OPEN,
            carryin => n12986,
            carryout => n12987,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_15_lut_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39909\,
            in3 => \N__38613\,
            lcout => n20,
            ltout => OPEN,
            carryin => n12987,
            carryout => n12988,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_16_lut_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38610\,
            in3 => \N__38589\,
            lcout => n19,
            ltout => OPEN,
            carryin => n12988,
            carryout => n12989,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_17_lut_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38586\,
            in3 => \N__38562\,
            lcout => n18,
            ltout => OPEN,
            carryin => n12989,
            carryout => n12990,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_18_lut_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45732\,
            in3 => \N__38559\,
            lcout => n17,
            ltout => OPEN,
            carryin => \bfn_9_24_0_\,
            carryout => n12991,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_19_lut_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41904\,
            in3 => \N__38556\,
            lcout => n16,
            ltout => OPEN,
            carryin => n12991,
            carryout => n12992,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_20_lut_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40326\,
            in3 => \N__38553\,
            lcout => n15,
            ltout => OPEN,
            carryin => n12992,
            carryout => n12993,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_21_lut_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38550\,
            in3 => \N__38529\,
            lcout => n14,
            ltout => OPEN,
            carryin => n12993,
            carryout => n12994,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_22_lut_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39864\,
            in3 => \N__38526\,
            lcout => n13,
            ltout => OPEN,
            carryin => n12994,
            carryout => n12995,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_23_lut_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__52389\,
            in3 => \N__38664\,
            lcout => n12,
            ltout => OPEN,
            carryin => n12995,
            carryout => n12996,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_24_lut_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45645\,
            in3 => \N__38661\,
            lcout => n11,
            ltout => OPEN,
            carryin => n12996,
            carryout => n12997,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_25_lut_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43719\,
            in3 => \N__38658\,
            lcout => n10,
            ltout => OPEN,
            carryin => n12997,
            carryout => n12998,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_26_lut_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40065\,
            in3 => \N__38655\,
            lcout => n9,
            ltout => OPEN,
            carryin => \bfn_9_25_0_\,
            carryout => n12999,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_27_lut_LC_9_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40251\,
            in3 => \N__38652\,
            lcout => n8,
            ltout => OPEN,
            carryin => n12999,
            carryout => n13000,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_28_lut_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41889\,
            in3 => \N__38649\,
            lcout => n7,
            ltout => OPEN,
            carryin => n13000,
            carryout => n13001,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_29_lut_LC_9_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40317\,
            in3 => \N__38646\,
            lcout => n6,
            ltout => OPEN,
            carryin => n13001,
            carryout => n13002,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_30_lut_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40242\,
            in3 => \N__38643\,
            lcout => n5,
            ltout => OPEN,
            carryin => n13002,
            carryout => n13003,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_31_lut_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38640\,
            in2 => \_gnd_net_\,
            in3 => \N__38628\,
            lcout => n4,
            ltout => OPEN,
            carryin => n13003,
            carryout => n13004,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_32_lut_LC_9_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41874\,
            in3 => \N__38733\,
            lcout => n3,
            ltout => OPEN,
            carryin => n13004,
            carryout => n13005,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_add_3_33_lut_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40083\,
            in2 => \_gnd_net_\,
            in3 => \N__38730\,
            lcout => n2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i9_1_lut_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38727\,
            lcout => n17_adj_559,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i11_1_lut_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44231\,
            lcout => n15_adj_587,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i15_1_lut_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38718\,
            lcout => n11_adj_565,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i11_1_lut_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38709\,
            lcout => n15_adj_561,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i13_1_lut_LC_9_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38700\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n13_adj_563,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i14_1_lut_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38691\,
            lcout => n12_adj_564,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i16_1_lut_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38682\,
            lcout => n10_adj_566,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12778_1_lut_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49877\,
            lcout => n15508,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i19_1_lut_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38763\,
            lcout => n7_adj_569,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9552_2_lut_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__46659\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46615\,
            lcout => n11526,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9553_1_lut_2_lut_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46614\,
            in2 => \_gnd_net_\,
            in3 => \N__46658\,
            lcout => n1377,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i24_1_lut_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38754\,
            lcout => n2_adj_574,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i18_1_lut_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38745\,
            lcout => n8_adj_568,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i17_1_lut_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44450\,
            lcout => n9_adj_581,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12768_2_lut_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46616\,
            in2 => \_gnd_net_\,
            in3 => \N__46660\,
            lcout => OPEN,
            ltout => \dti_N_333_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111101111"
        )
    port map (
            in0 => \N__39188\,
            in1 => \N__46692\,
            in2 => \N__38736\,
            in3 => \N__56517\,
            lcout => n5187,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12403_2_lut_4_lut_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000010000"
        )
    port map (
            in0 => \N__46693\,
            in1 => \N__56518\,
            in2 => \N__39077\,
            in3 => \N__39189\,
            lcout => n15072,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \debounce.reg_out_i0_i1_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46988\,
            in1 => \N__38895\,
            in2 => \_gnd_net_\,
            in3 => \N__38874\,
            lcout => h2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_662__i0_LC_9_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__38985\,
            in1 => \N__39002\,
            in2 => \N__38841\,
            in3 => \N__38829\,
            lcout => dti_counter_0,
            ltout => OPEN,
            carryin => \bfn_9_29_0_\,
            carryout => n13006,
            clk => \N__56223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_662__i1_LC_9_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__39198\,
            in1 => \N__38787\,
            in2 => \N__39224\,
            in3 => \N__38826\,
            lcout => dti_counter_1,
            ltout => OPEN,
            carryin => n13006,
            carryout => n13007,
            clk => \N__56223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_662__i2_LC_9_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__39090\,
            in1 => \N__39027\,
            in2 => \N__38800\,
            in3 => \N__38823\,
            lcout => dti_counter_2,
            ltout => OPEN,
            carryin => n13007,
            carryout => n13008,
            clk => \N__56223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_662__i3_LC_9_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__38961\,
            in1 => \N__38791\,
            in2 => \N__38979\,
            in3 => \N__38820\,
            lcout => dti_counter_3,
            ltout => OPEN,
            carryin => n13008,
            carryout => n13009,
            clk => \N__56223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_662__i4_LC_9_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__38937\,
            in1 => \N__38954\,
            in2 => \N__38801\,
            in3 => \N__38817\,
            lcout => dti_counter_4,
            ltout => OPEN,
            carryin => n13009,
            carryout => n13010,
            clk => \N__56223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_662__i5_LC_9_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__38814\,
            in1 => \N__38795\,
            in2 => \N__39078\,
            in3 => \N__38808\,
            lcout => dti_counter_5,
            ltout => OPEN,
            carryin => n13010,
            carryout => n13011,
            clk => \N__56223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_662__i6_LC_9_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__39084\,
            in1 => \N__39052\,
            in2 => \N__38802\,
            in3 => \N__38805\,
            lcout => dti_counter_6,
            ltout => OPEN,
            carryin => n13011,
            carryout => n13012,
            clk => \N__56223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_counter_662__i7_LC_9_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100001110100"
        )
    port map (
            in0 => \N__38927\,
            in1 => \N__38799\,
            in2 => \N__38907\,
            in3 => \N__38766\,
            lcout => dti_counter_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12406_2_lut_4_lut_LC_9_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100000000"
        )
    port map (
            in0 => \N__39184\,
            in1 => \N__56522\,
            in2 => \N__46722\,
            in3 => \N__39026\,
            lcout => n15075,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12390_2_lut_4_lut_LC_9_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010010000"
        )
    port map (
            in0 => \N__56519\,
            in1 => \N__39185\,
            in2 => \N__39054\,
            in3 => \N__46718\,
            lcout => n15071,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_79_LC_9_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39070\,
            in1 => \N__38950\,
            in2 => \N__39053\,
            in3 => \N__38923\,
            lcout => OPEN,
            ltout => \n14_adj_705_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_LC_9_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38974\,
            in1 => \N__39001\,
            in2 => \N__39030\,
            in3 => \N__39012\,
            lcout => n5137,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_adj_78_LC_9_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39214\,
            in2 => \_gnd_net_\,
            in3 => \N__39025\,
            lcout => n10_adj_706,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12360_2_lut_4_lut_LC_9_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010010000"
        )
    port map (
            in0 => \N__56523\,
            in1 => \N__39187\,
            in2 => \N__39006\,
            in3 => \N__46720\,
            lcout => n15081,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12405_2_lut_4_lut_LC_9_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100000000"
        )
    port map (
            in0 => \N__39183\,
            in1 => \N__56521\,
            in2 => \N__46721\,
            in3 => \N__38975\,
            lcout => n15074,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12404_2_lut_4_lut_LC_9_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010010000"
        )
    port map (
            in0 => \N__56520\,
            in1 => \N__39186\,
            in2 => \N__38955\,
            in3 => \N__46719\,
            lcout => n15073,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12418_2_lut_4_lut_LC_9_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000010000"
        )
    port map (
            in0 => \N__56509\,
            in1 => \N__46711\,
            in2 => \N__38931\,
            in3 => \N__39182\,
            lcout => n15070,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_3_lut_LC_9_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111101110"
        )
    port map (
            in0 => \N__47000\,
            in1 => \N__46955\,
            in2 => \_gnd_net_\,
            in3 => \N__46892\,
            lcout => n6_adj_721,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12199_4_lut_LC_9_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011011000"
        )
    port map (
            in0 => \N__40764\,
            in1 => \N__40784\,
            in2 => \N__40746\,
            in3 => \N__40992\,
            lcout => n14929,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12198_4_lut_LC_9_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011010000"
        )
    port map (
            in0 => \N__40991\,
            in1 => \N__40763\,
            in2 => \N__40785\,
            in3 => \N__40742\,
            lcout => n14928,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12407_2_lut_4_lut_LC_9_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000010000"
        )
    port map (
            in0 => \N__56508\,
            in1 => \N__46710\,
            in2 => \N__39225\,
            in3 => \N__39181\,
            lcout => n15076,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \commutation_state_prev_i0_LC_9_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56510\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => commutation_state_prev_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56235\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i18_LC_9_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50899\,
            in1 => \N__44553\,
            in2 => \_gnd_net_\,
            in3 => \N__42669\,
            lcout => pwm_setpoint_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56241\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12200_3_lut_LC_9_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__40971\,
            in1 => \N__39150\,
            in2 => \_gnd_net_\,
            in3 => \N__39144\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1183_3_lut_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43287\,
            in2 => \N__43317\,
            in3 => \N__45500\,
            lcout => n1831,
            ltout => \n1831_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1250_3_lut_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40836\,
            in2 => \N__39126\,
            in3 => \N__41490\,
            lcout => n1930,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1251_3_lut_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40883\,
            in2 => \N__40863\,
            in3 => \N__41494\,
            lcout => n1931,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1253_3_lut_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40950\,
            in2 => \N__41514\,
            in3 => \N__40920\,
            lcout => n1933,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1249_3_lut_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41055\,
            in2 => \N__43119\,
            in3 => \N__41489\,
            lcout => n1929,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1243_3_lut_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__43057\,
            in1 => \_gnd_net_\,
            in2 => \N__41019\,
            in3 => \N__41482\,
            lcout => n1923,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1245_3_lut_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43083\,
            in2 => \N__41512\,
            in3 => \N__41031\,
            lcout => n1925,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_137_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43027\,
            in2 => \N__43059\,
            in3 => \N__42858\,
            lcout => OPEN,
            ltout => \n14524_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_138_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__41665\,
            in1 => \N__43112\,
            in2 => \N__39255\,
            in3 => \N__40956\,
            lcout => OPEN,
            ltout => \n14526_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12925_4_lut_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41227\,
            in1 => \N__41067\,
            in2 => \N__39252\,
            in3 => \N__43748\,
            lcout => n1851,
            ltout => \n1851_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1248_3_lut_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__41666\,
            in1 => \_gnd_net_\,
            in2 => \N__39249\,
            in3 => \N__41046\,
            lcout => n1928,
            ltout => \n1928_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_141_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39601\,
            in2 => \N__39585\,
            in3 => \N__39571\,
            lcout => n14440,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1252_3_lut_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40893\,
            in2 => \N__41513\,
            in3 => \N__40911\,
            lcout => n1932,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i0_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39505\,
            in2 => \_gnd_net_\,
            in3 => \N__39483\,
            lcout => encoder0_position_0,
            ltout => OPEN,
            carryin => \bfn_10_18_0_\,
            carryout => \quad_counter0.n13095\,
            clk => \N__56201\,
            ce => \N__40308\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i1_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40455\,
            in2 => \N__45799\,
            in3 => \N__39480\,
            lcout => encoder0_position_1,
            ltout => OPEN,
            carryin => \quad_counter0.n13095\,
            carryout => \quad_counter0.n13096\,
            clk => \N__56201\,
            ce => \N__40308\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i2_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39473\,
            in2 => \N__40514\,
            in3 => \N__39453\,
            lcout => encoder0_position_2,
            ltout => OPEN,
            carryin => \quad_counter0.n13096\,
            carryout => \quad_counter0.n13097\,
            clk => \N__56201\,
            ce => \N__40308\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i3_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40459\,
            in2 => \N__41600\,
            in3 => \N__39450\,
            lcout => encoder0_position_3,
            ltout => OPEN,
            carryin => \quad_counter0.n13097\,
            carryout => \quad_counter0.n13098\,
            clk => \N__56201\,
            ce => \N__40308\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i4_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39439\,
            in2 => \N__40515\,
            in3 => \N__39417\,
            lcout => encoder0_position_4,
            ltout => OPEN,
            carryin => \quad_counter0.n13098\,
            carryout => \quad_counter0.n13099\,
            clk => \N__56201\,
            ce => \N__40308\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i5_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40463\,
            in2 => \N__39413\,
            in3 => \N__39387\,
            lcout => encoder0_position_5,
            ltout => OPEN,
            carryin => \quad_counter0.n13099\,
            carryout => \quad_counter0.n13100\,
            clk => \N__56201\,
            ce => \N__40308\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i6_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39379\,
            in2 => \N__40516\,
            in3 => \N__39357\,
            lcout => encoder0_position_6,
            ltout => OPEN,
            carryin => \quad_counter0.n13100\,
            carryout => \quad_counter0.n13101\,
            clk => \N__56201\,
            ce => \N__40308\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i7_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40467\,
            in2 => \N__39764\,
            in3 => \N__39738\,
            lcout => encoder0_position_7,
            ltout => OPEN,
            carryin => \quad_counter0.n13101\,
            carryout => \quad_counter0.n13102\,
            clk => \N__56201\,
            ce => \N__40308\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i8_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40468\,
            in2 => \N__39731\,
            in3 => \N__39702\,
            lcout => encoder0_position_8,
            ltout => OPEN,
            carryin => \bfn_10_19_0_\,
            carryout => \quad_counter0.n13103\,
            clk => \N__56202\,
            ce => \N__40303\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i9_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39695\,
            in2 => \N__40517\,
            in3 => \N__39675\,
            lcout => encoder0_position_9,
            ltout => OPEN,
            carryin => \quad_counter0.n13103\,
            carryout => \quad_counter0.n13104\,
            clk => \N__56202\,
            ce => \N__40303\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i10_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40472\,
            in2 => \N__39672\,
            in3 => \N__39648\,
            lcout => encoder0_position_10,
            ltout => OPEN,
            carryin => \quad_counter0.n13104\,
            carryout => \quad_counter0.n13105\,
            clk => \N__56202\,
            ce => \N__40303\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i11_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40001\,
            in2 => \N__40518\,
            in3 => \N__39645\,
            lcout => encoder0_position_11,
            ltout => OPEN,
            carryin => \quad_counter0.n13105\,
            carryout => \quad_counter0.n13106\,
            clk => \N__56202\,
            ce => \N__40303\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i12_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40476\,
            in2 => \N__39970\,
            in3 => \N__39642\,
            lcout => encoder0_position_12,
            ltout => OPEN,
            carryin => \quad_counter0.n13106\,
            carryout => \quad_counter0.n13107\,
            clk => \N__56202\,
            ce => \N__40303\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i13_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39929\,
            in2 => \N__40519\,
            in3 => \N__39639\,
            lcout => encoder0_position_13,
            ltout => OPEN,
            carryin => \quad_counter0.n13107\,
            carryout => \quad_counter0.n13108\,
            clk => \N__56202\,
            ce => \N__40303\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i14_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40480\,
            in2 => \N__39636\,
            in3 => \N__39615\,
            lcout => encoder0_position_14,
            ltout => OPEN,
            carryin => \quad_counter0.n13108\,
            carryout => \quad_counter0.n13109\,
            clk => \N__56202\,
            ce => \N__40303\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i15_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39828\,
            in2 => \N__40520\,
            in3 => \N__39813\,
            lcout => encoder0_position_15,
            ltout => OPEN,
            carryin => \quad_counter0.n13109\,
            carryout => \quad_counter0.n13110\,
            clk => \N__56202\,
            ce => \N__40303\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i16_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40484\,
            in2 => \N__45757\,
            in3 => \N__39810\,
            lcout => encoder0_position_16,
            ltout => OPEN,
            carryin => \bfn_10_20_0_\,
            carryout => \quad_counter0.n13111\,
            clk => \N__56205\,
            ce => \N__40304\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i17_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41919\,
            in2 => \N__40521\,
            in3 => \N__39807\,
            lcout => encoder0_position_17,
            ltout => OPEN,
            carryin => \quad_counter0.n13111\,
            carryout => \quad_counter0.n13112\,
            clk => \N__56205\,
            ce => \N__40304\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i18_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40488\,
            in2 => \N__43656\,
            in3 => \N__39804\,
            lcout => encoder0_position_18,
            ltout => OPEN,
            carryin => \quad_counter0.n13112\,
            carryout => \quad_counter0.n13113\,
            clk => \N__56205\,
            ce => \N__40304\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i19_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39800\,
            in2 => \N__40522\,
            in3 => \N__39780\,
            lcout => encoder0_position_19,
            ltout => OPEN,
            carryin => \quad_counter0.n13113\,
            carryout => \quad_counter0.n13114\,
            clk => \N__56205\,
            ce => \N__40304\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i20_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40492\,
            in2 => \N__47711\,
            in3 => \N__39777\,
            lcout => encoder0_position_20,
            ltout => OPEN,
            carryin => \quad_counter0.n13114\,
            carryout => \quad_counter0.n13115\,
            clk => \N__56205\,
            ce => \N__40304\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i21_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52408\,
            in2 => \N__40523\,
            in3 => \N__39774\,
            lcout => encoder0_position_21,
            ltout => OPEN,
            carryin => \quad_counter0.n13115\,
            carryout => \quad_counter0.n13116\,
            clk => \N__56205\,
            ce => \N__40304\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i22_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40496\,
            in2 => \N__47369\,
            in3 => \N__39771\,
            lcout => encoder0_position_22,
            ltout => OPEN,
            carryin => \quad_counter0.n13116\,
            carryout => \quad_counter0.n13117\,
            clk => \N__56205\,
            ce => \N__40304\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i23_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43837\,
            in2 => \N__40524\,
            in3 => \N__39768\,
            lcout => encoder0_position_23,
            ltout => OPEN,
            carryin => \quad_counter0.n13117\,
            carryout => \quad_counter0.n13118\,
            clk => \N__56205\,
            ce => \N__40304\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i24_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40500\,
            in2 => \N__43809\,
            in3 => \N__39855\,
            lcout => encoder0_position_24,
            ltout => OPEN,
            carryin => \bfn_10_21_0_\,
            carryout => \quad_counter0.n13119\,
            clk => \N__56206\,
            ce => \N__40302\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i25_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43909\,
            in2 => \N__40525\,
            in3 => \N__39852\,
            lcout => encoder0_position_25,
            ltout => OPEN,
            carryin => \quad_counter0.n13119\,
            carryout => \quad_counter0.n13120\,
            clk => \N__56206\,
            ce => \N__40302\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i26_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40504\,
            in2 => \N__41828\,
            in3 => \N__39849\,
            lcout => encoder0_position_26,
            ltout => OPEN,
            carryin => \quad_counter0.n13120\,
            carryout => \quad_counter0.n13121\,
            clk => \N__56206\,
            ce => \N__40302\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i27_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41785\,
            in2 => \N__40526\,
            in3 => \N__39846\,
            lcout => encoder0_position_27,
            ltout => OPEN,
            carryin => \quad_counter0.n13121\,
            carryout => \quad_counter0.n13122\,
            clk => \N__56206\,
            ce => \N__40302\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i28_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40508\,
            in2 => \N__42073\,
            in3 => \N__39843\,
            lcout => encoder0_position_28,
            ltout => OPEN,
            carryin => \quad_counter0.n13122\,
            carryout => \quad_counter0.n13123\,
            clk => \N__56206\,
            ce => \N__40302\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i29_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41954\,
            in2 => \N__40527\,
            in3 => \N__39840\,
            lcout => encoder0_position_29,
            ltout => OPEN,
            carryin => \quad_counter0.n13123\,
            carryout => \quad_counter0.n13124\,
            clk => \N__56206\,
            ce => \N__40302\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i30_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40512\,
            in2 => \N__42019\,
            in3 => \N__39837\,
            lcout => encoder0_position_30,
            ltout => OPEN,
            carryin => \quad_counter0.n13124\,
            carryout => \quad_counter0.n13125\,
            clk => \N__56206\,
            ce => \N__40302\,
            sr => \_gnd_net_\
        );

    \quad_counter0.position_659__i31_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__40513\,
            in1 => \N__49540\,
            in2 => \_gnd_net_\,
            in3 => \N__39834\,
            lcout => encoder0_position_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56206\,
            ce => \N__40302\,
            sr => \_gnd_net_\
        );

    \add_741_2_lut_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42282\,
            in3 => \N__39831\,
            lcout => n2566,
            ltout => OPEN,
            carryin => \bfn_10_22_0_\,
            carryout => n12496,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_741_3_lut_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54700\,
            in2 => \N__40029\,
            in3 => \N__39900\,
            lcout => n2565,
            ltout => OPEN,
            carryin => n12496,
            carryout => n12497,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_741_4_lut_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40047\,
            in3 => \N__39897\,
            lcout => n2564,
            ltout => OPEN,
            carryin => n12497,
            carryout => n12498,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_741_5_lut_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54701\,
            in2 => \N__41928\,
            in3 => \N__39894\,
            lcout => n2563,
            ltout => OPEN,
            carryin => n12498,
            carryout => n12499,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_741_6_lut_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__39873\,
            in3 => \N__39891\,
            lcout => n2562,
            ltout => OPEN,
            carryin => n12499,
            carryout => n12500,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_741_7_lut_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40038\,
            in3 => \N__39888\,
            lcout => n2561,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10984_3_lut_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49496\,
            in2 => \N__41955\,
            in3 => \N__39879\,
            lcout => n830,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10983_3_lut_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42193\,
            in2 => \N__42318\,
            in3 => \N__39885\,
            lcout => n13656,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i31_3_lut_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__49547\,
            in1 => \_gnd_net_\,
            in2 => \N__42020\,
            in3 => \N__42220\,
            lcout => n403,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i27_3_lut_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49542\,
            in2 => \N__41829\,
            in3 => \N__41846\,
            lcout => n40,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47707\,
            lcout => n13_adj_631,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i29_3_lut_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49546\,
            in2 => \N__42075\,
            in3 => \N__42256\,
            lcout => n38,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_152_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42231\,
            in2 => \N__49598\,
            in3 => \N__42221\,
            lcout => n14568,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2181_2_lut_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49548\,
            in2 => \_gnd_net_\,
            in3 => \N__42428\,
            lcout => n402,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i28_3_lut_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41787\,
            in2 => \N__49597\,
            in3 => \N__42340\,
            lcout => n39,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10981_3_lut_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42194\,
            in2 => \N__42225\,
            in3 => \N__40020\,
            lcout => n13654,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dti_163_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46601\,
            in2 => \_gnd_net_\,
            in3 => \N__46665\,
            lcout => dti,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56212\,
            ce => \N__40014\,
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40002\,
            lcout => n22_adj_640,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39971\,
            lcout => n21_adj_639,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39930\,
            lcout => n20_adj_638,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43648\,
            lcout => n15_adj_633,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41786\,
            lcout => n6_adj_624,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.debounce_cnt_I_0_4_lut_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010101000"
        )
    port map (
            in0 => \N__46306\,
            in1 => \N__40362\,
            in2 => \N__46401\,
            in3 => \N__40542\,
            lcout => \direction_N_537\,
            ltout => \direction_N_537_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.direction_57_LC_10_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110010101100"
        )
    port map (
            in0 => \N__46400\,
            in1 => \N__40257\,
            in2 => \N__40260\,
            in3 => \N__46278\,
            lcout => n1302,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56215\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43916\,
            lcout => n8_adj_626,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut_LC_10_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42074\,
            in3 => \_gnd_net_\,
            lcout => n5_adj_623,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49541\,
            lcout => n2_adj_620,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43801\,
            lcout => n9_adj_627,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i6_1_lut_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40056\,
            lcout => n20_adj_556,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i2_1_lut_LC_10_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40371\,
            lcout => n24_adj_552,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i8_3_lut_3_lut_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__42803\,
            in1 => \N__47979\,
            in2 => \_gnd_net_\,
            in3 => \N__40563\,
            lcout => n8_adj_657,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_prev_I_0_65_2_lut_LC_10_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46340\,
            in2 => \_gnd_net_\,
            in3 => \N__46277\,
            lcout => \quad_counter0.direction_N_540\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i10_1_lut_LC_10_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40356\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n16_adj_560,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i5_LC_10_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43968\,
            in1 => \N__42459\,
            in2 => \_gnd_net_\,
            in3 => \N__50907\,
            lcout => pwm_setpoint_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i21_1_lut_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40347\,
            lcout => n5_adj_571,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i7_LC_10_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42441\,
            in1 => \N__50908\,
            in2 => \_gnd_net_\,
            in3 => \N__44340\,
            lcout => pwm_setpoint_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i4_LC_10_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50906\,
            in1 => \N__42474\,
            in2 => \_gnd_net_\,
            in3 => \N__43998\,
            lcout => pwm_setpoint_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i12_1_lut_LC_10_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40335\,
            lcout => n14_adj_562,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i13_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50868\,
            in1 => \N__44151\,
            in2 => \_gnd_net_\,
            in3 => \N__42558\,
            lcout => pwm_setpoint_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i22_1_lut_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40581\,
            lcout => n4_adj_572,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i20_1_lut_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40572\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n6_adj_570,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i9_2_lut_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40562\,
            in2 => \_gnd_net_\,
            in3 => \N__48102\,
            lcout => n9_adj_658,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i23_1_lut_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40551\,
            lcout => n3_adj_573,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i14_1_lut_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44150\,
            lcout => n12_adj_584,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i11_LC_10_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50867\,
            in1 => \N__44201\,
            in2 => \_gnd_net_\,
            in3 => \N__42576\,
            lcout => pwm_setpoint_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i8_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44309\,
            in1 => \N__42627\,
            in2 => \_gnd_net_\,
            in3 => \N__50869\,
            lcout => pwm_setpoint_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.a_prev_51_LC_10_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__46395\,
            in1 => \N__40541\,
            in2 => \N__46308\,
            in3 => \N__46356\,
            lcout => \quad_counter0.a_prev\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56220\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_prev_I_0_63_2_lut_LC_10_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46394\,
            in2 => \_gnd_net_\,
            in3 => \N__46270\,
            lcout => \quad_counter0.direction_N_536\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.debounce_cnt_50_LC_10_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__46396\,
            in1 => \N__46457\,
            in2 => \N__46347\,
            in3 => \N__46428\,
            lcout => \quad_counter0.debounce_cnt\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56220\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i0_LC_10_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40644\,
            in2 => \_gnd_net_\,
            in3 => \N__40638\,
            lcout => n26_adj_703,
            ltout => OPEN,
            carryin => \bfn_10_29_0_\,
            carryout => n13070,
            clk => \N__56224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i1_LC_10_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40635\,
            in2 => \_gnd_net_\,
            in3 => \N__40629\,
            lcout => n25_adj_702,
            ltout => OPEN,
            carryin => n13070,
            carryout => n13071,
            clk => \N__56224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i2_LC_10_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40626\,
            in2 => \_gnd_net_\,
            in3 => \N__40620\,
            lcout => n24_adj_701,
            ltout => OPEN,
            carryin => n13071,
            carryout => n13072,
            clk => \N__56224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i3_LC_10_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40617\,
            in2 => \_gnd_net_\,
            in3 => \N__40611\,
            lcout => n23_adj_700,
            ltout => OPEN,
            carryin => n13072,
            carryout => n13073,
            clk => \N__56224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i4_LC_10_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40608\,
            in2 => \_gnd_net_\,
            in3 => \N__40602\,
            lcout => n22_adj_699,
            ltout => OPEN,
            carryin => n13073,
            carryout => n13074,
            clk => \N__56224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i5_LC_10_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40599\,
            in2 => \_gnd_net_\,
            in3 => \N__40593\,
            lcout => n21_adj_698,
            ltout => OPEN,
            carryin => n13074,
            carryout => n13075,
            clk => \N__56224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i6_LC_10_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40590\,
            in2 => \_gnd_net_\,
            in3 => \N__40584\,
            lcout => n20_adj_697,
            ltout => OPEN,
            carryin => n13075,
            carryout => n13076,
            clk => \N__56224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i7_LC_10_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40725\,
            in2 => \_gnd_net_\,
            in3 => \N__40719\,
            lcout => n19_adj_696,
            ltout => OPEN,
            carryin => n13076,
            carryout => n13077,
            clk => \N__56224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i8_LC_10_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40716\,
            in2 => \_gnd_net_\,
            in3 => \N__40710\,
            lcout => n18_adj_695,
            ltout => OPEN,
            carryin => \bfn_10_30_0_\,
            carryout => n13078,
            clk => \N__56229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i9_LC_10_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40707\,
            in2 => \_gnd_net_\,
            in3 => \N__40701\,
            lcout => n17_adj_694,
            ltout => OPEN,
            carryin => n13078,
            carryout => n13079,
            clk => \N__56229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i10_LC_10_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40698\,
            in2 => \_gnd_net_\,
            in3 => \N__40692\,
            lcout => n16_adj_693,
            ltout => OPEN,
            carryin => n13079,
            carryout => n13080,
            clk => \N__56229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i11_LC_10_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40689\,
            in2 => \_gnd_net_\,
            in3 => \N__40683\,
            lcout => n15_adj_692,
            ltout => OPEN,
            carryin => n13080,
            carryout => n13081,
            clk => \N__56229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i12_LC_10_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40680\,
            in2 => \_gnd_net_\,
            in3 => \N__40674\,
            lcout => n14_adj_691,
            ltout => OPEN,
            carryin => n13081,
            carryout => n13082,
            clk => \N__56229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i13_LC_10_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40671\,
            in2 => \_gnd_net_\,
            in3 => \N__40665\,
            lcout => n13_adj_690,
            ltout => OPEN,
            carryin => n13082,
            carryout => n13083,
            clk => \N__56229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i14_LC_10_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40662\,
            in2 => \_gnd_net_\,
            in3 => \N__40656\,
            lcout => n12_adj_689,
            ltout => OPEN,
            carryin => n13083,
            carryout => n13084,
            clk => \N__56229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i15_LC_10_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40653\,
            in2 => \_gnd_net_\,
            in3 => \N__40647\,
            lcout => n11_adj_688,
            ltout => OPEN,
            carryin => n13084,
            carryout => n13085,
            clk => \N__56229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i16_LC_10_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40830\,
            in2 => \_gnd_net_\,
            in3 => \N__40824\,
            lcout => n10_adj_687,
            ltout => OPEN,
            carryin => \bfn_10_31_0_\,
            carryout => n13086,
            clk => \N__56236\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i17_LC_10_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40821\,
            in2 => \_gnd_net_\,
            in3 => \N__40815\,
            lcout => n9_adj_686,
            ltout => OPEN,
            carryin => n13086,
            carryout => n13087,
            clk => \N__56236\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i18_LC_10_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40812\,
            in2 => \_gnd_net_\,
            in3 => \N__40806\,
            lcout => n8_adj_685,
            ltout => OPEN,
            carryin => n13087,
            carryout => n13088,
            clk => \N__56236\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i19_LC_10_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40803\,
            in2 => \_gnd_net_\,
            in3 => \N__40797\,
            lcout => n7_adj_684,
            ltout => OPEN,
            carryin => n13088,
            carryout => n13089,
            clk => \N__56236\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i20_LC_10_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40794\,
            in2 => \_gnd_net_\,
            in3 => \N__40788\,
            lcout => n6_adj_683,
            ltout => OPEN,
            carryin => n13089,
            carryout => n13090,
            clk => \N__56236\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i21_LC_10_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40780\,
            in2 => \_gnd_net_\,
            in3 => \N__40767\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n13090,
            carryout => n13091,
            clk => \N__56236\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i22_LC_10_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40762\,
            in2 => \_gnd_net_\,
            in3 => \N__40749\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n13091,
            carryout => n13092,
            clk => \N__56236\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i23_LC_10_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40741\,
            in2 => \_gnd_net_\,
            in3 => \N__40728\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n13092,
            carryout => n13093,
            clk => \N__56236\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i24_LC_10_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40990\,
            in2 => \_gnd_net_\,
            in3 => \N__40977\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_10_32_0_\,
            carryout => n13094,
            clk => \N__56242\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_663__i25_LC_10_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40970\,
            in2 => \_gnd_net_\,
            in3 => \N__40974\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56242\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1185_3_lut_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43692\,
            in1 => \N__43347\,
            in2 => \_gnd_net_\,
            in3 => \N__45476\,
            lcout => n1833,
            ltout => \n1833_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10012_4_lut_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__40949\,
            in1 => \N__40847\,
            in2 => \N__40959\,
            in3 => \N__40879\,
            lcout => n11989,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1184_3_lut_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43332\,
            in2 => \N__45499\,
            in3 => \N__45537\,
            lcout => n1832,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_2_lut_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40948\,
            in2 => \_gnd_net_\,
            in3 => \N__40914\,
            lcout => n1901,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => n12606,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_3_lut_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55285\,
            in2 => \N__40910\,
            in3 => \N__40887\,
            lcout => n1900,
            ltout => OPEN,
            carryin => n12606,
            carryout => n12607,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_4_lut_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40884\,
            in3 => \N__40854\,
            lcout => n1899,
            ltout => OPEN,
            carryin => n12607,
            carryout => n12608,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_5_lut_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55286\,
            in2 => \N__40851\,
            in3 => \N__41058\,
            lcout => n1898,
            ltout => OPEN,
            carryin => n12608,
            carryout => n12609,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_6_lut_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43111\,
            in3 => \N__41049\,
            lcout => n1897,
            ltout => OPEN,
            carryin => n12609,
            carryout => n12610,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_7_lut_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41667\,
            in3 => \N__41040\,
            lcout => n1896,
            ltout => OPEN,
            carryin => n12610,
            carryout => n12611,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_8_lut_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55087\,
            in2 => \N__42848\,
            in3 => \N__41037\,
            lcout => n1895,
            ltout => OPEN,
            carryin => n12611,
            carryout => n12612,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_9_lut_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55287\,
            in2 => \N__43169\,
            in3 => \N__41034\,
            lcout => n1894,
            ltout => OPEN,
            carryin => n12612,
            carryout => n12613,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_10_lut_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55281\,
            in2 => \N__43082\,
            in3 => \N__41025\,
            lcout => n1893,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => n12614,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_11_lut_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54955\,
            in2 => \N__42878\,
            in3 => \N__41022\,
            lcout => n1892,
            ltout => OPEN,
            carryin => n12614,
            carryout => n12615,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_12_lut_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55282\,
            in2 => \N__43058\,
            in3 => \N__41010\,
            lcout => n1891,
            ltout => OPEN,
            carryin => n12615,
            carryout => n12616,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_13_lut_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54956\,
            in2 => \N__43031\,
            in3 => \N__40995\,
            lcout => n1890,
            ltout => OPEN,
            carryin => n12616,
            carryout => n12617,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_14_lut_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55283\,
            in2 => \N__41087\,
            in3 => \N__41181\,
            lcout => n1889,
            ltout => OPEN,
            carryin => n12617,
            carryout => n12618,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_15_lut_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54957\,
            in2 => \N__43142\,
            in3 => \N__41178\,
            lcout => n1888,
            ltout => OPEN,
            carryin => n12618,
            carryout => n12619,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_16_lut_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55284\,
            in2 => \N__43193\,
            in3 => \N__41163\,
            lcout => n1887,
            ltout => OPEN,
            carryin => n12619,
            carryout => n12620,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_17_lut_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54958\,
            in2 => \N__41228\,
            in3 => \N__41148\,
            lcout => n1886,
            ltout => OPEN,
            carryin => n12620,
            carryout => n12621,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1235_18_lut_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__55280\,
            in1 => \_gnd_net_\,
            in2 => \N__43749\,
            in3 => \N__41145\,
            lcout => n1885,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1244_3_lut_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42879\,
            in2 => \N__41142\,
            in3 => \N__41503\,
            lcout => n1924,
            ltout => \n1924_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_140_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41725\,
            in2 => \N__41106\,
            in3 => \N__41683\,
            lcout => n14438,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1174_3_lut_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__43467\,
            in1 => \_gnd_net_\,
            in2 => \N__45506\,
            in3 => \N__43487\,
            lcout => n1822,
            ltout => \n1822_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_139_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43186\,
            in2 => \N__41070\,
            in3 => \N__43135\,
            lcout => n14534,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1247_3_lut_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42849\,
            in2 => \N__41757\,
            in3 => \N__41502\,
            lcout => n1927,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1246_3_lut_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41712\,
            in2 => \N__43170\,
            in3 => \N__41501\,
            lcout => n1926,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1181_3_lut_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43242\,
            in2 => \N__45501\,
            in3 => \N__45702\,
            lcout => n1829,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1237_3_lut_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43735\,
            in2 => \N__41646\,
            in3 => \N__41505\,
            lcout => n1917,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i4_3_lut_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__41613\,
            in1 => \_gnd_net_\,
            in2 => \N__41601\,
            in3 => \N__49539\,
            lcout => n316,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1240_3_lut_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41532\,
            in2 => \N__43143\,
            in3 => \N__41504\,
            lcout => n1920,
            ltout => \n1920_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1307_3_lut_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41397\,
            in2 => \N__41385\,
            in3 => \N__41378\,
            lcout => n2019,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1171_3_lut_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43368\,
            in2 => \N__43395\,
            in3 => \N__45502\,
            lcout => n1819,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i18_3_lut_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__41918\,
            in1 => \_gnd_net_\,
            in2 => \N__49553\,
            in3 => \N__41967\,
            lcout => n302,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i30_3_lut_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41950\,
            in2 => \N__49552\,
            in3 => \N__42316\,
            lcout => n404,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41917\,
            lcout => n16_adj_634,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41817\,
            lcout => n7_adj_625,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42003\,
            lcout => n3_adj_621,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10989_3_lut_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41859\,
            in2 => \N__41853\,
            in3 => \N__42188\,
            lcout => OPEN,
            ltout => \n13662_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12421_3_lut_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49493\,
            in2 => \N__41832\,
            in3 => \N__41821\,
            lcout => n833,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10987_3_lut_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42348\,
            in2 => \N__41796\,
            in3 => \N__42189\,
            lcout => OPEN,
            ltout => \n13660_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10988_3_lut_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__41784\,
            in1 => \_gnd_net_\,
            in2 => \N__41760\,
            in3 => \N__49494\,
            lcout => n832,
            ltout => \n832_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10050_4_lut_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__43585\,
            in1 => \N__43875\,
            in2 => \N__42087\,
            in3 => \N__42151\,
            lcout => n12027,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10985_3_lut_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42264\,
            in2 => \N__42195\,
            in3 => \N__42084\,
            lcout => OPEN,
            ltout => \n13658_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10986_3_lut_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__49495\,
            in1 => \_gnd_net_\,
            in2 => \N__42078\,
            in3 => \N__42063\,
            lcout => n831,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i5_1_lut_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__42036\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n21_adj_555,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i569_3_lut_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44089\,
            in2 => \N__42125\,
            in3 => \N__42099\,
            lcout => n929,
            ltout => \n929_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_85_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42024\,
            in3 => \N__46096\,
            lcout => n14460,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10982_3_lut_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__49600\,
            in1 => \_gnd_net_\,
            in2 => \N__42021\,
            in3 => \N__41985\,
            lcout => n829,
            ltout => \n829_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10150_4_lut_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__42118\,
            in1 => \N__42377\,
            in2 => \N__41979\,
            in3 => \N__41976\,
            lcout => n861,
            ltout => \n861_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i570_3_lut_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42155\,
            in2 => \N__41970\,
            in3 => \N__42135\,
            lcout => n930,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_83_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__42347\,
            in1 => \N__42317\,
            in2 => \N__42281\,
            in3 => \N__42263\,
            lcout => n5_adj_682,
            ltout => \n5_adj_682_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_84_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42219\,
            in2 => \N__42198\,
            in3 => \N__42427\,
            lcout => n13653,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_2_lut_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43874\,
            in2 => \_gnd_net_\,
            in3 => \N__42168\,
            lcout => n901,
            ltout => OPEN,
            carryin => \bfn_11_24_0_\,
            carryout => n12501,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_3_lut_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53813\,
            in2 => \N__43592\,
            in3 => \N__42165\,
            lcout => n900,
            ltout => OPEN,
            carryin => n12501,
            carryout => n12502,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_4_lut_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43620\,
            in3 => \N__42162\,
            lcout => n899,
            ltout => OPEN,
            carryin => n12502,
            carryout => n12503,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_5_lut_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53814\,
            in2 => \N__42159\,
            in3 => \N__42129\,
            lcout => n898,
            ltout => OPEN,
            carryin => n12503,
            carryout => n12504,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_6_lut_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42126\,
            in3 => \N__42093\,
            lcout => n897,
            ltout => OPEN,
            carryin => n12504,
            carryout => n12505,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_7_lut_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__44063\,
            in3 => \N__42090\,
            lcout => n896,
            ltout => OPEN,
            carryin => n12505,
            carryout => n12506,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_565_8_lut_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__53815\,
            in1 => \N__44093\,
            in2 => \N__42381\,
            in3 => \N__42432\,
            lcout => n927,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i500_4_lut_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__42429\,
            in1 => \N__49560\,
            in2 => \N__42399\,
            in3 => \N__42390\,
            lcout => n828,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i4_1_lut_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42366\,
            lcout => n22_adj_554,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i7_1_lut_LC_11_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__42357\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n19_adj_557,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i4_1_lut_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46142\,
            lcout => n22_adj_594,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i8_1_lut_LC_11_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44333\,
            lcout => n18_adj_590,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i1_1_lut_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44501\,
            lcout => n25_adj_597,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i6_1_lut_LC_11_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43958\,
            lcout => n20_adj_592,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i5_1_lut_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43991\,
            lcout => n21_adj_593,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i3_1_lut_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42513\,
            lcout => n23_adj_553,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_2_lut_LC_11_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42504\,
            in2 => \_gnd_net_\,
            in3 => \N__42498\,
            lcout => \pwm_setpoint_23_N_171_0\,
            ltout => OPEN,
            carryin => \bfn_11_26_0_\,
            carryout => n12426,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_3_lut_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47850\,
            in2 => \_gnd_net_\,
            in3 => \N__42495\,
            lcout => \pwm_setpoint_23_N_171_1\,
            ltout => OPEN,
            carryin => n12426,
            carryout => n12427,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_4_lut_LC_11_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46512\,
            in2 => \_gnd_net_\,
            in3 => \N__42492\,
            lcout => \pwm_setpoint_23_N_171_2\,
            ltout => OPEN,
            carryin => n12427,
            carryout => n12428,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_5_lut_LC_11_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42489\,
            in2 => \_gnd_net_\,
            in3 => \N__42483\,
            lcout => \pwm_setpoint_23_N_171_3\,
            ltout => OPEN,
            carryin => n12428,
            carryout => n12429,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_6_lut_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42480\,
            in2 => \_gnd_net_\,
            in3 => \N__42468\,
            lcout => \pwm_setpoint_23_N_171_4\,
            ltout => OPEN,
            carryin => n12429,
            carryout => n12430,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_7_lut_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42465\,
            in2 => \_gnd_net_\,
            in3 => \N__42453\,
            lcout => \pwm_setpoint_23_N_171_5\,
            ltout => OPEN,
            carryin => n12430,
            carryout => n12431,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_8_lut_LC_11_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47301\,
            in2 => \_gnd_net_\,
            in3 => \N__42450\,
            lcout => \pwm_setpoint_23_N_171_6\,
            ltout => OPEN,
            carryin => n12431,
            carryout => n12432,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_9_lut_LC_11_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42447\,
            in2 => \_gnd_net_\,
            in3 => \N__42435\,
            lcout => \pwm_setpoint_23_N_171_7\,
            ltout => OPEN,
            carryin => n12432,
            carryout => n12433,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_10_lut_LC_11_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42639\,
            in2 => \_gnd_net_\,
            in3 => \N__42621\,
            lcout => \pwm_setpoint_23_N_171_8\,
            ltout => OPEN,
            carryin => \bfn_11_27_0_\,
            carryout => n12434,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_11_lut_LC_11_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42618\,
            in2 => \_gnd_net_\,
            in3 => \N__42606\,
            lcout => \pwm_setpoint_23_N_171_9\,
            ltout => OPEN,
            carryin => n12434,
            carryout => n12435,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_12_lut_LC_11_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42603\,
            in2 => \_gnd_net_\,
            in3 => \N__42591\,
            lcout => \pwm_setpoint_23_N_171_10\,
            ltout => OPEN,
            carryin => n12435,
            carryout => n12436,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_13_lut_LC_11_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42588\,
            in2 => \_gnd_net_\,
            in3 => \N__42570\,
            lcout => \pwm_setpoint_23_N_171_11\,
            ltout => OPEN,
            carryin => n12436,
            carryout => n12437,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_14_lut_LC_11_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44937\,
            in2 => \_gnd_net_\,
            in3 => \N__42567\,
            lcout => \pwm_setpoint_23_N_171_12\,
            ltout => OPEN,
            carryin => n12437,
            carryout => n12438,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_15_lut_LC_11_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42564\,
            in2 => \_gnd_net_\,
            in3 => \N__42552\,
            lcout => \pwm_setpoint_23_N_171_13\,
            ltout => OPEN,
            carryin => n12438,
            carryout => n12439,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_16_lut_LC_11_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42549\,
            in2 => \_gnd_net_\,
            in3 => \N__42537\,
            lcout => \pwm_setpoint_23_N_171_14\,
            ltout => OPEN,
            carryin => n12439,
            carryout => n12440,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_17_lut_LC_11_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42534\,
            in2 => \_gnd_net_\,
            in3 => \N__42516\,
            lcout => \pwm_setpoint_23_N_171_15\,
            ltout => OPEN,
            carryin => n12440,
            carryout => n12441,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_18_lut_LC_11_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42684\,
            in2 => \_gnd_net_\,
            in3 => \N__42675\,
            lcout => \pwm_setpoint_23_N_171_16\,
            ltout => OPEN,
            carryin => \bfn_11_28_0_\,
            carryout => n12442,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_19_lut_LC_11_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44580\,
            in2 => \_gnd_net_\,
            in3 => \N__42672\,
            lcout => \pwm_setpoint_23_N_171_17\,
            ltout => OPEN,
            carryin => n12442,
            carryout => n12443,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_20_lut_LC_11_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44532\,
            in2 => \_gnd_net_\,
            in3 => \N__42657\,
            lcout => \pwm_setpoint_23_N_171_18\,
            ltout => OPEN,
            carryin => n12443,
            carryout => n12444,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_21_lut_LC_11_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46737\,
            in2 => \_gnd_net_\,
            in3 => \N__42654\,
            lcout => \pwm_setpoint_23_N_171_19\,
            ltout => OPEN,
            carryin => n12444,
            carryout => n12445,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_22_lut_LC_11_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44475\,
            in2 => \_gnd_net_\,
            in3 => \N__42651\,
            lcout => \pwm_setpoint_23_N_171_20\,
            ltout => OPEN,
            carryin => n12445,
            carryout => n12446,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_23_lut_LC_11_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44559\,
            in2 => \_gnd_net_\,
            in3 => \N__42648\,
            lcout => \pwm_setpoint_23_N_171_21\,
            ltout => OPEN,
            carryin => n12446,
            carryout => n12447,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_add_3_24_lut_LC_11_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44625\,
            in2 => \_gnd_net_\,
            in3 => \N__42645\,
            lcout => \pwm_setpoint_23_N_171_22\,
            ltout => OPEN,
            carryin => n12447,
            carryout => n12448,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i23_LC_11_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47837\,
            in2 => \_gnd_net_\,
            in3 => \N__42642\,
            lcout => pwm_setpoint_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56225\,
            ce => 'H',
            sr => \N__47838\
        );

    \LessThan_299_i19_2_lut_LC_11_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42703\,
            in2 => \_gnd_net_\,
            in3 => \N__48395\,
            lcout => n19_adj_666,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i16_3_lut_3_lut_LC_11_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__42704\,
            in1 => \N__48475\,
            in2 => \_gnd_net_\,
            in3 => \N__44878\,
            lcout => OPEN,
            ltout => \n16_adj_664_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i24_3_lut_LC_11_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44715\,
            in2 => \N__42747\,
            in3 => \N__44677\,
            lcout => OPEN,
            ltout => \n24_adj_669_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12493_4_lut_LC_11_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__44678\,
            in1 => \N__42729\,
            in2 => \N__42744\,
            in3 => \N__42741\,
            lcout => n15223,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12414_2_lut_4_lut_LC_11_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__44879\,
            in1 => \N__42705\,
            in2 => \N__48477\,
            in3 => \N__48396\,
            lcout => n15144,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i23_2_lut_LC_11_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42929\,
            in2 => \_gnd_net_\,
            in3 => \N__48344\,
            lcout => n23_adj_668,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i21_LC_11_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42723\,
            in1 => \N__50892\,
            in2 => \_gnd_net_\,
            in3 => \N__44574\,
            lcout => pwm_setpoint_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i9_LC_11_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50893\,
            in1 => \_gnd_net_\,
            in2 => \N__42717\,
            in3 => \N__44271\,
            lcout => pwm_setpoint_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12448_4_lut_LC_11_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001101"
        )
    port map (
            in0 => \N__42815\,
            in1 => \N__46809\,
            in2 => \N__46239\,
            in3 => \N__44747\,
            lcout => n15178,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i14_LC_11_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50894\,
            in1 => \N__44120\,
            in2 => \_gnd_net_\,
            in3 => \N__42693\,
            lcout => pwm_setpoint_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56237\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i22_LC_11_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__44643\,
            in1 => \N__50895\,
            in2 => \_gnd_net_\,
            in3 => \N__42825\,
            lcout => pwm_setpoint_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56237\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12380_4_lut_LC_11_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__47144\,
            in1 => \N__42780\,
            in2 => \N__42789\,
            in3 => \N__42816\,
            lcout => n15110,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i15_2_lut_LC_11_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48017\,
            in2 => \_gnd_net_\,
            in3 => \N__42965\,
            lcout => n15_adj_663,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i17_2_lut_LC_11_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42804\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47978\,
            lcout => n17_adj_665,
            ltout => \n17_adj_665_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12444_4_lut_LC_11_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111011"
        )
    port map (
            in0 => \N__42779\,
            in1 => \N__42771\,
            in2 => \N__42765\,
            in3 => \N__44733\,
            lcout => n15174,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i33_2_lut_LC_11_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__42981\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48213\,
            lcout => n33_adj_675,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12367_2_lut_4_lut_LC_11_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__48212\,
            in1 => \N__42980\,
            in2 => \N__42969\,
            in3 => \N__48018\,
            lcout => n15097,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12435_3_lut_LC_11_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__44808\,
            in1 => \N__44820\,
            in2 => \_gnd_net_\,
            in3 => \N__42906\,
            lcout => n15165,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i16_LC_11_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42762\,
            in1 => \N__50900\,
            in2 => \_gnd_net_\,
            in3 => \N__44454\,
            lcout => pwm_setpoint_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56243\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12507_4_lut_LC_11_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42753\,
            in1 => \N__44789\,
            in2 => \N__47145\,
            in3 => \N__44807\,
            lcout => n15237,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i17_LC_11_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50901\,
            in1 => \N__44598\,
            in2 => \_gnd_net_\,
            in3 => \N__42990\,
            lcout => pwm_setpoint_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56243\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i12_3_lut_3_lut_LC_11_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__48211\,
            in1 => \N__42979\,
            in2 => \_gnd_net_\,
            in3 => \N__42964\,
            lcout => n12_adj_661,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i10_LC_11_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50910\,
            in1 => \N__42939\,
            in2 => \_gnd_net_\,
            in3 => \N__44235\,
            lcout => pwm_setpoint_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56249\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12474_3_lut_LC_11_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47094\,
            in1 => \N__42930\,
            in2 => \_gnd_net_\,
            in3 => \N__44790\,
            lcout => n15204,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i35_2_lut_LC_11_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42896\,
            in2 => \_gnd_net_\,
            in3 => \N__48582\,
            lcout => n35,
            ltout => \n35_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i30_3_lut_LC_11_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__42897\,
            in1 => \_gnd_net_\,
            in2 => \N__42888\,
            in3 => \N__42885\,
            lcout => n30_adj_673,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1177_3_lut_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43553\,
            in2 => \N__43539\,
            in3 => \N__45457\,
            lcout => n1825,
            ltout => \n1825_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_136_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43075\,
            in1 => \N__42841\,
            in2 => \N__42861\,
            in3 => \N__43162\,
            lcout => n14520,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1180_3_lut_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43233\,
            in2 => \N__45681\,
            in3 => \N__45456\,
            lcout => n1828,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1182_3_lut_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__43272\,
            in1 => \_gnd_net_\,
            in2 => \N__45486\,
            in3 => \N__43254\,
            lcout => n1830,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12904_4_lut_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43418\,
            in1 => \N__43390\,
            in2 => \N__45341\,
            in3 => \N__42996\,
            lcout => n1752,
            ltout => \n1752_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12480_3_lut_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45314\,
            in2 => \N__43086\,
            in3 => \N__43206\,
            lcout => n1826,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1176_3_lut_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43521\,
            in2 => \N__45210\,
            in3 => \N__45461\,
            lcout => n1824,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1175_3_lut_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45245\,
            in2 => \N__45485\,
            in3 => \N__43506\,
            lcout => n1823,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12478_3_lut_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45135\,
            in2 => \N__47211\,
            in3 => \N__45608\,
            lcout => n1726,
            ltout => \n1726_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_132_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__45277\,
            in1 => \_gnd_net_\,
            in2 => \N__43005\,
            in3 => \N__45310\,
            lcout => OPEN,
            ltout => \n14244_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_133_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45235\,
            in1 => \N__45196\,
            in2 => \N__43002\,
            in3 => \N__43483\,
            lcout => OPEN,
            ltout => \n14250_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_135_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__43448\,
            in1 => \N__43353\,
            in2 => \N__42999\,
            in3 => \N__45654\,
            lcout => n14254,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1105_3_lut_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47181\,
            in2 => \N__45099\,
            in3 => \N__45609\,
            lcout => n1721,
            ltout => \n1721_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1172_3_lut_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__45455\,
            in1 => \_gnd_net_\,
            in2 => \N__43197\,
            in3 => \N__43407\,
            lcout => n1820,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1179_3_lut_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45278\,
            in2 => \N__43221\,
            in3 => \N__45454\,
            lcout => n1827,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1104_3_lut_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__45087\,
            in1 => \_gnd_net_\,
            in2 => \N__45372\,
            in3 => \N__45604\,
            lcout => n1720,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1107_3_lut_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__45602\,
            in1 => \_gnd_net_\,
            in2 => \N__47283\,
            in3 => \N__45120\,
            lcout => n1723,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1106_3_lut_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45603\,
            in2 => \N__45111\,
            in3 => \N__47253\,
            lcout => n1722,
            ltout => \n1722_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1173_3_lut_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__45484\,
            in1 => \_gnd_net_\,
            in2 => \N__43146\,
            in3 => \N__43437\,
            lcout => n1821,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1116_3_lut_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44985\,
            in2 => \N__48756\,
            in3 => \N__45598\,
            lcout => n1732,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1115_3_lut_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__44973\,
            in1 => \_gnd_net_\,
            in2 => \N__45616\,
            in3 => \N__48810\,
            lcout => n1731,
            ltout => \n1731_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10014_4_lut_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__43687\,
            in1 => \N__43303\,
            in2 => \N__43356\,
            in3 => \N__45526\,
            lcout => n11991,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_2_lut_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43688\,
            in2 => \_gnd_net_\,
            in3 => \N__43335\,
            lcout => n1801,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => n12591,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_3_lut_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54881\,
            in2 => \N__45533\,
            in3 => \N__43320\,
            lcout => n1800,
            ltout => OPEN,
            carryin => n12591,
            carryout => n12592,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_4_lut_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43310\,
            in3 => \N__43275\,
            lcout => n1799,
            ltout => OPEN,
            carryin => n12592,
            carryout => n12593,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_5_lut_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54882\,
            in2 => \N__43271\,
            in3 => \N__43245\,
            lcout => n1798,
            ltout => OPEN,
            carryin => n12593,
            carryout => n12594,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_6_lut_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45701\,
            in3 => \N__43236\,
            lcout => n1797,
            ltout => OPEN,
            carryin => n12594,
            carryout => n12595,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_7_lut_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45677\,
            in3 => \N__43224\,
            lcout => n1796,
            ltout => OPEN,
            carryin => n12595,
            carryout => n12596,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_8_lut_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55086\,
            in2 => \N__45282\,
            in3 => \N__43209\,
            lcout => n1795,
            ltout => OPEN,
            carryin => n12596,
            carryout => n12597,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_9_lut_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54883\,
            in2 => \N__45318\,
            in3 => \N__43563\,
            lcout => n1794,
            ltout => OPEN,
            carryin => n12597,
            carryout => n12598,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_10_lut_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54586\,
            in2 => \N__43560\,
            in3 => \N__43524\,
            lcout => n1793,
            ltout => OPEN,
            carryin => \bfn_12_21_0_\,
            carryout => n12599,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_11_lut_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54590\,
            in2 => \N__45209\,
            in3 => \N__43509\,
            lcout => n1792,
            ltout => OPEN,
            carryin => n12599,
            carryout => n12600,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_12_lut_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54587\,
            in2 => \N__45246\,
            in3 => \N__43494\,
            lcout => n1791,
            ltout => OPEN,
            carryin => n12600,
            carryout => n12601,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_13_lut_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54591\,
            in2 => \N__43491\,
            in3 => \N__43458\,
            lcout => n1790,
            ltout => OPEN,
            carryin => n12601,
            carryout => n12602,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_14_lut_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54588\,
            in2 => \N__43455\,
            in3 => \N__43428\,
            lcout => n1789,
            ltout => OPEN,
            carryin => n12602,
            carryout => n12603,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_15_lut_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54592\,
            in2 => \N__43425\,
            in3 => \N__43398\,
            lcout => n1788,
            ltout => OPEN,
            carryin => n12603,
            carryout => n12604,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_16_lut_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43391\,
            in2 => \N__54880\,
            in3 => \N__43362\,
            lcout => n1787,
            ltout => OPEN,
            carryin => n12604,
            carryout => n12605,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1168_17_lut_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__54589\,
            in1 => \N__45345\,
            in2 => \N__45389\,
            in3 => \N__43359\,
            lcout => n1818,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43838\,
            lcout => n10_adj_628,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i17_3_lut_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49611\,
            in1 => \N__43704\,
            in2 => \_gnd_net_\,
            in3 => \N__45759\,
            lcout => n303,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i19_3_lut_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43668\,
            in1 => \N__49610\,
            in2 => \_gnd_net_\,
            in3 => \N__43655\,
            lcout => n301,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i571_3_lut_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43626\,
            in2 => \N__43619\,
            in3 => \N__44090\,
            lcout => n931,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i636_3_lut_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46064\,
            in2 => \N__46013\,
            in3 => \N__46050\,
            lcout => n1028,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i572_3_lut_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43599\,
            in2 => \N__43593\,
            in3 => \N__44092\,
            lcout => n932,
            ltout => \n932_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i639_3_lut_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__46004\,
            in1 => \_gnd_net_\,
            in2 => \N__43566\,
            in3 => \N__45864\,
            lcout => n1031,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i641_3_lut_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45924\,
            in1 => \N__45912\,
            in2 => \_gnd_net_\,
            in3 => \N__46002\,
            lcout => n1033,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i26_3_lut_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49599\,
            in2 => \N__43920\,
            in3 => \N__43887\,
            lcout => n41,
            ltout => \n41_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i573_3_lut_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__43863\,
            in1 => \_gnd_net_\,
            in2 => \N__43857\,
            in3 => \N__44091\,
            lcout => n933,
            ltout => \n933_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i640_3_lut_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__46003\,
            in1 => \_gnd_net_\,
            in2 => \N__43854\,
            in3 => \N__45888\,
            lcout => n1032,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i635_rep_47_3_lut_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46037\,
            in2 => \N__46014\,
            in3 => \N__46023\,
            lcout => n1027,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i24_3_lut_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49602\,
            in2 => \N__43851\,
            in3 => \N__43839\,
            lcout => n296,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i25_3_lut_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__43808\,
            in1 => \N__49601\,
            in2 => \_gnd_net_\,
            in3 => \N__43779\,
            lcout => n295,
            ltout => \n295_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9978_4_lut_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__45850\,
            in1 => \N__45899\,
            in2 => \N__43764\,
            in3 => \N__45875\,
            lcout => OPEN,
            ltout => \n11955_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_86_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__46036\,
            in1 => \N__45968\,
            in2 => \N__43761\,
            in3 => \N__43758\,
            lcout => n960,
            ltout => \n960_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i637_3_lut_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__46100\,
            in1 => \_gnd_net_\,
            in2 => \N__43752\,
            in3 => \N__46080\,
            lcout => n1029,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i568_3_lut_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44094\,
            in2 => \N__44064\,
            in3 => \N__44046\,
            lcout => n928,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i0_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45945\,
            in2 => \N__49770\,
            in3 => \N__44040\,
            lcout => duty_0,
            ltout => OPEN,
            carryin => \bfn_12_25_0_\,
            carryout => n12473,
            clk => \N__56218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i1_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44037\,
            in2 => \N__49740\,
            in3 => \N__44028\,
            lcout => duty_1,
            ltout => OPEN,
            carryin => n12473,
            carryout => n12474,
            clk => \N__56218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i2_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44025\,
            in2 => \N__49704\,
            in3 => \N__44019\,
            lcout => duty_2,
            ltout => OPEN,
            carryin => n12474,
            carryout => n12475,
            clk => \N__56218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i3_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44016\,
            in2 => \N__50352\,
            in3 => \N__44010\,
            lcout => duty_3,
            ltout => OPEN,
            carryin => n12475,
            carryout => n12476,
            clk => \N__56218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i4_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44007\,
            in2 => \N__50319\,
            in3 => \N__43980\,
            lcout => duty_4,
            ltout => OPEN,
            carryin => n12476,
            carryout => n12477,
            clk => \N__56218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i5_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43977\,
            in2 => \N__50274\,
            in3 => \N__43947\,
            lcout => duty_5,
            ltout => OPEN,
            carryin => n12477,
            carryout => n12478,
            clk => \N__56218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i6_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43944\,
            in2 => \N__50238\,
            in3 => \N__43938\,
            lcout => duty_6,
            ltout => OPEN,
            carryin => n12478,
            carryout => n12479,
            clk => \N__56218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i7_LC_12_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43935\,
            in2 => \N__50202\,
            in3 => \N__44322\,
            lcout => duty_7,
            ltout => OPEN,
            carryin => n12479,
            carryout => n12480,
            clk => \N__56218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i8_LC_12_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44319\,
            in2 => \N__50157\,
            in3 => \N__44283\,
            lcout => duty_8,
            ltout => OPEN,
            carryin => \bfn_12_26_0_\,
            carryout => n12481,
            clk => \N__56221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i9_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44280\,
            in2 => \N__50118\,
            in3 => \N__44247\,
            lcout => duty_9,
            ltout => OPEN,
            carryin => n12481,
            carryout => n12482,
            clk => \N__56221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i10_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44244\,
            in2 => \N__50076\,
            in3 => \N__44214\,
            lcout => duty_10,
            ltout => OPEN,
            carryin => n12482,
            carryout => n12483,
            clk => \N__56221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i11_LC_12_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44211\,
            in2 => \N__50709\,
            in3 => \N__44178\,
            lcout => duty_11,
            ltout => OPEN,
            carryin => n12483,
            carryout => n12484,
            clk => \N__56221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i12_LC_12_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50674\,
            in2 => \N__44175\,
            in3 => \N__44163\,
            lcout => duty_12,
            ltout => OPEN,
            carryin => n12484,
            carryout => n12485,
            clk => \N__56221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i13_LC_12_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44160\,
            in2 => \N__50637\,
            in3 => \N__44133\,
            lcout => duty_13,
            ltout => OPEN,
            carryin => n12485,
            carryout => n12486,
            clk => \N__56221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i14_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44130\,
            in2 => \N__50598\,
            in3 => \N__44097\,
            lcout => duty_14,
            ltout => OPEN,
            carryin => n12486,
            carryout => n12487,
            clk => \N__56221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i15_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44469\,
            in2 => \N__50565\,
            in3 => \N__44457\,
            lcout => duty_15,
            ltout => OPEN,
            carryin => n12487,
            carryout => n12488,
            clk => \N__56221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i16_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47883\,
            in2 => \N__50517\,
            in3 => \N__44433\,
            lcout => duty_16,
            ltout => OPEN,
            carryin => \bfn_12_27_0_\,
            carryout => n12489,
            clk => \N__56226\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i17_LC_12_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44430\,
            in2 => \N__50481\,
            in3 => \N__44418\,
            lcout => duty_17,
            ltout => OPEN,
            carryin => n12489,
            carryout => n12490,
            clk => \N__56226\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i18_LC_12_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44415\,
            in2 => \N__50436\,
            in3 => \N__44406\,
            lcout => duty_18,
            ltout => OPEN,
            carryin => n12490,
            carryout => n12491,
            clk => \N__56226\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i19_LC_12_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44403\,
            in2 => \N__50396\,
            in3 => \N__44394\,
            lcout => duty_19,
            ltout => OPEN,
            carryin => n12491,
            carryout => n12492,
            clk => \N__56226\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i20_LC_12_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44391\,
            in2 => \N__51300\,
            in3 => \N__44379\,
            lcout => duty_20,
            ltout => OPEN,
            carryin => n12492,
            carryout => n12493,
            clk => \N__56226\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i21_LC_12_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44376\,
            in2 => \N__51270\,
            in3 => \N__44367\,
            lcout => duty_21,
            ltout => OPEN,
            carryin => n12493,
            carryout => n12494,
            clk => \N__56226\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i22_LC_12_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44364\,
            in2 => \N__51228\,
            in3 => \N__44355\,
            lcout => duty_22,
            ltout => OPEN,
            carryin => n12494,
            carryout => n12495,
            clk => \N__56226\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \duty_i23_LC_12_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__51054\,
            in1 => \N__44352\,
            in2 => \_gnd_net_\,
            in3 => \N__44343\,
            lcout => duty_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56226\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i18_1_lut_LC_12_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44591\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n8_adj_580,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i22_1_lut_LC_12_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44570\,
            lcout => n4_adj_576,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i19_1_lut_LC_12_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44543\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n7_adj_579,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i19_LC_12_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__50833\,
            in1 => \_gnd_net_\,
            in2 => \N__46752\,
            in3 => \N__44526\,
            lcout => pwm_setpoint_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i20_LC_12_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__44484\,
            in1 => \N__50834\,
            in2 => \_gnd_net_\,
            in3 => \N__44520\,
            lcout => pwm_setpoint_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i4_4_lut_LC_12_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__48156\,
            in1 => \N__47940\,
            in2 => \N__48177\,
            in3 => \N__44490\,
            lcout => n4_adj_655,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i0_LC_12_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44514\,
            in1 => \N__50832\,
            in2 => \_gnd_net_\,
            in3 => \N__44505\,
            lcout => pwm_setpoint_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i21_1_lut_LC_12_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44483\,
            lcout => n5_adj_577,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i45_2_lut_LC_12_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44711\,
            in2 => \_gnd_net_\,
            in3 => \N__48432\,
            lcout => n45,
            ltout => \n45_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12515_4_lut_LC_12_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__44649\,
            in1 => \N__44838\,
            in2 => \N__44700\,
            in3 => \N__44685\,
            lcout => n15245,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i41_2_lut_LC_12_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44696\,
            in2 => \_gnd_net_\,
            in3 => \N__48504\,
            lcout => n41_adj_678,
            ltout => \n41_adj_678_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12522_3_lut_LC_12_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__44697\,
            in1 => \_gnd_net_\,
            in2 => \N__44688\,
            in3 => \N__44604\,
            lcout => n40_adj_677,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12513_4_lut_LC_12_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__44679\,
            in1 => \N__44664\,
            in2 => \N__44757\,
            in3 => \N__44658\,
            lcout => n15243,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i23_1_lut_LC_12_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44639\,
            lcout => n3_adj_575,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i13_2_lut_LC_12_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__46208\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48056\,
            lcout => n13_adj_662,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i39_2_lut_LC_12_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44618\,
            in2 => \_gnd_net_\,
            in3 => \N__48528\,
            lcout => n39_adj_676,
            ltout => \n39_adj_676_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12524_3_lut_LC_12_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__44619\,
            in1 => \_gnd_net_\,
            in2 => \N__44607\,
            in3 => \N__44997\,
            lcout => n15254,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i43_2_lut_LC_12_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48476\,
            in2 => \_gnd_net_\,
            in3 => \N__44880\,
            lcout => n43,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i12_LC_12_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50873\,
            in1 => \N__44955\,
            in2 => \_gnd_net_\,
            in3 => \N__44865\,
            lcout => pwm_setpoint_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12361_4_lut_LC_12_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__44766\,
            in1 => \N__44856\,
            in2 => \N__44850\,
            in3 => \N__44907\,
            lcout => n15091,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12499_3_lut_LC_12_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__46575\,
            in1 => \N__46540\,
            in2 => \_gnd_net_\,
            in3 => \N__44829\,
            lcout => n15229,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i25_2_lut_LC_12_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44819\,
            in2 => \_gnd_net_\,
            in3 => \N__48318\,
            lcout => n25_adj_670,
            ltout => \n25_adj_670_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12416_4_lut_LC_12_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__44799\,
            in1 => \N__44788\,
            in2 => \N__44769\,
            in3 => \N__44765\,
            lcout => n15146,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \commutation_state_i1_LC_12_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001100100010"
        )
    port map (
            in0 => \N__47005\,
            in1 => \N__46957\,
            in2 => \N__46905\,
            in3 => \N__56319\,
            lcout => commutation_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56250\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12374_4_lut_LC_12_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__46547\,
            in1 => \N__44748\,
            in2 => \N__46805\,
            in3 => \N__44732\,
            lcout => n15104,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12500_3_lut_LC_12_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__46784\,
            in1 => \N__46765\,
            in2 => \_gnd_net_\,
            in3 => \N__44721\,
            lcout => n15230,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i10_3_lut_3_lut_LC_12_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__46830\,
            in1 => \N__46212\,
            in2 => \_gnd_net_\,
            in3 => \N__48057\,
            lcout => n10_adj_659,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i13_1_lut_LC_12_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44954\,
            lcout => n13_adj_585,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_LC_12_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__46956\,
            in1 => \N__47004\,
            in2 => \_gnd_net_\,
            in3 => \N__46899\,
            lcout => \commutation_state_7__N_261\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i31_2_lut_LC_12_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46475\,
            in2 => \_gnd_net_\,
            in3 => \N__48242\,
            lcout => n31_adj_674,
            ltout => \n31_adj_674_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12490_3_lut_LC_12_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__46476\,
            in1 => \_gnd_net_\,
            in2 => \N__44925\,
            in3 => \N__44922\,
            lcout => n15220,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12465_4_lut_LC_12_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__45060\,
            in1 => \N__44916\,
            in2 => \N__46770\,
            in3 => \N__46548\,
            lcout => OPEN,
            ltout => \n15195_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12511_4_lut_LC_12_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45078\,
            in1 => \N__45006\,
            in2 => \N__44910\,
            in3 => \N__45050\,
            lcout => n15241,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i37_2_lut_LC_12_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45020\,
            in2 => \_gnd_net_\,
            in3 => \N__48555\,
            lcout => n37,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12517_4_lut_LC_12_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__44898\,
            in1 => \N__44892\,
            in2 => \N__45051\,
            in3 => \N__44886\,
            lcout => n15247,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12369_4_lut_LC_12_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__45077\,
            in1 => \N__46766\,
            in2 => \N__45069\,
            in3 => \N__45059\,
            lcout => OPEN,
            ltout => \n15099_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12527_4_lut_LC_12_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__45049\,
            in1 => \N__45036\,
            in2 => \N__45030\,
            in3 => \N__45027\,
            lcout => OPEN,
            ltout => \n15257_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12528_3_lut_LC_12_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45021\,
            in2 => \N__45009\,
            in3 => \N__45005\,
            lcout => n15258,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_2_lut_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48788\,
            in2 => \_gnd_net_\,
            in3 => \N__44988\,
            lcout => n1701,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => n12577,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_3_lut_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53850\,
            in2 => \N__48749\,
            in3 => \N__44976\,
            lcout => n1700,
            ltout => OPEN,
            carryin => n12577,
            carryout => n12578,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_4_lut_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__48809\,
            in3 => \N__44964\,
            lcout => n1699,
            ltout => OPEN,
            carryin => n12578,
            carryout => n12579,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_5_lut_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53851\,
            in2 => \N__48926\,
            in3 => \N__44961\,
            lcout => n1698,
            ltout => OPEN,
            carryin => n12579,
            carryout => n12580,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_6_lut_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__47081\,
            in3 => \N__44958\,
            lcout => n1697,
            ltout => OPEN,
            carryin => n12580,
            carryout => n12581,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_7_lut_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__47063\,
            in3 => \N__45141\,
            lcout => n1696,
            ltout => OPEN,
            carryin => n12581,
            carryout => n12582,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_8_lut_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47406\,
            in2 => \N__54246\,
            in3 => \N__45138\,
            lcout => n1695,
            ltout => OPEN,
            carryin => n12582,
            carryout => n12583,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_9_lut_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53855\,
            in2 => \N__47207\,
            in3 => \N__45129\,
            lcout => n1694,
            ltout => OPEN,
            carryin => n12583,
            carryout => n12584,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_10_lut_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53841\,
            in2 => \N__47340\,
            in3 => \N__45126\,
            lcout => n1693_adj_614,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => n12585,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_11_lut_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54953\,
            in2 => \N__45156\,
            in3 => \N__45123\,
            lcout => n1692,
            ltout => OPEN,
            carryin => n12585,
            carryout => n12586,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_12_lut_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53842\,
            in2 => \N__47276\,
            in3 => \N__45114\,
            lcout => n1691,
            ltout => OPEN,
            carryin => n12586,
            carryout => n12587,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_13_lut_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47246\,
            in2 => \N__54244\,
            in3 => \N__45102\,
            lcout => n1690,
            ltout => OPEN,
            carryin => n12587,
            carryout => n12588,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_14_lut_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53846\,
            in2 => \N__47180\,
            in3 => \N__45090\,
            lcout => n1689,
            ltout => OPEN,
            carryin => n12588,
            carryout => n12589,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_15_lut_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45371\,
            in2 => \N__54245\,
            in3 => \N__45081\,
            lcout => n1688,
            ltout => OPEN,
            carryin => n12589,
            carryout => n12590,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1101_16_lut_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__54954\,
            in1 => \N__45167\,
            in2 => \N__52443\,
            in3 => \N__45348\,
            lcout => n1719,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1111_3_lut_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45324\,
            in2 => \N__45617\,
            in3 => \N__47405\,
            lcout => n1727,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12884_4_lut_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47173\,
            in1 => \N__45364\,
            in2 => \N__47220\,
            in3 => \N__52439\,
            lcout => n1653,
            ltout => \n1653_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1112_3_lut_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45294\,
            in2 => \N__45285\,
            in3 => \N__47064\,
            lcout => n1728,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1113_3_lut_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47082\,
            in2 => \N__45264\,
            in3 => \N__45586\,
            lcout => n1729,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1108_3_lut_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__45252\,
            in1 => \N__45155\,
            in2 => \N__45613\,
            in3 => \_gnd_net_\,
            lcout => n1724,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1109_3_lut_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47336\,
            in2 => \N__45219\,
            in3 => \N__45587\,
            lcout => n1725,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12881_1_lut_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45614\,
            in3 => \_gnd_net_\,
            lcout => n15611,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1041_3_lut_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__51969\,
            in1 => \_gnd_net_\,
            in2 => \N__51999\,
            in3 => \N__48877\,
            lcout => n1625_adj_605,
            ltout => \n1625_adj_605_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_122_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47335\,
            in1 => \N__47200\,
            in2 => \N__45714\,
            in3 => \N__47401\,
            lcout => n14502,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1114_3_lut_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45711\,
            in2 => \N__48930\,
            in3 => \N__45597\,
            lcout => n1730,
            ltout => \n1730_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_134_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45684\,
            in3 => \N__45670\,
            lcout => n14514,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47365\,
            lcout => n11_adj_629,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1117_3_lut_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45630\,
            in2 => \N__45615\,
            in3 => \N__48789\,
            lcout => n1733,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12900_1_lut_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45480\,
            lcout => n15630,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1037_3_lut_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__52536\,
            in1 => \N__52509\,
            in2 => \N__48893\,
            in3 => \_gnd_net_\,
            lcout => n1621_adj_601,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_new_i1_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46417\,
            lcout => \quad_counter0.b_new_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56213\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_new_i0_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45822\,
            lcout => \quad_counter0.b_new_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56213\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i707_3_lut_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53017\,
            in2 => \N__49860\,
            in3 => \N__52995\,
            lcout => n1131,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45800\,
            lcout => n32_adj_650,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45758\,
            lcout => n17_adj_635,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i705_3_lut_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__49842\,
            in1 => \_gnd_net_\,
            in2 => \N__52937\,
            in3 => \N__52911\,
            lcout => n1129,
            ltout => \n1129_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_99_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45717\,
            in3 => \N__47536\,
            lcout => n14464,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i706_3_lut_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49841\,
            in2 => \N__52979\,
            in3 => \N__52953\,
            lcout => n1130,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i702_3_lut_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55592\,
            in2 => \N__49868\,
            in3 => \N__55575\,
            lcout => n1126,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i638_3_lut_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45854\,
            in2 => \N__45834\,
            in3 => \N__46008\,
            lcout => n1030,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9957_3_lut_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53083\,
            in2 => \N__53021\,
            in3 => \N__53050\,
            lcout => OPEN,
            ltout => \n11933_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_92_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__52885\,
            in1 => \N__52972\,
            in2 => \N__45936\,
            in3 => \N__52930\,
            lcout => OPEN,
            ltout => \n13728_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12781_4_lut_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__52852\,
            in1 => \N__53377\,
            in2 => \N__45933\,
            in3 => \N__55591\,
            lcout => n1059,
            ltout => \n1059_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i709_3_lut_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__53084\,
            in1 => \_gnd_net_\,
            in2 => \N__45930\,
            in3 => \N__53070\,
            lcout => n1133,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i708_3_lut_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53034\,
            in2 => \N__49867\,
            in3 => \N__53051\,
            lcout => n1132,
            ltout => \n1132_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10042_4_lut_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__47572\,
            in1 => \N__47647\,
            in2 => \N__45927\,
            in3 => \N__47611\,
            lcout => n12019,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_2_lut_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45923\,
            in2 => \_gnd_net_\,
            in3 => \N__45906\,
            lcout => n1001,
            ltout => OPEN,
            carryin => \bfn_13_24_0_\,
            carryout => n12507,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_3_lut_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53785\,
            in2 => \N__45903\,
            in3 => \N__45882\,
            lcout => n1000,
            ltout => OPEN,
            carryin => n12507,
            carryout => n12508,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_4_lut_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__45879\,
            in3 => \N__45858\,
            lcout => n999,
            ltout => OPEN,
            carryin => n12508,
            carryout => n12509,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_5_lut_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53786\,
            in2 => \N__45855\,
            in3 => \N__46110\,
            lcout => n998,
            ltout => OPEN,
            carryin => n12509,
            carryout => n12510,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_6_lut_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__46107\,
            in3 => \N__46074\,
            lcout => n997,
            ltout => OPEN,
            carryin => n12510,
            carryout => n12511,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_7_lut_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__46071\,
            in3 => \N__46044\,
            lcout => n996,
            ltout => OPEN,
            carryin => n12511,
            carryout => n12512,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_8_lut_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53787\,
            in2 => \N__46041\,
            in3 => \N__46017\,
            lcout => n995,
            ltout => OPEN,
            carryin => n12512,
            carryout => n12513,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_632_9_lut_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__53788\,
            in1 => \N__46012\,
            in2 => \N__45975\,
            in3 => \N__45957\,
            lcout => n1026,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i1_1_lut_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45954\,
            lcout => n25_adj_551,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9898_2_lut_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50265\,
            in2 => \_gnd_net_\,
            in3 => \N__50310\,
            lcout => OPEN,
            ltout => \n11872_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_adj_52_LC_13_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__50071\,
            in1 => \N__50191\,
            in2 => \N__45939\,
            in3 => \N__50232\,
            lcout => n10_adj_681,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__49763\,
            in1 => \N__50347\,
            in2 => \N__49736\,
            in3 => \N__49699\,
            lcout => OPEN,
            ltout => \n14034_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__50266\,
            in1 => \_gnd_net_\,
            in2 => \N__46173\,
            in3 => \N__50318\,
            lcout => OPEN,
            ltout => \n14116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_51_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__50117\,
            in1 => \N__50476\,
            in2 => \N__46170\,
            in3 => \N__46167\,
            lcout => n15_adj_680,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_LC_13_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50072\,
            in1 => \N__50233\,
            in2 => \N__50198\,
            in3 => \N__50153\,
            lcout => n10_adj_598,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__51266\,
            in1 => \N__50557\,
            in2 => \N__50397\,
            in3 => \N__51050\,
            lcout => n24_adj_653,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i2_LC_13_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50836\,
            in1 => \N__46161\,
            in2 => \_gnd_net_\,
            in3 => \N__46526\,
            lcout => pwm_setpoint_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i3_LC_13_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50837\,
            in1 => \N__46152\,
            in2 => \_gnd_net_\,
            in3 => \N__46143\,
            lcout => pwm_setpoint_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_70_LC_13_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__50392\,
            in1 => \N__50107\,
            in2 => \N__46131\,
            in3 => \N__50151\,
            lcout => n15_adj_711,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_adj_53_LC_13_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__50670\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51265\,
            lcout => OPEN,
            ltout => \n16_adj_710_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_4_lut_adj_73_LC_13_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50630\,
            in1 => \N__51227\,
            in2 => \N__46122\,
            in3 => \N__46119\,
            lcout => n25_adj_707,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i3_1_lut_LC_13_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46527\,
            lcout => n23_adj_595,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i15_LC_13_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50835\,
            in1 => \N__46499\,
            in2 => \_gnd_net_\,
            in3 => \N__46485\,
            lcout => pwm_setpoint_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.a_new_i1_LC_13_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46461\,
            lcout => a_new_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.i12534_4_lut_LC_13_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__46456\,
            in1 => \N__46424\,
            in2 => \N__46393\,
            in3 => \N__46332\,
            lcout => \quad_counter0.a_prev_N_543\,
            ltout => \quad_counter0.a_prev_N_543_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \quad_counter0.b_prev_52_LC_13_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__46333\,
            in1 => \N__46307\,
            in2 => \N__46281\,
            in3 => \N__46269\,
            lcout => b_prev,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56238\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i2_3_lut_LC_13_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__48080\,
            in1 => \N__48048\,
            in2 => \_gnd_net_\,
            in3 => \N__48009\,
            lcout => \PWM.n13991\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12391_3_lut_4_lut_LC_13_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__46196\,
            in1 => \N__46184\,
            in2 => \N__48138\,
            in3 => \N__48118\,
            lcout => n15121,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i6_LC_13_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50838\,
            in1 => \N__46224\,
            in2 => \_gnd_net_\,
            in3 => \N__47321\,
            lcout => pwm_setpoint_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56238\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i6_3_lut_3_lut_LC_13_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__46197\,
            in1 => \N__46185\,
            in2 => \_gnd_net_\,
            in3 => \N__48119\,
            lcout => n6_adj_656,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i20_1_lut_LC_13_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__46748\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n6_adj_578,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i1_4_lut_LC_13_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__48526\,
            in1 => \N__48394\,
            in2 => \N__47977\,
            in3 => \N__46728\,
            lcout => \PWM.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_80_LC_13_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__47013\,
            in1 => \N__56320\,
            in2 => \N__56405\,
            in3 => \N__46671\,
            lcout => n4_adj_599,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \commutation_state_prev_i1_LC_13_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__56322\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => commutation_state_prev_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56245\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12529_4_lut_LC_13_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111011"
        )
    port map (
            in0 => \N__46664\,
            in1 => \N__46622\,
            in2 => \N__56406\,
            in3 => \N__56321\,
            lcout => n5201,
            ltout => \n5201_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3271_2_lut_LC_13_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__46623\,
            in1 => \_gnd_net_\,
            in2 => \N__46578\,
            in3 => \_gnd_net_\,
            lcout => n5253,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i27_2_lut_LC_13_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46571\,
            in2 => \_gnd_net_\,
            in3 => \N__48289\,
            lcout => n27_adj_671,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i11_4_lut_LC_13_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__48345\,
            in1 => \N__48367\,
            in2 => \N__48270\,
            in3 => \N__48499\,
            lcout => \PWM.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i12_4_lut_LC_13_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50980\,
            in1 => \N__48291\,
            in2 => \N__48210\,
            in3 => \N__48577\,
            lcout => \PWM.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i10_4_lut_LC_13_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__48427\,
            in1 => \N__48550\,
            in2 => \N__48243\,
            in3 => \N__48462\,
            lcout => OPEN,
            ltout => \PWM.n26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i13_4_lut_LC_13_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__48314\,
            in1 => \N__47037\,
            in2 => \N__47031\,
            in3 => \N__50934\,
            lcout => OPEN,
            ltout => \PWM.n29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.i9630_4_lut_LC_13_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__47028\,
            in1 => \N__50951\,
            in2 => \N__47022\,
            in3 => \N__47019\,
            lcout => \PWM.pwm_counter_31__N_407\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \commutation_state_i2_LC_13_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111100000100"
        )
    port map (
            in0 => \N__47007\,
            in1 => \N__56404\,
            in2 => \N__46904\,
            in3 => \N__46959\,
            lcout => commutation_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56251\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \commutation_state_prev_i2_LC_13_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__56403\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => commutation_state_prev_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56251\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \commutation_state_i0_LC_13_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__47006\,
            in1 => \N__46958\,
            in2 => \_gnd_net_\,
            in3 => \N__46903\,
            lcout => commutation_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56255\,
            ce => \N__46845\,
            sr => \N__46836\
        );

    \LessThan_299_i11_2_lut_LC_13_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46829\,
            in2 => \_gnd_net_\,
            in3 => \N__48081\,
            lcout => n11_adj_660,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i29_2_lut_LC_13_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__48266\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46788\,
            lcout => n29_adj_672,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_13_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LessThan_299_i21_2_lut_LC_13_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__48369\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47117\,
            lcout => n21_adj_667,
            ltout => \n21_adj_667_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12473_3_lut_LC_13_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__47118\,
            in1 => \_gnd_net_\,
            in2 => \N__47106\,
            in3 => \N__47103\,
            lcout => n15203,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1039_3_lut_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51905\,
            in2 => \N__48884\,
            in3 => \N__51891\,
            lcout => n1623_adj_603,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1045_3_lut_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52125\,
            in2 => \N__52149\,
            in3 => \N__48861\,
            lcout => n1629_adj_609,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_112_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__52075\,
            in3 => \N__52027\,
            lcout => OPEN,
            ltout => \n14420_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_118_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__51985\,
            in1 => \N__51943\,
            in2 => \N__47085\,
            in3 => \N__51904\,
            lcout => n14426,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1046_3_lut_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51573\,
            in2 => \N__51594\,
            in3 => \N__48862\,
            lcout => n1630_adj_610,
            ltout => \n1630_adj_610_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_123_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__48913\,
            in1 => \N__47056\,
            in2 => \N__47040\,
            in3 => \N__48726\,
            lcout => n13748,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1049_3_lut_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__51678\,
            in1 => \N__51710\,
            in2 => \_gnd_net_\,
            in3 => \N__48860\,
            lcout => n1633_adj_613,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1040_3_lut_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51927\,
            in2 => \N__51953\,
            in3 => \N__48875\,
            lcout => n1624_adj_604,
            ltout => \n1624_adj_604_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_124_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47259\,
            in1 => \N__47245\,
            in2 => \N__47229\,
            in3 => \N__47226\,
            lcout => n14508,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12477_3_lut_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52050\,
            in2 => \N__52077\,
            in3 => \N__48874\,
            lcout => n1627_adj_607,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i971_3_lut_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__51804\,
            in1 => \_gnd_net_\,
            in2 => \N__51834\,
            in3 => \N__48993\,
            lcout => n1523,
            ltout => \n1523_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1038_3_lut_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52554\,
            in2 => \N__47184\,
            in3 => \N__48876\,
            lcout => n1622_adj_602,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_119_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__52141\,
            in1 => \N__52105\,
            in2 => \N__49023\,
            in3 => \N__47157\,
            lcout => OPEN,
            ltout => \n14428_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12864_4_lut_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__52525\,
            in1 => \N__51866\,
            in2 => \N__47151\,
            in3 => \N__52496\,
            lcout => n1554,
            ltout => \n1554_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12861_1_lut_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__47148\,
            in3 => \_gnd_net_\,
            lcout => n15591,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i908_3_lut_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47445\,
            in2 => \N__49188\,
            in3 => \N__52332\,
            lcout => n1428,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i907_3_lut_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49287\,
            in2 => \N__52348\,
            in3 => \N__47436\,
            lcout => n1427,
            ltout => \n1427_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_107_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__47409\,
            in3 => \N__51388\,
            lcout => n14484,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1044_rep_29_3_lut_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__52109\,
            in1 => \N__52089\,
            in2 => \N__48886\,
            in3 => \_gnd_net_\,
            lcout => n1628_adj_608,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i904_3_lut_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47421\,
            in2 => \N__49668\,
            in3 => \N__52336\,
            lcout => n1424,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i23_3_lut_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47385\,
            in1 => \N__49606\,
            in2 => \_gnd_net_\,
            in3 => \N__47370\,
            lcout => n297,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1042_3_lut_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52011\,
            in2 => \N__52035\,
            in3 => \N__48870\,
            lcout => n1626_adj_606,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i7_1_lut_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47322\,
            lcout => n19_adj_591,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_2_lut_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49138\,
            in2 => \_gnd_net_\,
            in3 => \N__47289\,
            lcout => n1401,
            ltout => OPEN,
            carryin => \bfn_14_20_0_\,
            carryout => n12541,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_3_lut_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54890\,
            in2 => \N__49080\,
            in3 => \N__47286\,
            lcout => n1400,
            ltout => OPEN,
            carryin => n12541,
            carryout => n12542,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_4_lut_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__49212\,
            in3 => \N__47454\,
            lcout => n1399,
            ltout => OPEN,
            carryin => n12542,
            carryout => n12543,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_5_lut_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54891\,
            in2 => \N__49233\,
            in3 => \N__47451\,
            lcout => n1398,
            ltout => OPEN,
            carryin => n12543,
            carryout => n12544,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_6_lut_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__53121\,
            in3 => \N__47448\,
            lcout => n1397,
            ltout => OPEN,
            carryin => n12544,
            carryout => n12545,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_7_lut_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__49184\,
            in3 => \N__47439\,
            lcout => n1396,
            ltout => OPEN,
            carryin => n12545,
            carryout => n12546,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_8_lut_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54893\,
            in2 => \N__49286\,
            in3 => \N__47430\,
            lcout => n1395,
            ltout => OPEN,
            carryin => n12546,
            carryout => n12547,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_9_lut_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54892\,
            in2 => \N__49256\,
            in3 => \N__47427\,
            lcout => n1394,
            ltout => OPEN,
            carryin => n12547,
            carryout => n12548,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_10_lut_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54661\,
            in2 => \N__49376\,
            in3 => \N__47424\,
            lcout => n1393,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => n12549,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_11_lut_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54657\,
            in2 => \N__49664\,
            in3 => \N__47412\,
            lcout => n1392,
            ltout => OPEN,
            carryin => n12549,
            carryout => n12550,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_12_lut_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50001\,
            in2 => \N__54952\,
            in3 => \N__47508\,
            lcout => n1391,
            ltout => OPEN,
            carryin => n12550,
            carryout => n12551,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_900_13_lut_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__54662\,
            in1 => \N__47489\,
            in2 => \N__52581\,
            in3 => \N__47505\,
            lcout => n1422,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12823_1_lut_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__52347\,
            in3 => \_gnd_net_\,
            lcout => n15553,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i774_3_lut_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47556\,
            in2 => \N__47580\,
            in3 => \N__49934\,
            lcout => n1230,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i845_3_lut_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__52230\,
            in1 => \N__52248\,
            in2 => \_gnd_net_\,
            in3 => \N__53174\,
            lcout => n1333,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i913_3_lut_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__49139\,
            in1 => \_gnd_net_\,
            in2 => \N__47478\,
            in3 => \N__52327\,
            lcout => n1433,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_96_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__49307\,
            in1 => \_gnd_net_\,
            in2 => \N__49805\,
            in3 => \N__50026\,
            lcout => OPEN,
            ltout => \n14406_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12795_4_lut_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__47469\,
            in1 => \N__47681\,
            in2 => \N__47463\,
            in3 => \N__47460\,
            lcout => n1158,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i773_3_lut_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47520\,
            in2 => \N__47544\,
            in3 => \N__49924\,
            lcout => n1229,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12765_2_lut_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55761\,
            in2 => \_gnd_net_\,
            in3 => \N__47661\,
            lcout => n5215,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i776_3_lut_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47615\,
            in2 => \N__47595\,
            in3 => \N__49923\,
            lcout => n1232,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i777_3_lut_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47625\,
            in1 => \N__47649\,
            in2 => \_gnd_net_\,
            in3 => \N__49922\,
            lcout => n1233,
            ltout => \n1233_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9951_3_lut_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__52246\,
            in1 => \_gnd_net_\,
            in2 => \N__47652\,
            in3 => \N__52177\,
            lcout => n11927,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_2_lut_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47648\,
            in2 => \_gnd_net_\,
            in3 => \N__47619\,
            lcout => n1201,
            ltout => OPEN,
            carryin => \bfn_14_23_0_\,
            carryout => n12522,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_3_lut_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54247\,
            in2 => \N__47616\,
            in3 => \N__47586\,
            lcout => n1200,
            ltout => OPEN,
            carryin => n12522,
            carryout => n12523,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_4_lut_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__49328\,
            in3 => \N__47583\,
            lcout => n1199,
            ltout => OPEN,
            carryin => n12523,
            carryout => n12524,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_5_lut_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54248\,
            in2 => \N__47579\,
            in3 => \N__47547\,
            lcout => n1198,
            ltout => OPEN,
            carryin => n12524,
            carryout => n12525,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_6_lut_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__47543\,
            in3 => \N__47514\,
            lcout => n1197,
            ltout => OPEN,
            carryin => n12525,
            carryout => n12526,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_7_lut_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__49979\,
            in3 => \N__47511\,
            lcout => n1196,
            ltout => OPEN,
            carryin => n12526,
            carryout => n12527,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_8_lut_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49801\,
            in2 => \N__54656\,
            in3 => \N__47757\,
            lcout => n1195,
            ltout => OPEN,
            carryin => n12527,
            carryout => n12528,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_9_lut_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54252\,
            in2 => \N__49311\,
            in3 => \N__47754\,
            lcout => n1194,
            ltout => OPEN,
            carryin => n12528,
            carryout => n12529,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_10_lut_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53789\,
            in2 => \N__50033\,
            in3 => \N__47751\,
            lcout => n1193,
            ltout => OPEN,
            carryin => \bfn_14_24_0_\,
            carryout => n12530,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_766_11_lut_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__53790\,
            in1 => \N__47738\,
            in2 => \N__47682\,
            in3 => \N__47748\,
            lcout => n1224,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12792_1_lut_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49941\,
            lcout => n15522,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i21_3_lut_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__47727\,
            in1 => \_gnd_net_\,
            in2 => \N__47715\,
            in3 => \N__49603\,
            lcout => n299,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i701_3_lut_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49854\,
            in2 => \N__53384\,
            in3 => \N__53355\,
            lcout => n1125,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_3_lut_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__53346\,
            in1 => \N__55716\,
            in2 => \_gnd_net_\,
            in3 => \N__53328\,
            lcout => OPEN,
            ltout => \n20_adj_618_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12_4_lut_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__55629\,
            in1 => \N__53247\,
            in2 => \N__47664\,
            in3 => \N__47904\,
            lcout => n13197,
            ltout => \n13197_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \direction_167_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011000110"
        )
    port map (
            in0 => \N__55760\,
            in1 => \N__51117\,
            in2 => \N__47823\,
            in3 => \N__47805\,
            lcout => direction_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56228\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9624_4_lut_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__47820\,
            in1 => \N__47772\,
            in2 => \N__51049\,
            in3 => \N__47919\,
            lcout => \direction_N_342\,
            ltout => \direction_N_342_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_303_i1_3_lut_LC_14_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47789\,
            in2 => \N__47814\,
            in3 => \N__51115\,
            lcout => n1693,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20_3_lut_LC_14_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51116\,
            in1 => \N__47790\,
            in2 => \_gnd_net_\,
            in3 => \N__47811\,
            lcout => n13675,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9_4_lut_adj_72_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50586\,
            in1 => \N__50418\,
            in2 => \N__50510\,
            in3 => \N__50544\,
            lcout => OPEN,
            ltout => \n23_adj_709_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i831_4_lut_LC_14_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__51039\,
            in1 => \N__47778\,
            in2 => \N__47799\,
            in3 => \N__47796\,
            lcout => \direction_N_340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_adj_71_LC_14_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__51038\,
            in1 => \N__50463\,
            in2 => \N__50705\,
            in3 => \N__51291\,
            lcout => n24_adj_708,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9_4_lut_LC_14_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__50625\,
            in1 => \N__50419\,
            in2 => \N__50676\,
            in3 => \N__50587\,
            lcout => n23_adj_654,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_setpoint_i1_LC_14_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50905\,
            in1 => \N__47766\,
            in2 => \_gnd_net_\,
            in3 => \N__47874\,
            lcout => pwm_setpoint_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56233\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_LC_14_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__50700\,
            in1 => \N__51216\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \n16_adj_679_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_4_lut_LC_14_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__51292\,
            in1 => \N__50505\,
            in2 => \N__47928\,
            in3 => \N__47925\,
            lcout => n25_adj_652,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9_4_lut_adj_76_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__53310\,
            in1 => \N__53289\,
            in2 => \N__55674\,
            in3 => \N__55938\,
            lcout => n22_adj_617,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_2_lut_LC_14_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55650\,
            in2 => \_gnd_net_\,
            in3 => \N__55959\,
            lcout => OPEN,
            ltout => \n16_adj_619_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_4_lut_adj_77_LC_14_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__55698\,
            in1 => \N__53268\,
            in2 => \N__47913\,
            in3 => \N__47910\,
            lcout => n24_adj_616,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_23__I_0_204_inv_0_i17_1_lut_LC_14_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47895\,
            lcout => n9_adj_567,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \unary_minus_13_inv_0_i2_1_lut_LC_14_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47873\,
            lcout => n24_adj_596,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2178_1_lut_LC_14_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__50863\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_setpoint_23__N_195\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM.pwm_counter_664__i0_LC_14_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48173\,
            in2 => \_gnd_net_\,
            in3 => \N__48159\,
            lcout => pwm_counter_0,
            ltout => OPEN,
            carryin => \bfn_14_28_0_\,
            carryout => \PWM.n13022\,
            clk => \N__56246\,
            ce => 'H',
            sr => \N__48702\
        );

    \PWM.pwm_counter_664__i1_LC_14_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48155\,
            in2 => \_gnd_net_\,
            in3 => \N__48141\,
            lcout => pwm_counter_1,
            ltout => OPEN,
            carryin => \PWM.n13022\,
            carryout => \PWM.n13023\,
            clk => \N__56246\,
            ce => 'H',
            sr => \N__48702\
        );

    \PWM.pwm_counter_664__i2_LC_14_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48137\,
            in2 => \_gnd_net_\,
            in3 => \N__48123\,
            lcout => pwm_counter_2,
            ltout => OPEN,
            carryin => \PWM.n13023\,
            carryout => \PWM.n13024\,
            clk => \N__56246\,
            ce => 'H',
            sr => \N__48702\
        );

    \PWM.pwm_counter_664__i3_LC_14_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48120\,
            in2 => \_gnd_net_\,
            in3 => \N__48105\,
            lcout => pwm_counter_3,
            ltout => OPEN,
            carryin => \PWM.n13024\,
            carryout => \PWM.n13025\,
            clk => \N__56246\,
            ce => 'H',
            sr => \N__48702\
        );

    \PWM.pwm_counter_664__i4_LC_14_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48098\,
            in2 => \_gnd_net_\,
            in3 => \N__48084\,
            lcout => pwm_counter_4,
            ltout => OPEN,
            carryin => \PWM.n13025\,
            carryout => \PWM.n13026\,
            clk => \N__56246\,
            ce => 'H',
            sr => \N__48702\
        );

    \PWM.pwm_counter_664__i5_LC_14_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48079\,
            in2 => \_gnd_net_\,
            in3 => \N__48060\,
            lcout => pwm_counter_5,
            ltout => OPEN,
            carryin => \PWM.n13026\,
            carryout => \PWM.n13027\,
            clk => \N__56246\,
            ce => 'H',
            sr => \N__48702\
        );

    \PWM.pwm_counter_664__i6_LC_14_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48049\,
            in2 => \_gnd_net_\,
            in3 => \N__48021\,
            lcout => pwm_counter_6,
            ltout => OPEN,
            carryin => \PWM.n13027\,
            carryout => \PWM.n13028\,
            clk => \N__56246\,
            ce => 'H',
            sr => \N__48702\
        );

    \PWM.pwm_counter_664__i7_LC_14_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48010\,
            in2 => \_gnd_net_\,
            in3 => \N__47982\,
            lcout => pwm_counter_7,
            ltout => OPEN,
            carryin => \PWM.n13028\,
            carryout => \PWM.n13029\,
            clk => \N__56246\,
            ce => 'H',
            sr => \N__48702\
        );

    \PWM.pwm_counter_664__i8_LC_14_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47967\,
            in2 => \_gnd_net_\,
            in3 => \N__47943\,
            lcout => pwm_counter_8,
            ltout => OPEN,
            carryin => \bfn_14_29_0_\,
            carryout => \PWM.n13030\,
            clk => \N__56252\,
            ce => 'H',
            sr => \N__48694\
        );

    \PWM.pwm_counter_664__i9_LC_14_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48393\,
            in2 => \_gnd_net_\,
            in3 => \N__48372\,
            lcout => pwm_counter_9,
            ltout => OPEN,
            carryin => \PWM.n13030\,
            carryout => \PWM.n13031\,
            clk => \N__56252\,
            ce => 'H',
            sr => \N__48694\
        );

    \PWM.pwm_counter_664__i10_LC_14_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48368\,
            in2 => \_gnd_net_\,
            in3 => \N__48348\,
            lcout => pwm_counter_10,
            ltout => OPEN,
            carryin => \PWM.n13031\,
            carryout => \PWM.n13032\,
            clk => \N__56252\,
            ce => 'H',
            sr => \N__48694\
        );

    \PWM.pwm_counter_664__i11_LC_14_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48340\,
            in2 => \_gnd_net_\,
            in3 => \N__48321\,
            lcout => pwm_counter_11,
            ltout => OPEN,
            carryin => \PWM.n13032\,
            carryout => \PWM.n13033\,
            clk => \N__56252\,
            ce => 'H',
            sr => \N__48694\
        );

    \PWM.pwm_counter_664__i12_LC_14_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48313\,
            in2 => \_gnd_net_\,
            in3 => \N__48294\,
            lcout => pwm_counter_12,
            ltout => OPEN,
            carryin => \PWM.n13033\,
            carryout => \PWM.n13034\,
            clk => \N__56252\,
            ce => 'H',
            sr => \N__48694\
        );

    \PWM.pwm_counter_664__i13_LC_14_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48290\,
            in2 => \_gnd_net_\,
            in3 => \N__48273\,
            lcout => pwm_counter_13,
            ltout => OPEN,
            carryin => \PWM.n13034\,
            carryout => \PWM.n13035\,
            clk => \N__56252\,
            ce => 'H',
            sr => \N__48694\
        );

    \PWM.pwm_counter_664__i14_LC_14_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48265\,
            in2 => \_gnd_net_\,
            in3 => \N__48246\,
            lcout => pwm_counter_14,
            ltout => OPEN,
            carryin => \PWM.n13035\,
            carryout => \PWM.n13036\,
            clk => \N__56252\,
            ce => 'H',
            sr => \N__48694\
        );

    \PWM.pwm_counter_664__i15_LC_14_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48235\,
            in2 => \_gnd_net_\,
            in3 => \N__48216\,
            lcout => pwm_counter_15,
            ltout => OPEN,
            carryin => \PWM.n13036\,
            carryout => \PWM.n13037\,
            clk => \N__56252\,
            ce => 'H',
            sr => \N__48694\
        );

    \PWM.pwm_counter_664__i16_LC_14_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48202\,
            in2 => \_gnd_net_\,
            in3 => \N__48180\,
            lcout => pwm_counter_16,
            ltout => OPEN,
            carryin => \bfn_14_30_0_\,
            carryout => \PWM.n13038\,
            clk => \N__56256\,
            ce => 'H',
            sr => \N__48693\
        );

    \PWM.pwm_counter_664__i17_LC_14_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48578\,
            in2 => \_gnd_net_\,
            in3 => \N__48558\,
            lcout => pwm_counter_17,
            ltout => OPEN,
            carryin => \PWM.n13038\,
            carryout => \PWM.n13039\,
            clk => \N__56256\,
            ce => 'H',
            sr => \N__48693\
        );

    \PWM.pwm_counter_664__i18_LC_14_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48554\,
            in2 => \_gnd_net_\,
            in3 => \N__48531\,
            lcout => pwm_counter_18,
            ltout => OPEN,
            carryin => \PWM.n13039\,
            carryout => \PWM.n13040\,
            clk => \N__56256\,
            ce => 'H',
            sr => \N__48693\
        );

    \PWM.pwm_counter_664__i19_LC_14_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48527\,
            in2 => \_gnd_net_\,
            in3 => \N__48507\,
            lcout => pwm_counter_19,
            ltout => OPEN,
            carryin => \PWM.n13040\,
            carryout => \PWM.n13041\,
            clk => \N__56256\,
            ce => 'H',
            sr => \N__48693\
        );

    \PWM.pwm_counter_664__i20_LC_14_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48500\,
            in2 => \_gnd_net_\,
            in3 => \N__48480\,
            lcout => pwm_counter_20,
            ltout => OPEN,
            carryin => \PWM.n13041\,
            carryout => \PWM.n13042\,
            clk => \N__56256\,
            ce => 'H',
            sr => \N__48693\
        );

    \PWM.pwm_counter_664__i21_LC_14_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48463\,
            in2 => \_gnd_net_\,
            in3 => \N__48435\,
            lcout => pwm_counter_21,
            ltout => OPEN,
            carryin => \PWM.n13042\,
            carryout => \PWM.n13043\,
            clk => \N__56256\,
            ce => 'H',
            sr => \N__48693\
        );

    \PWM.pwm_counter_664__i22_LC_14_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48428\,
            in2 => \_gnd_net_\,
            in3 => \N__48408\,
            lcout => pwm_counter_22,
            ltout => OPEN,
            carryin => \PWM.n13043\,
            carryout => \PWM.n13044\,
            clk => \N__56256\,
            ce => 'H',
            sr => \N__48693\
        );

    \PWM.pwm_counter_664__i23_LC_14_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50981\,
            in2 => \_gnd_net_\,
            in3 => \N__48405\,
            lcout => pwm_counter_23,
            ltout => OPEN,
            carryin => \PWM.n13044\,
            carryout => \PWM.n13045\,
            clk => \N__56256\,
            ce => 'H',
            sr => \N__48693\
        );

    \PWM.pwm_counter_664__i24_LC_14_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48672\,
            in2 => \_gnd_net_\,
            in3 => \N__48402\,
            lcout => pwm_counter_24,
            ltout => OPEN,
            carryin => \bfn_14_31_0_\,
            carryout => \PWM.n13046\,
            clk => \N__56257\,
            ce => 'H',
            sr => \N__48695\
        );

    \PWM.pwm_counter_664__i25_LC_14_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48609\,
            in2 => \_gnd_net_\,
            in3 => \N__48399\,
            lcout => pwm_counter_25,
            ltout => OPEN,
            carryin => \PWM.n13046\,
            carryout => \PWM.n13047\,
            clk => \N__56257\,
            ce => 'H',
            sr => \N__48695\
        );

    \PWM.pwm_counter_664__i26_LC_14_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48633\,
            in2 => \_gnd_net_\,
            in3 => \N__48720\,
            lcout => pwm_counter_26,
            ltout => OPEN,
            carryin => \PWM.n13047\,
            carryout => \PWM.n13048\,
            clk => \N__56257\,
            ce => 'H',
            sr => \N__48695\
        );

    \PWM.pwm_counter_664__i27_LC_14_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48647\,
            in2 => \_gnd_net_\,
            in3 => \N__48717\,
            lcout => pwm_counter_27,
            ltout => OPEN,
            carryin => \PWM.n13048\,
            carryout => \PWM.n13049\,
            clk => \N__56257\,
            ce => 'H',
            sr => \N__48695\
        );

    \PWM.pwm_counter_664__i28_LC_14_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48594\,
            in2 => \_gnd_net_\,
            in3 => \N__48714\,
            lcout => pwm_counter_28,
            ltout => OPEN,
            carryin => \PWM.n13049\,
            carryout => \PWM.n13050\,
            clk => \N__56257\,
            ce => 'H',
            sr => \N__48695\
        );

    \PWM.pwm_counter_664__i29_LC_14_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48660\,
            in2 => \_gnd_net_\,
            in3 => \N__48711\,
            lcout => pwm_counter_29,
            ltout => OPEN,
            carryin => \PWM.n13050\,
            carryout => \PWM.n13051\,
            clk => \N__56257\,
            ce => 'H',
            sr => \N__48695\
        );

    \PWM.pwm_counter_664__i30_LC_14_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48621\,
            in2 => \_gnd_net_\,
            in3 => \N__48708\,
            lcout => pwm_counter_30,
            ltout => OPEN,
            carryin => \PWM.n13051\,
            carryout => \PWM.n13052\,
            clk => \N__56257\,
            ce => 'H',
            sr => \N__48695\
        );

    \PWM.pwm_counter_664__i31_LC_14_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50952\,
            in2 => \_gnd_net_\,
            in3 => \N__48705\,
            lcout => pwm_counter_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56257\,
            ce => 'H',
            sr => \N__48695\
        );

    \i5_4_lut_LC_14_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__48671\,
            in1 => \N__48659\,
            in2 => \N__48648\,
            in3 => \N__48632\,
            lcout => OPEN,
            ltout => \n12_adj_615_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_LC_14_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__48620\,
            in1 => \N__48608\,
            in2 => \N__48597\,
            in3 => \N__48593\,
            lcout => n5180,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1047_3_lut_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51606\,
            in2 => \N__48885\,
            in3 => \N__51626\,
            lcout => n1631_adj_611,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i973_3_lut_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51333\,
            in2 => \N__49007\,
            in3 => \N__51309\,
            lcout => n1525,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i1048_3_lut_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51662\,
            in2 => \N__51642\,
            in3 => \N__48866\,
            lcout => n1632_adj_612,
            ltout => \n1632_adj_612_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9943_3_lut_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48787\,
            in2 => \N__48759\,
            in3 => \N__48742\,
            lcout => n11919,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i981_3_lut_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50754\,
            in1 => \N__50718\,
            in2 => \_gnd_net_\,
            in3 => \N__48976\,
            lcout => n1533,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i972_3_lut_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__51855\,
            in1 => \_gnd_net_\,
            in2 => \N__48999\,
            in3 => \N__51843\,
            lcout => n1524,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i970_3_lut_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51791\,
            in2 => \N__51765\,
            in3 => \N__48987\,
            lcout => n1522,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i978_3_lut_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51476\,
            in2 => \N__49000\,
            in3 => \N__51450\,
            lcout => n1530,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i976_rep_49_3_lut_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48972\,
            in2 => \N__52281\,
            in3 => \N__51408\,
            lcout => n1528,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i974_3_lut_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__51356\,
            in1 => \_gnd_net_\,
            in2 => \N__48998\,
            in3 => \N__51342\,
            lcout => n1526,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i980_3_lut_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__51519\,
            in1 => \_gnd_net_\,
            in2 => \N__51557\,
            in3 => \N__48980\,
            lcout => n1532,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i975_3_lut_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51392\,
            in2 => \N__48997\,
            in3 => \N__51372\,
            lcout => n1527,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12842_1_lut_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48991\,
            lcout => n15572,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i905_3_lut_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49050\,
            in2 => \N__49380\,
            in3 => \N__52343\,
            lcout => n1425,
            ltout => \n1425_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_110_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__51325\,
            in1 => \N__51815\,
            in2 => \N__49041\,
            in3 => \N__49038\,
            lcout => OPEN,
            ltout => \n14490_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12845_4_lut_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__51728\,
            in1 => \N__51781\,
            in2 => \N__49032\,
            in3 => \N__49101\,
            lcout => n1455,
            ltout => \n1455_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i979_3_lut_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__51489\,
            in1 => \_gnd_net_\,
            in2 => \N__49029\,
            in3 => \N__51503\,
            lcout => n1531,
            ltout => \n1531_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10020_4_lut_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__51658\,
            in1 => \N__51706\,
            in2 => \N__49026\,
            in3 => \N__51622\,
            lcout => n11997,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i977_3_lut_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51420\,
            in2 => \N__51440\,
            in3 => \N__48992\,
            lcout => n1529,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i906_3_lut_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49152\,
            in2 => \N__49260\,
            in3 => \N__52342\,
            lcout => n1426,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i903_3_lut_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50000\,
            in2 => \N__52349\,
            in3 => \N__49146\,
            lcout => n1423,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9949_3_lut_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49140\,
            in2 => \N__49079\,
            in3 => \N__49208\,
            lcout => OPEN,
            ltout => \n11925_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_106_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__53113\,
            in1 => \N__49225\,
            in2 => \N__49113\,
            in3 => \N__49177\,
            lcout => n13720,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i910_3_lut_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49110\,
            in2 => \N__49232\,
            in3 => \N__52338\,
            lcout => n1430,
            ltout => \n1430_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_108_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__52276\,
            in1 => \N__51466\,
            in2 => \N__49104\,
            in3 => \N__49056\,
            lcout => n13739,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12826_4_lut_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__49999\,
            in1 => \N__49266\,
            in2 => \N__52577\,
            in3 => \N__49095\,
            lcout => n1356,
            ltout => \n1356_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i912_3_lut_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49089\,
            in2 => \N__49083\,
            in3 => \N__49075\,
            lcout => n1432,
            ltout => \n1432_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9947_3_lut_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50743\,
            in2 => \N__49059\,
            in3 => \N__51538\,
            lcout => n11923,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i840_3_lut_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__52755\,
            in1 => \_gnd_net_\,
            in2 => \N__53180\,
            in3 => \N__52781\,
            lcout => n1328,
            ltout => \n1328_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_105_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__49249\,
            in1 => \N__49369\,
            in2 => \N__49269\,
            in3 => \N__49657\,
            lcout => n14414,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i839_3_lut_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52719\,
            in2 => \N__52746\,
            in3 => \N__53166\,
            lcout => n1327,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i843_3_lut_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52178\,
            in2 => \N__53179\,
            in3 => \N__52158\,
            lcout => n1331,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i844_3_lut_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52194\,
            in2 => \N__52214\,
            in3 => \N__53162\,
            lcout => n1332,
            ltout => \n1332_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i911_3_lut_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__49197\,
            in1 => \_gnd_net_\,
            in2 => \N__49191\,
            in3 => \N__52331\,
            lcout => n1431,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i841_3_lut_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52794\,
            in2 => \N__52821\,
            in3 => \N__53167\,
            lcout => n1329,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_101_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__52813\,
            in1 => \N__52774\,
            in2 => \N__53221\,
            in3 => \N__49161\,
            lcout => OPEN,
            ltout => \n13723_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12810_4_lut_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__52652\,
            in1 => \N__49344\,
            in2 => \N__49155\,
            in3 => \N__52601\,
            lcout => n1257,
            ltout => \n1257_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i837_3_lut_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__52679\,
            in1 => \_gnd_net_\,
            in2 => \N__49671\,
            in3 => \N__52665\,
            lcout => n1325,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12807_1_lut_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53171\,
            lcout => n15537,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_mux_3_i22_3_lut_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__49641\,
            in1 => \N__49622\,
            in2 => \_gnd_net_\,
            in3 => \N__52416\,
            lcout => n298,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i838_3_lut_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52692\,
            in2 => \N__52710\,
            in3 => \N__53172\,
            lcout => n1326,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i771_3_lut_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49806\,
            in2 => \N__49943\,
            in3 => \N__49353\,
            lcout => n1227,
            ltout => \n1227_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_100_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52732\,
            in2 => \N__49347\,
            in3 => \N__52678\,
            lcout => n14476,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i775_3_lut_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49338\,
            in2 => \N__49332\,
            in3 => \N__49928\,
            lcout => n1231,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i703_3_lut_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52859\,
            in2 => \N__49876\,
            in3 => \N__52833\,
            lcout => n1127,
            ltout => \n1127_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i770_3_lut_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49296\,
            in2 => \N__49290\,
            in3 => \N__49929\,
            lcout => n1226,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i769_3_lut_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50034\,
            in2 => \N__49942\,
            in3 => \N__50010\,
            lcout => n1225,
            ltout => \n1225_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i836_3_lut_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__53175\,
            in1 => \N__52641\,
            in2 => \N__50004\,
            in3 => \_gnd_net_\,
            lcout => n1324,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i772_3_lut_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49983\,
            in2 => \N__49962\,
            in3 => \N__49930\,
            lcout => n1228,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i704_3_lut_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52895\,
            in2 => \N__49875\,
            in3 => \N__52869\,
            lcout => n1128,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_305_1_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51118\,
            in2 => \N__51164\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_25_0_\,
            carryout => n12449,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i0_LC_15_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49762\,
            in2 => \N__49782\,
            in3 => \N__49743\,
            lcout => encoder0_position_target_0,
            ltout => OPEN,
            carryin => n12449,
            carryout => n12450,
            clk => \N__56234\,
            ce => \N__55881\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i1_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51119\,
            in2 => \N__49735\,
            in3 => \N__49707\,
            lcout => encoder0_position_target_1,
            ltout => OPEN,
            carryin => n12450,
            carryout => n12451,
            clk => \N__56234\,
            ce => \N__55881\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i2_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51125\,
            in2 => \N__49703\,
            in3 => \N__49674\,
            lcout => encoder0_position_target_2,
            ltout => OPEN,
            carryin => n12451,
            carryout => n12452,
            clk => \N__56234\,
            ce => \N__55881\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i3_LC_15_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51120\,
            in2 => \N__50351\,
            in3 => \N__50322\,
            lcout => encoder0_position_target_3,
            ltout => OPEN,
            carryin => n12452,
            carryout => n12453,
            clk => \N__56234\,
            ce => \N__55881\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i4_LC_15_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51126\,
            in2 => \N__50317\,
            in3 => \N__50277\,
            lcout => encoder0_position_target_4,
            ltout => OPEN,
            carryin => n12453,
            carryout => n12454,
            clk => \N__56234\,
            ce => \N__55881\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i5_LC_15_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51121\,
            in2 => \N__50270\,
            in3 => \N__50241\,
            lcout => encoder0_position_target_5,
            ltout => OPEN,
            carryin => n12454,
            carryout => n12455,
            clk => \N__56234\,
            ce => \N__55881\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i6_LC_15_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51127\,
            in2 => \N__50237\,
            in3 => \N__50205\,
            lcout => encoder0_position_target_6,
            ltout => OPEN,
            carryin => n12455,
            carryout => n12456,
            clk => \N__56234\,
            ce => \N__55881\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i7_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50181\,
            in2 => \N__51165\,
            in3 => \N__50160\,
            lcout => encoder0_position_target_7,
            ltout => OPEN,
            carryin => \bfn_15_26_0_\,
            carryout => n12457,
            clk => \N__56239\,
            ce => \N__55916\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i8_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51131\,
            in2 => \N__50152\,
            in3 => \N__50121\,
            lcout => encoder0_position_target_8,
            ltout => OPEN,
            carryin => n12457,
            carryout => n12458,
            clk => \N__56239\,
            ce => \N__55916\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i9_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50106\,
            in2 => \N__51166\,
            in3 => \N__50079\,
            lcout => encoder0_position_target_9,
            ltout => OPEN,
            carryin => n12458,
            carryout => n12459,
            clk => \N__56239\,
            ce => \N__55916\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i10_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51135\,
            in2 => \N__50070\,
            in3 => \N__50037\,
            lcout => encoder0_position_target_10,
            ltout => OPEN,
            carryin => n12459,
            carryout => n12460,
            clk => \N__56239\,
            ce => \N__55916\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i11_LC_15_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50704\,
            in2 => \N__51167\,
            in3 => \N__50679\,
            lcout => encoder0_position_target_11,
            ltout => OPEN,
            carryin => n12460,
            carryout => n12461,
            clk => \N__56239\,
            ce => \N__55916\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i12_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51139\,
            in2 => \N__50675\,
            in3 => \N__50640\,
            lcout => encoder0_position_target_12,
            ltout => OPEN,
            carryin => n12461,
            carryout => n12462,
            clk => \N__56239\,
            ce => \N__55916\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i13_LC_15_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50629\,
            in2 => \N__51168\,
            in3 => \N__50601\,
            lcout => encoder0_position_target_13,
            ltout => OPEN,
            carryin => n12462,
            carryout => n12463,
            clk => \N__56239\,
            ce => \N__55916\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i14_LC_15_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51143\,
            in2 => \N__50597\,
            in3 => \N__50568\,
            lcout => encoder0_position_target_14,
            ltout => OPEN,
            carryin => n12463,
            carryout => n12464,
            clk => \N__56239\,
            ce => \N__55916\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i15_LC_15_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51169\,
            in2 => \N__50558\,
            in3 => \N__50520\,
            lcout => encoder0_position_target_15,
            ltout => OPEN,
            carryin => \bfn_15_27_0_\,
            carryout => n12465,
            clk => \N__56247\,
            ce => \N__55898\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i16_LC_15_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50509\,
            in2 => \N__51186\,
            in3 => \N__50484\,
            lcout => encoder0_position_target_16,
            ltout => OPEN,
            carryin => n12465,
            carryout => n12466,
            clk => \N__56247\,
            ce => \N__55898\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i17_LC_15_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51173\,
            in2 => \N__50477\,
            in3 => \N__50439\,
            lcout => encoder0_position_target_17,
            ltout => OPEN,
            carryin => n12466,
            carryout => n12467,
            clk => \N__56247\,
            ce => \N__55898\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i18_LC_15_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50429\,
            in2 => \N__51187\,
            in3 => \N__50400\,
            lcout => encoder0_position_target_18,
            ltout => OPEN,
            carryin => n12467,
            carryout => n12468,
            clk => \N__56247\,
            ce => \N__55898\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i19_LC_15_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51177\,
            in2 => \N__50391\,
            in3 => \N__50355\,
            lcout => encoder0_position_target_19,
            ltout => OPEN,
            carryin => n12468,
            carryout => n12469,
            clk => \N__56247\,
            ce => \N__55898\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i20_LC_15_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51296\,
            in2 => \N__51188\,
            in3 => \N__51273\,
            lcout => encoder0_position_target_20,
            ltout => OPEN,
            carryin => n12469,
            carryout => n12470,
            clk => \N__56247\,
            ce => \N__55898\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i21_LC_15_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51181\,
            in2 => \N__51264\,
            in3 => \N__51231\,
            lcout => encoder0_position_target_21,
            ltout => OPEN,
            carryin => n12470,
            carryout => n12471,
            clk => \N__56247\,
            ce => \N__55898\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i22_LC_15_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51220\,
            in2 => \N__51189\,
            in3 => \N__51192\,
            lcout => encoder0_position_target_22,
            ltout => OPEN,
            carryin => n12471,
            carryout => n12472,
            clk => \N__56247\,
            ce => \N__55898\,
            sr => \_gnd_net_\
        );

    \encoder0_position_target_i0_i23_LC_15_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__51185\,
            in1 => \N__51037\,
            in2 => \_gnd_net_\,
            in3 => \N__51057\,
            lcout => encoder0_position_target_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56253\,
            ce => \N__55911\,
            sr => \_gnd_net_\
        );

    \PWM.pwm_out_12_LC_15_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__50997\,
            in1 => \N__50982\,
            in2 => \_gnd_net_\,
            in3 => \N__50964\,
            lcout => pwm_out,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56258\,
            ce => 'H',
            sr => \N__50919\
        );

    \i1_2_lut_adj_44_LC_15_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50950\,
            in2 => \_gnd_net_\,
            in3 => \N__50933\,
            lcout => n5182,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dir_160_LC_15_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50909\,
            lcout => dir,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56259\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_2_lut_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50750\,
            in2 => \_gnd_net_\,
            in3 => \N__50712\,
            lcout => n1501,
            ltout => OPEN,
            carryin => \bfn_16_17_0_\,
            carryout => n12552,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_3_lut_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55128\,
            in2 => \N__51558\,
            in3 => \N__51513\,
            lcout => n1500,
            ltout => OPEN,
            carryin => n12552,
            carryout => n12553,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_4_lut_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51510\,
            in3 => \N__51480\,
            lcout => n1499,
            ltout => OPEN,
            carryin => n12553,
            carryout => n12554,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_5_lut_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55129\,
            in2 => \N__51477\,
            in3 => \N__51444\,
            lcout => n1498,
            ltout => OPEN,
            carryin => n12554,
            carryout => n12555,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_6_lut_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51441\,
            in3 => \N__51411\,
            lcout => n1497,
            ltout => OPEN,
            carryin => n12555,
            carryout => n12556,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_7_lut_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__52280\,
            in3 => \N__51402\,
            lcout => n1496,
            ltout => OPEN,
            carryin => n12556,
            carryout => n12557,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_8_lut_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55131\,
            in2 => \N__51399\,
            in3 => \N__51366\,
            lcout => n1495,
            ltout => OPEN,
            carryin => n12557,
            carryout => n12558,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_9_lut_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55130\,
            in2 => \N__51363\,
            in3 => \N__51336\,
            lcout => n1494,
            ltout => OPEN,
            carryin => n12558,
            carryout => n12559,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_10_lut_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55121\,
            in2 => \N__51332\,
            in3 => \N__51303\,
            lcout => n1493,
            ltout => OPEN,
            carryin => \bfn_16_18_0_\,
            carryout => n12560,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_11_lut_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51854\,
            in2 => \N__55288\,
            in3 => \N__51837\,
            lcout => n1492,
            ltout => OPEN,
            carryin => n12560,
            carryout => n12561,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_12_lut_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55125\,
            in2 => \N__51833\,
            in3 => \N__51795\,
            lcout => n1491,
            ltout => OPEN,
            carryin => n12561,
            carryout => n12562,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_13_lut_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55126\,
            in2 => \N__51792\,
            in3 => \N__51756\,
            lcout => n1490,
            ltout => OPEN,
            carryin => n12562,
            carryout => n12563,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_967_14_lut_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__55127\,
            in1 => \N__51746\,
            in2 => \N__51735\,
            in3 => \N__51714\,
            lcout => n1521,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_2_lut_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51711\,
            in2 => \_gnd_net_\,
            in3 => \N__51666\,
            lcout => n1601,
            ltout => OPEN,
            carryin => \bfn_16_19_0_\,
            carryout => n12564,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_3_lut_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55117\,
            in2 => \N__51663\,
            in3 => \N__51630\,
            lcout => n1600,
            ltout => OPEN,
            carryin => n12564,
            carryout => n12565,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_4_lut_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__51627\,
            in3 => \N__51597\,
            lcout => n1599,
            ltout => OPEN,
            carryin => n12565,
            carryout => n12566,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_5_lut_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55118\,
            in2 => \N__51590\,
            in3 => \N__51561\,
            lcout => n1598,
            ltout => OPEN,
            carryin => n12566,
            carryout => n12567,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_6_lut_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__52148\,
            in3 => \N__52113\,
            lcout => n1597,
            ltout => OPEN,
            carryin => n12567,
            carryout => n12568,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_7_lut_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__52110\,
            in3 => \N__52080\,
            lcout => n1596,
            ltout => OPEN,
            carryin => n12568,
            carryout => n12569,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_8_lut_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55120\,
            in2 => \N__52076\,
            in3 => \N__52038\,
            lcout => n1595,
            ltout => OPEN,
            carryin => n12569,
            carryout => n12570,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_9_lut_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55119\,
            in2 => \N__52034\,
            in3 => \N__52002\,
            lcout => n1594,
            ltout => OPEN,
            carryin => n12570,
            carryout => n12571,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_10_lut_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51992\,
            in2 => \N__55278\,
            in3 => \N__51957\,
            lcout => n1593,
            ltout => OPEN,
            carryin => \bfn_16_20_0_\,
            carryout => n12572,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_11_lut_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55091\,
            in2 => \N__51954\,
            in3 => \N__51915\,
            lcout => n1592,
            ltout => OPEN,
            carryin => n12572,
            carryout => n12573,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_12_lut_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55096\,
            in2 => \N__51912\,
            in3 => \N__51879\,
            lcout => n1591,
            ltout => OPEN,
            carryin => n12573,
            carryout => n12574,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_13_lut_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55092\,
            in2 => \N__51876\,
            in3 => \N__52539\,
            lcout => n1590,
            ltout => OPEN,
            carryin => n12574,
            carryout => n12575,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_14_lut_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52532\,
            in2 => \N__55279\,
            in3 => \N__52500\,
            lcout => n1589,
            ltout => OPEN,
            carryin => n12575,
            carryout => n12576,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_1034_15_lut_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__55097\,
            in1 => \N__52497\,
            in2 => \N__52475\,
            in3 => \N__52446\,
            lcout => n1620_adj_600,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52409\,
            lcout => n12_adj_630,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i909_3_lut_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53114\,
            in2 => \N__52371\,
            in3 => \N__52337\,
            lcout => n1429,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_2_lut_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52247\,
            in2 => \_gnd_net_\,
            in3 => \N__52221\,
            lcout => n1301,
            ltout => OPEN,
            carryin => \bfn_16_21_0_\,
            carryout => n12531,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_3_lut_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54650\,
            in2 => \N__52218\,
            in3 => \N__52188\,
            lcout => n1300,
            ltout => OPEN,
            carryin => n12531,
            carryout => n12532,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_4_lut_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__52185\,
            in3 => \N__52152\,
            lcout => n1299,
            ltout => OPEN,
            carryin => n12532,
            carryout => n12533,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_5_lut_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54651\,
            in2 => \N__53223\,
            in3 => \N__52824\,
            lcout => n1298,
            ltout => OPEN,
            carryin => n12533,
            carryout => n12534,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_6_lut_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__52820\,
            in3 => \N__52788\,
            lcout => n1297,
            ltout => OPEN,
            carryin => n12534,
            carryout => n12535,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_7_lut_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__52785\,
            in3 => \N__52749\,
            lcout => n1296,
            ltout => OPEN,
            carryin => n12535,
            carryout => n12536,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_8_lut_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54653\,
            in2 => \N__52745\,
            in3 => \N__52713\,
            lcout => n1295,
            ltout => OPEN,
            carryin => n12536,
            carryout => n12537,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_9_lut_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54652\,
            in2 => \N__52709\,
            in3 => \N__52686\,
            lcout => n1294,
            ltout => OPEN,
            carryin => n12537,
            carryout => n12538,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_10_lut_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54647\,
            in2 => \N__52683\,
            in3 => \N__52659\,
            lcout => n1293,
            ltout => OPEN,
            carryin => \bfn_16_22_0_\,
            carryout => n12539,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_11_lut_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54648\,
            in2 => \N__52656\,
            in3 => \N__52635\,
            lcout => n1292,
            ltout => OPEN,
            carryin => n12539,
            carryout => n12540,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_833_12_lut_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__54649\,
            in1 => \N__52619\,
            in2 => \N__52608\,
            in3 => \N__52584\,
            lcout => n1323,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_i842_3_lut_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53229\,
            in2 => \N__53222\,
            in3 => \N__53173\,
            lcout => n1330,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_2_lut_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53091\,
            in2 => \_gnd_net_\,
            in3 => \N__53058\,
            lcout => n1101,
            ltout => OPEN,
            carryin => \bfn_16_23_0_\,
            carryout => n12514,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_3_lut_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54643\,
            in2 => \N__53055\,
            in3 => \N__53025\,
            lcout => n1100,
            ltout => OPEN,
            carryin => n12514,
            carryout => n12515,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_4_lut_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__53022\,
            in3 => \N__52983\,
            lcout => n1099,
            ltout => OPEN,
            carryin => n12515,
            carryout => n12516,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_5_lut_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54644\,
            in2 => \N__52980\,
            in3 => \N__52941\,
            lcout => n1098,
            ltout => OPEN,
            carryin => n12516,
            carryout => n12517,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_6_lut_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__52938\,
            in3 => \N__52899\,
            lcout => n1097,
            ltout => OPEN,
            carryin => n12517,
            carryout => n12518,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_7_lut_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__52896\,
            in3 => \N__52863\,
            lcout => n1096,
            ltout => OPEN,
            carryin => n12518,
            carryout => n12519,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_8_lut_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54646\,
            in2 => \N__52860\,
            in3 => \N__52827\,
            lcout => n1095,
            ltout => OPEN,
            carryin => n12519,
            carryout => n12520,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_9_lut_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54645\,
            in2 => \N__55599\,
            in3 => \N__55566\,
            lcout => n1094,
            ltout => OPEN,
            carryin => n12520,
            carryout => n12521,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \encoder0_position_31__I_0_add_699_10_lut_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53791\,
            in2 => \N__53385\,
            in3 => \N__53358\,
            lcout => n1093,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sweep_counter_660_661__i1_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53345\,
            in2 => \_gnd_net_\,
            in3 => \N__53331\,
            lcout => sweep_counter_0,
            ltout => OPEN,
            carryin => \bfn_16_25_0_\,
            carryout => n13053,
            clk => \N__56240\,
            ce => 'H',
            sr => \N__55897\
        );

    \sweep_counter_660_661__i2_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53327\,
            in2 => \_gnd_net_\,
            in3 => \N__53313\,
            lcout => sweep_counter_1,
            ltout => OPEN,
            carryin => n13053,
            carryout => n13054,
            clk => \N__56240\,
            ce => 'H',
            sr => \N__55897\
        );

    \sweep_counter_660_661__i3_LC_16_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53309\,
            in2 => \_gnd_net_\,
            in3 => \N__53292\,
            lcout => sweep_counter_2,
            ltout => OPEN,
            carryin => n13054,
            carryout => n13055,
            clk => \N__56240\,
            ce => 'H',
            sr => \N__55897\
        );

    \sweep_counter_660_661__i4_LC_16_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53285\,
            in2 => \_gnd_net_\,
            in3 => \N__53271\,
            lcout => sweep_counter_3,
            ltout => OPEN,
            carryin => n13055,
            carryout => n13056,
            clk => \N__56240\,
            ce => 'H',
            sr => \N__55897\
        );

    \sweep_counter_660_661__i5_LC_16_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53264\,
            in2 => \_gnd_net_\,
            in3 => \N__53250\,
            lcout => sweep_counter_4,
            ltout => OPEN,
            carryin => n13056,
            carryout => n13057,
            clk => \N__56240\,
            ce => 'H',
            sr => \N__55897\
        );

    \sweep_counter_660_661__i6_LC_16_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53246\,
            in2 => \_gnd_net_\,
            in3 => \N__53232\,
            lcout => sweep_counter_5,
            ltout => OPEN,
            carryin => n13057,
            carryout => n13058,
            clk => \N__56240\,
            ce => 'H',
            sr => \N__55897\
        );

    \sweep_counter_660_661__i7_LC_16_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55715\,
            in2 => \_gnd_net_\,
            in3 => \N__55701\,
            lcout => sweep_counter_6,
            ltout => OPEN,
            carryin => n13058,
            carryout => n13059,
            clk => \N__56240\,
            ce => 'H',
            sr => \N__55897\
        );

    \sweep_counter_660_661__i8_LC_16_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55694\,
            in2 => \_gnd_net_\,
            in3 => \N__55680\,
            lcout => sweep_counter_7,
            ltout => OPEN,
            carryin => n13059,
            carryout => n13060,
            clk => \N__56240\,
            ce => 'H',
            sr => \N__55897\
        );

    \sweep_counter_660_661__i9_LC_16_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55835\,
            in2 => \_gnd_net_\,
            in3 => \N__55677\,
            lcout => sweep_counter_8,
            ltout => OPEN,
            carryin => \bfn_16_26_0_\,
            carryout => n13061,
            clk => \N__56248\,
            ce => 'H',
            sr => \N__55912\
        );

    \sweep_counter_660_661__i10_LC_16_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55667\,
            in2 => \_gnd_net_\,
            in3 => \N__55653\,
            lcout => sweep_counter_9,
            ltout => OPEN,
            carryin => n13061,
            carryout => n13062,
            clk => \N__56248\,
            ce => 'H',
            sr => \N__55912\
        );

    \sweep_counter_660_661__i11_LC_16_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55646\,
            in2 => \_gnd_net_\,
            in3 => \N__55632\,
            lcout => sweep_counter_10,
            ltout => OPEN,
            carryin => n13062,
            carryout => n13063,
            clk => \N__56248\,
            ce => 'H',
            sr => \N__55912\
        );

    \sweep_counter_660_661__i12_LC_16_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55625\,
            in2 => \_gnd_net_\,
            in3 => \N__55611\,
            lcout => sweep_counter_11,
            ltout => OPEN,
            carryin => n13063,
            carryout => n13064,
            clk => \N__56248\,
            ce => 'H',
            sr => \N__55912\
        );

    \sweep_counter_660_661__i13_LC_16_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55775\,
            in2 => \_gnd_net_\,
            in3 => \N__55608\,
            lcout => sweep_counter_12,
            ltout => OPEN,
            carryin => n13064,
            carryout => n13065,
            clk => \N__56248\,
            ce => 'H',
            sr => \N__55912\
        );

    \sweep_counter_660_661__i14_LC_16_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55805\,
            in2 => \_gnd_net_\,
            in3 => \N__55605\,
            lcout => sweep_counter_13,
            ltout => OPEN,
            carryin => n13065,
            carryout => n13066,
            clk => \N__56248\,
            ce => 'H',
            sr => \N__55912\
        );

    \sweep_counter_660_661__i15_LC_16_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55820\,
            in2 => \_gnd_net_\,
            in3 => \N__55602\,
            lcout => sweep_counter_14,
            ltout => OPEN,
            carryin => n13066,
            carryout => n13067,
            clk => \N__56248\,
            ce => 'H',
            sr => \N__55912\
        );

    \sweep_counter_660_661__i16_LC_16_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55955\,
            in2 => \_gnd_net_\,
            in3 => \N__55941\,
            lcout => sweep_counter_15,
            ltout => OPEN,
            carryin => n13067,
            carryout => n13068,
            clk => \N__56248\,
            ce => 'H',
            sr => \N__55912\
        );

    \sweep_counter_660_661__i17_LC_16_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55937\,
            in2 => \_gnd_net_\,
            in3 => \N__55923\,
            lcout => sweep_counter_16,
            ltout => OPEN,
            carryin => \bfn_16_27_0_\,
            carryout => n13069,
            clk => \N__56254\,
            ce => 'H',
            sr => \N__55917\
        );

    \sweep_counter_660_661__i18_LC_16_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55791\,
            in2 => \_gnd_net_\,
            in3 => \N__55920\,
            lcout => sweep_counter_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56254\,
            ce => 'H',
            sr => \N__55917\
        );

    \i1_2_lut_adj_74_LC_16_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55836\,
            in2 => \_gnd_net_\,
            in3 => \N__55821\,
            lcout => OPEN,
            ltout => \n6_adj_712_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_adj_75_LC_16_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__55806\,
            in1 => \N__55790\,
            in2 => \N__55779\,
            in3 => \N__55776\,
            lcout => n13968,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GHC_174_LC_16_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110000010"
        )
    port map (
            in0 => \N__56353\,
            in1 => \N__56516\,
            in2 => \N__56439\,
            in3 => \N__56328\,
            lcout => \GHC\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56260\,
            ce => \N__56056\,
            sr => \N__56029\
        );

    \GHB_172_LC_17_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100000000011"
        )
    port map (
            in0 => \N__56515\,
            in1 => \N__56323\,
            in2 => \N__56440\,
            in3 => \N__56354\,
            lcout => \GHB\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56261\,
            ce => \N__56063\,
            sr => \N__56030\
        );

    \i9546_2_lut_LC_17_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55994\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55734\,
            lcout => \INHC_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9545_2_lut_LC_17_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55993\,
            in2 => \_gnd_net_\,
            in3 => \N__56571\,
            lcout => \INHB_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GHA_170_LC_18_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010010011000"
        )
    port map (
            in0 => \N__56324\,
            in1 => \N__56355\,
            in2 => \N__56441\,
            in3 => \N__56513\,
            lcout => \GHA\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56262\,
            ce => \N__56064\,
            sr => \N__56034\
        );

    \GLA_171_LC_18_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111000010"
        )
    port map (
            in0 => \N__56512\,
            in1 => \N__56431\,
            in2 => \N__56363\,
            in3 => \N__56326\,
            lcout => \INLA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56262\,
            ce => \N__56064\,
            sr => \N__56034\
        );

    \GLB_173_LC_18_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011000010100"
        )
    port map (
            in0 => \N__56325\,
            in1 => \N__56359\,
            in2 => \N__56442\,
            in3 => \N__56514\,
            lcout => \INLB_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56262\,
            ce => \N__56064\,
            sr => \N__56034\
        );

    \GLC_175_LC_18_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000001001"
        )
    port map (
            in0 => \N__56511\,
            in1 => \N__56432\,
            in2 => \N__56364\,
            in3 => \N__56327\,
            lcout => \INLC_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56262\,
            ce => \N__56064\,
            sr => \N__56034\
        );

    \i9544_2_lut_LC_18_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__56001\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55995\,
            lcout => \INHA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
