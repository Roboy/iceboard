-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Jan 29 2020 19:23:48

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    TX : out std_logic;
    SDA : inout std_logic;
    SCL : inout std_logic;
    RX : in std_logic;
    NEOPXL : out std_logic;
    LED : out std_logic;
    INLC : out std_logic;
    INLB : out std_logic;
    INLA : out std_logic;
    INHC : out std_logic;
    INHB : out std_logic;
    INHA : out std_logic;
    HALL3 : in std_logic;
    HALL2 : in std_logic;
    HALL1 : in std_logic;
    FAULT_N : in std_logic;
    ENCODER1_B : in std_logic;
    ENCODER1_A : in std_logic;
    ENCODER0_B : in std_logic;
    ENCODER0_A : in std_logic;
    DE : out std_logic;
    CS_MISO : in std_logic;
    CS_CLK : out std_logic;
    CS : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__5901\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3254\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2788\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2705\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2699\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2630\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2579\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2507\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2483\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal n26 : std_logic;
signal \bfn_13_21_0_\ : std_logic;
signal n25 : std_logic;
signal n2535 : std_logic;
signal n24 : std_logic;
signal n2536 : std_logic;
signal n23 : std_logic;
signal n2537 : std_logic;
signal n22 : std_logic;
signal n2538 : std_logic;
signal n21 : std_logic;
signal n2539 : std_logic;
signal n20 : std_logic;
signal n2540 : std_logic;
signal n19 : std_logic;
signal n2541 : std_logic;
signal n2542 : std_logic;
signal n18 : std_logic;
signal \bfn_13_22_0_\ : std_logic;
signal n17_adj_394 : std_logic;
signal n2543 : std_logic;
signal n16_adj_393 : std_logic;
signal n2544 : std_logic;
signal n15_adj_392 : std_logic;
signal n2545 : std_logic;
signal n14_adj_391 : std_logic;
signal n2546 : std_logic;
signal n13_adj_390 : std_logic;
signal n2547 : std_logic;
signal n12_adj_389 : std_logic;
signal n2548 : std_logic;
signal n11 : std_logic;
signal n2549 : std_logic;
signal n2550 : std_logic;
signal n10 : std_logic;
signal \bfn_13_23_0_\ : std_logic;
signal n9 : std_logic;
signal n2551 : std_logic;
signal n8_adj_388 : std_logic;
signal n2552 : std_logic;
signal n7_adj_387 : std_logic;
signal n2553 : std_logic;
signal n6 : std_logic;
signal n2554 : std_logic;
signal n2555 : std_logic;
signal n2556 : std_logic;
signal n2557 : std_logic;
signal n2558 : std_logic;
signal \bfn_13_24_0_\ : std_logic;
signal n2559 : std_logic;
signal blink_counter_21 : std_logic;
signal blink_counter_24 : std_logic;
signal blink_counter_23 : std_logic;
signal blink_counter_22 : std_logic;
signal n2730 : std_logic;
signal \n2731_cascade_\ : std_logic;
signal blink_counter_25 : std_logic;
signal \LED_c\ : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal n2478 : std_logic;
signal n2479 : std_logic;
signal n2480 : std_logic;
signal n2481 : std_logic;
signal n2482 : std_logic;
signal n2483 : std_logic;
signal n2484 : std_logic;
signal n2485 : std_logic;
signal \bfn_14_22_0_\ : std_logic;
signal n2486 : std_logic;
signal n2487 : std_logic;
signal n2488 : std_logic;
signal n2489 : std_logic;
signal n2490 : std_logic;
signal n2491 : std_logic;
signal n2492 : std_logic;
signal n2493 : std_logic;
signal \bfn_14_23_0_\ : std_logic;
signal n2494 : std_logic;
signal n2495 : std_logic;
signal n2496 : std_logic;
signal n2497 : std_logic;
signal n2498 : std_logic;
signal n2499 : std_logic;
signal n2500 : std_logic;
signal n2501 : std_logic;
signal \bfn_14_24_0_\ : std_logic;
signal n2502 : std_logic;
signal n2503 : std_logic;
signal n2504 : std_logic;
signal n2505 : std_logic;
signal n2506 : std_logic;
signal n2507 : std_logic;
signal n2508 : std_logic;
signal delay_counter_6 : std_logic;
signal delay_counter_0 : std_logic;
signal delay_counter_9 : std_logic;
signal delay_counter_4 : std_logic;
signal delay_counter_2 : std_logic;
signal delay_counter_7 : std_logic;
signal delay_counter_5 : std_logic;
signal delay_counter_3 : std_logic;
signal delay_counter_8 : std_logic;
signal delay_counter_1 : std_logic;
signal n17 : std_logic;
signal n16 : std_logic;
signal delay_counter_11 : std_logic;
signal delay_counter_10 : std_logic;
signal \n2722_cascade_\ : std_logic;
signal delay_counter_12 : std_logic;
signal delay_counter_17 : std_logic;
signal delay_counter_15 : std_logic;
signal delay_counter_14 : std_logic;
signal n8 : std_logic;
signal delay_counter_16 : std_logic;
signal delay_counter_13 : std_logic;
signal n2715 : std_logic;
signal delay_counter_18 : std_logic;
signal delay_counter_19 : std_logic;
signal \n2721_cascade_\ : std_logic;
signal delay_counter_22 : std_logic;
signal delay_counter_21 : std_logic;
signal delay_counter_23 : std_logic;
signal \n7_cascade_\ : std_logic;
signal delay_counter_20 : std_logic;
signal delay_counter_29 : std_logic;
signal delay_counter_25 : std_logic;
signal \n2695_cascade_\ : std_logic;
signal delay_counter_28 : std_logic;
signal \n13_cascade_\ : std_logic;
signal \addr_10__N_70\ : std_logic;
signal delay_counter_31 : std_logic;
signal n13 : std_logic;
signal delay_counter_26 : std_logic;
signal delay_counter_30 : std_logic;
signal delay_counter_27 : std_logic;
signal delay_counter_24 : std_logic;
signal n14 : std_logic;
signal \n2077_cascade_\ : std_logic;
signal n2077 : std_logic;
signal \n12_cascade_\ : std_logic;
signal \bfn_17_19_0_\ : std_logic;
signal \eeprom.n2516\ : std_logic;
signal \eeprom.n2517\ : std_logic;
signal \eeprom.n2518\ : std_logic;
signal \eeprom.n2519\ : std_logic;
signal \eeprom.n2520\ : std_logic;
signal \eeprom.n2521\ : std_logic;
signal \eeprom.n2522\ : std_logic;
signal \eeprom.n2523\ : std_logic;
signal \bfn_17_20_0_\ : std_logic;
signal \eeprom.n2524\ : std_logic;
signal \eeprom.n2525\ : std_logic;
signal \eeprom.n2526\ : std_logic;
signal \eeprom.n2527\ : std_logic;
signal \eeprom.n2528\ : std_logic;
signal \eeprom.n2529\ : std_logic;
signal \eeprom.n2530\ : std_logic;
signal \n6_adj_397_cascade_\ : std_logic;
signal \n2662_cascade_\ : std_logic;
signal n2668 : std_logic;
signal \eeprom.delay_counter_0\ : std_logic;
signal \eeprom.delay_counter_2\ : std_logic;
signal \eeprom.delay_counter_5\ : std_logic;
signal \eeprom.delay_counter_10\ : std_logic;
signal \eeprom.n24_cascade_\ : std_logic;
signal \eeprom.n1338_cascade_\ : std_logic;
signal \eeprom.n575\ : std_logic;
signal \eeprom.n1435\ : std_logic;
signal \eeprom.n1435_cascade_\ : std_logic;
signal \eeprom.n1503\ : std_logic;
signal \eeprom.delay_counter_6\ : std_logic;
signal \eeprom.delay_counter_12\ : std_logic;
signal \eeprom.n16\ : std_logic;
signal \n624_cascade_\ : std_logic;
signal \eeprom.delay_counter_14\ : std_logic;
signal \eeprom.delay_counter_11\ : std_logic;
signal \eeprom.delay_counter_15\ : std_logic;
signal \eeprom.delay_counter_9\ : std_logic;
signal \eeprom.delay_counter_1\ : std_logic;
signal \eeprom.delay_counter_7\ : std_logic;
signal \eeprom.n2685_cascade_\ : std_logic;
signal \eeprom.delay_counter_3\ : std_logic;
signal \eeprom.n22\ : std_logic;
signal \eeprom.delay_counter_13\ : std_logic;
signal \eeprom.delay_counter_8\ : std_logic;
signal \eeprom.delay_counter_4\ : std_logic;
signal \eeprom.n20\ : std_logic;
signal \eeprom.i2c.n6_cascade_\ : std_logic;
signal \eeprom.i2c.counter2_7__N_256_cascade_\ : std_logic;
signal \eeprom.i2c.n1384\ : std_logic;
signal \eeprom.i2c.counter2_0\ : std_logic;
signal \bfn_19_17_0_\ : std_logic;
signal \eeprom.i2c.counter2_1\ : std_logic;
signal \eeprom.i2c.n2531\ : std_logic;
signal \eeprom.i2c.counter2_2\ : std_logic;
signal \eeprom.i2c.n2532\ : std_logic;
signal \eeprom.i2c.counter2_3\ : std_logic;
signal \eeprom.i2c.n2533\ : std_logic;
signal \eeprom.i2c.n2534\ : std_logic;
signal \eeprom.i2c.counter2_4\ : std_logic;
signal \eeprom.i2c.counter2_7__N_256\ : std_logic;
signal read : std_logic;
signal state_0 : std_logic;
signal \eeprom.n1338\ : std_logic;
signal \CLK_c\ : std_logic;
signal state_1 : std_logic;
signal \eeprom.i2c.n2740_cascade_\ : std_logic;
signal \eeprom.i2c.n970\ : std_logic;
signal \eeprom.i2c.n2747_cascade_\ : std_logic;
signal \eeprom.i2c.n15_adj_381_cascade_\ : std_logic;
signal \eeprom.i2c.n2671\ : std_logic;
signal \eeprom.i2c.n2671_cascade_\ : std_logic;
signal rw : std_logic;
signal n15 : std_logic;
signal \state_7_N_269_0\ : std_logic;
signal \n15_cascade_\ : std_logic;
signal \eeprom.i2c.n37\ : std_logic;
signal n7_adj_385 : std_logic;
signal \bfn_21_14_0_\ : std_logic;
signal \eeprom.i2c.n2509\ : std_logic;
signal \eeprom.i2c.n2510\ : std_logic;
signal \eeprom.i2c.n2511\ : std_logic;
signal \eeprom.i2c.n2512\ : std_logic;
signal \eeprom.i2c.n2513\ : std_logic;
signal \eeprom.i2c.n2514\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \eeprom.i2c.n2515\ : std_logic;
signal \eeprom.i2c.n1413\ : std_logic;
signal \eeprom.i2c.n1495\ : std_logic;
signal \eeprom.i2c.n2734\ : std_logic;
signal \INVeeprom.i2c.sda_out_133C_net\ : std_logic;
signal \eeprom.enable\ : std_logic;
signal \INVeeprom.i2c.write_enable_132C_net\ : std_logic;
signal \eeprom.i2c.n2736\ : std_logic;
signal \eeprom.i2c.n2664\ : std_logic;
signal \eeprom.i2c.n39_cascade_\ : std_logic;
signal \eeprom.i2c.n952\ : std_logic;
signal \eeprom.i2c.n33_cascade_\ : std_logic;
signal \eeprom.i2c.n16\ : std_logic;
signal \eeprom.i2c.n34_cascade_\ : std_logic;
signal \eeprom.i2c.n2616\ : std_logic;
signal \eeprom.i2c.n36\ : std_logic;
signal \eeprom.i2c.n33\ : std_logic;
signal \eeprom.i2c.n36_cascade_\ : std_logic;
signal \eeprom.i2c.n1493\ : std_logic;
signal \state_7_N_285_3\ : std_logic;
signal \eeprom.i2c.n11\ : std_logic;
signal saved_addr_0 : std_logic;
signal \eeprom.i2c.n11_adj_377\ : std_logic;
signal \eeprom.i2c.n11_adj_378\ : std_logic;
signal \eeprom.i2c.counter_4\ : std_logic;
signal \eeprom.i2c.counter_6\ : std_logic;
signal \eeprom.i2c.counter_7\ : std_logic;
signal \eeprom.i2c.counter_5\ : std_logic;
signal \eeprom.i2c.counter_3\ : std_logic;
signal \eeprom.i2c.n10_adj_380_cascade_\ : std_logic;
signal \eeprom.i2c.counter_2\ : std_logic;
signal \eeprom.i2c.n2706\ : std_logic;
signal \eeprom.i2c.n2654\ : std_logic;
signal \eeprom.i2c.counter_1\ : std_logic;
signal \eeprom.i2c.n2063_cascade_\ : std_logic;
signal \eeprom.i2c.counter_0\ : std_logic;
signal \eeprom.i2c.n1358_cascade_\ : std_logic;
signal \eeprom.i2c.n2726\ : std_logic;
signal \eeprom.i2c.n876_cascade_\ : std_logic;
signal \eeprom.i2c.n2078\ : std_logic;
signal \eeprom.i2c.n11_adj_376\ : std_logic;
signal \eeprom.i2c.n21\ : std_logic;
signal \eeprom.i2c.n2714\ : std_logic;
signal \eeprom.i2c.n2741_cascade_\ : std_logic;
signal \eeprom.i2c.n10_adj_379\ : std_logic;
signal \eeprom.i2c.n2018\ : std_logic;
signal sda_enable : std_logic;
signal \eeprom.i2c.n10\ : std_logic;
signal \eeprom.i2c.sda_out\ : std_logic;
signal \eeprom.i2c.n876\ : std_logic;
signal \eeprom.i2c.n2008\ : std_logic;
signal \INVeeprom.i2c.i2c_scl_enable_124C_net\ : std_logic;
signal \eeprom.i2c.n9\ : std_logic;
signal \eeprom.state_3\ : std_logic;
signal state_0_adj_386 : std_logic;
signal \eeprom.state_1_adj_383\ : std_logic;
signal \eeprom.state_2\ : std_logic;
signal \eeprom.i2c.n11_adj_382\ : std_logic;
signal scl_enable : std_logic;
signal \eeprom.i2c.i2c_clk\ : std_logic;
signal scl_c : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CS_CLK_wire\ : std_logic;
signal \CS_wire\ : std_logic;
signal \DE_wire\ : std_logic;
signal \INHA_wire\ : std_logic;
signal \INHB_wire\ : std_logic;
signal \INHC_wire\ : std_logic;
signal \INLA_wire\ : std_logic;
signal \INLB_wire\ : std_logic;
signal \INLC_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \NEOPXL_wire\ : std_logic;
signal \TX_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    CS_CLK <= \CS_CLK_wire\;
    CS <= \CS_wire\;
    DE <= \DE_wire\;
    INHA <= \INHA_wire\;
    INHB <= \INHB_wire\;
    INHC <= \INHC_wire\;
    INLA <= \INLA_wire\;
    INLB <= \INLB_wire\;
    INLC <= \INLC_wire\;
    LED <= \LED_wire\;
    NEOPXL <= \NEOPXL_wire\;
    TX <= \TX_wire\;
    USBPU <= \USBPU_wire\;
    \CLK_wire\ <= CLK;

    \CS_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5901\,
            DIN => \N__5900\,
            DOUT => \N__5899\,
            PACKAGEPIN => \CS_CLK_wire\
        );

    \CS_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5901\,
            PADOUT => \N__5900\,
            PADIN => \N__5899\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \CS_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5892\,
            DIN => \N__5891\,
            DOUT => \N__5890\,
            PACKAGEPIN => \CS_wire\
        );

    \CS_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5892\,
            PADOUT => \N__5891\,
            PADIN => \N__5890\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \DE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5883\,
            DIN => \N__5882\,
            DOUT => \N__5881\,
            PACKAGEPIN => \DE_wire\
        );

    \DE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5883\,
            PADOUT => \N__5882\,
            PADIN => \N__5881\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHA_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5874\,
            DIN => \N__5873\,
            DOUT => \N__5872\,
            PACKAGEPIN => \INHA_wire\
        );

    \INHA_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5874\,
            PADOUT => \N__5873\,
            PADIN => \N__5872\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHB_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5865\,
            DIN => \N__5864\,
            DOUT => \N__5863\,
            PACKAGEPIN => \INHB_wire\
        );

    \INHB_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5865\,
            PADOUT => \N__5864\,
            PADIN => \N__5863\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5856\,
            DIN => \N__5855\,
            DOUT => \N__5854\,
            PACKAGEPIN => \INHC_wire\
        );

    \INHC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5856\,
            PADOUT => \N__5855\,
            PADIN => \N__5854\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLA_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5847\,
            DIN => \N__5846\,
            DOUT => \N__5845\,
            PACKAGEPIN => \INLA_wire\
        );

    \INLA_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5847\,
            PADOUT => \N__5846\,
            PADIN => \N__5845\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLB_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5838\,
            DIN => \N__5837\,
            DOUT => \N__5836\,
            PACKAGEPIN => \INLB_wire\
        );

    \INLB_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5838\,
            PADOUT => \N__5837\,
            PADIN => \N__5836\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5829\,
            DIN => \N__5828\,
            DOUT => \N__5827\,
            PACKAGEPIN => \INLC_wire\
        );

    \INLC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5829\,
            PADOUT => \N__5828\,
            PADIN => \N__5827\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5820\,
            DIN => \N__5819\,
            DOUT => \N__5818\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5820\,
            PADOUT => \N__5819\,
            PADIN => \N__5818\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__2723\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \NEOPXL_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5811\,
            DIN => \N__5810\,
            DOUT => \N__5809\,
            PACKAGEPIN => \NEOPXL_wire\
        );

    \NEOPXL_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5811\,
            PADOUT => \N__5810\,
            PADIN => \N__5809\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \TX_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5802\,
            DIN => \N__5801\,
            DOUT => \N__5800\,
            PACKAGEPIN => \TX_wire\
        );

    \TX_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5802\,
            PADOUT => \N__5801\,
            PADIN => \N__5800\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5793\,
            DIN => \N__5792\,
            DOUT => \N__5791\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5793\,
            PADOUT => \N__5792\,
            PADIN => \N__5791\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \scl_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__5784\,
            DIN => \N__5783\,
            DOUT => \N__5782\,
            PACKAGEPIN => SCL
        );

    \scl_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5784\,
            PADOUT => \N__5783\,
            PADIN => \N__5782\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__4859\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__5000\
        );

    \sda_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__5775\,
            DIN => \N__5774\,
            DOUT => \N__5773\,
            PACKAGEPIN => SDA
        );

    \sda_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5775\,
            PADOUT => \N__5774\,
            PADIN => \N__5773\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__4493\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__5717\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5766\,
            DIN => \N__5765\,
            DOUT => \N__5764\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5766\,
            PADOUT => \N__5765\,
            PADIN => \N__5764\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__1302\ : InMux
    port map (
            O => \N__5747\,
            I => \N__5743\
        );

    \I__1301\ : InMux
    port map (
            O => \N__5746\,
            I => \N__5740\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__5743\,
            I => \N__5737\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__5740\,
            I => \eeprom.i2c.n10_adj_379\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__5737\,
            I => \eeprom.i2c.n10_adj_379\
        );

    \I__1297\ : InMux
    port map (
            O => \N__5732\,
            I => \N__5728\
        );

    \I__1296\ : InMux
    port map (
            O => \N__5731\,
            I => \N__5725\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__5728\,
            I => \N__5720\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__5725\,
            I => \N__5720\
        );

    \I__1293\ : Odrv4
    port map (
            O => \N__5720\,
            I => \eeprom.i2c.n2018\
        );

    \I__1292\ : IoInMux
    port map (
            O => \N__5717\,
            I => \N__5714\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__5714\,
            I => \N__5710\
        );

    \I__1290\ : InMux
    port map (
            O => \N__5713\,
            I => \N__5707\
        );

    \I__1289\ : Span12Mux_s11_h
    port map (
            O => \N__5710\,
            I => \N__5702\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__5707\,
            I => \N__5699\
        );

    \I__1287\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5696\
        );

    \I__1286\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5693\
        );

    \I__1285\ : Odrv12
    port map (
            O => \N__5702\,
            I => sda_enable
        );

    \I__1284\ : Odrv4
    port map (
            O => \N__5699\,
            I => sda_enable
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__5696\,
            I => sda_enable
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__5693\,
            I => sda_enable
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__5684\,
            I => \N__5679\
        );

    \I__1280\ : InMux
    port map (
            O => \N__5683\,
            I => \N__5676\
        );

    \I__1279\ : InMux
    port map (
            O => \N__5682\,
            I => \N__5673\
        );

    \I__1278\ : InMux
    port map (
            O => \N__5679\,
            I => \N__5670\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__5676\,
            I => \N__5667\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__5673\,
            I => \N__5664\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__5670\,
            I => \eeprom.i2c.n10\
        );

    \I__1274\ : Odrv4
    port map (
            O => \N__5667\,
            I => \eeprom.i2c.n10\
        );

    \I__1273\ : Odrv4
    port map (
            O => \N__5664\,
            I => \eeprom.i2c.n10\
        );

    \I__1272\ : InMux
    port map (
            O => \N__5657\,
            I => \N__5654\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__5654\,
            I => \N__5651\
        );

    \I__1270\ : Span4Mux_h
    port map (
            O => \N__5651\,
            I => \N__5646\
        );

    \I__1269\ : InMux
    port map (
            O => \N__5650\,
            I => \N__5643\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5649\,
            I => \N__5640\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__5646\,
            I => \eeprom.i2c.sda_out\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__5643\,
            I => \eeprom.i2c.sda_out\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__5640\,
            I => \eeprom.i2c.sda_out\
        );

    \I__1264\ : CascadeMux
    port map (
            O => \N__5633\,
            I => \N__5627\
        );

    \I__1263\ : CEMux
    port map (
            O => \N__5632\,
            I => \N__5622\
        );

    \I__1262\ : CEMux
    port map (
            O => \N__5631\,
            I => \N__5619\
        );

    \I__1261\ : CEMux
    port map (
            O => \N__5630\,
            I => \N__5616\
        );

    \I__1260\ : InMux
    port map (
            O => \N__5627\,
            I => \N__5613\
        );

    \I__1259\ : InMux
    port map (
            O => \N__5626\,
            I => \N__5608\
        );

    \I__1258\ : InMux
    port map (
            O => \N__5625\,
            I => \N__5608\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__5622\,
            I => \eeprom.i2c.n876\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__5619\,
            I => \eeprom.i2c.n876\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__5616\,
            I => \eeprom.i2c.n876\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__5613\,
            I => \eeprom.i2c.n876\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__5608\,
            I => \eeprom.i2c.n876\
        );

    \I__1252\ : SRMux
    port map (
            O => \N__5597\,
            I => \N__5594\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__5594\,
            I => \N__5591\
        );

    \I__1250\ : Odrv4
    port map (
            O => \N__5591\,
            I => \eeprom.i2c.n2008\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__5588\,
            I => \N__5585\
        );

    \I__1248\ : InMux
    port map (
            O => \N__5585\,
            I => \N__5582\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__5582\,
            I => \eeprom.i2c.n9\
        );

    \I__1246\ : InMux
    port map (
            O => \N__5579\,
            I => \N__5575\
        );

    \I__1245\ : InMux
    port map (
            O => \N__5578\,
            I => \N__5570\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__5575\,
            I => \N__5559\
        );

    \I__1243\ : InMux
    port map (
            O => \N__5574\,
            I => \N__5556\
        );

    \I__1242\ : InMux
    port map (
            O => \N__5573\,
            I => \N__5553\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__5570\,
            I => \N__5550\
        );

    \I__1240\ : InMux
    port map (
            O => \N__5569\,
            I => \N__5547\
        );

    \I__1239\ : InMux
    port map (
            O => \N__5568\,
            I => \N__5539\
        );

    \I__1238\ : InMux
    port map (
            O => \N__5567\,
            I => \N__5539\
        );

    \I__1237\ : InMux
    port map (
            O => \N__5566\,
            I => \N__5539\
        );

    \I__1236\ : InMux
    port map (
            O => \N__5565\,
            I => \N__5536\
        );

    \I__1235\ : InMux
    port map (
            O => \N__5564\,
            I => \N__5532\
        );

    \I__1234\ : CascadeMux
    port map (
            O => \N__5563\,
            I => \N__5527\
        );

    \I__1233\ : InMux
    port map (
            O => \N__5562\,
            I => \N__5521\
        );

    \I__1232\ : Span4Mux_h
    port map (
            O => \N__5559\,
            I => \N__5514\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__5556\,
            I => \N__5514\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__5553\,
            I => \N__5514\
        );

    \I__1229\ : Span4Mux_h
    port map (
            O => \N__5550\,
            I => \N__5509\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__5547\,
            I => \N__5509\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5546\,
            I => \N__5506\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__5539\,
            I => \N__5501\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__5536\,
            I => \N__5501\
        );

    \I__1224\ : InMux
    port map (
            O => \N__5535\,
            I => \N__5493\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__5532\,
            I => \N__5490\
        );

    \I__1222\ : InMux
    port map (
            O => \N__5531\,
            I => \N__5483\
        );

    \I__1221\ : InMux
    port map (
            O => \N__5530\,
            I => \N__5483\
        );

    \I__1220\ : InMux
    port map (
            O => \N__5527\,
            I => \N__5483\
        );

    \I__1219\ : InMux
    port map (
            O => \N__5526\,
            I => \N__5476\
        );

    \I__1218\ : InMux
    port map (
            O => \N__5525\,
            I => \N__5476\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5476\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__5521\,
            I => \N__5473\
        );

    \I__1215\ : Span4Mux_v
    port map (
            O => \N__5514\,
            I => \N__5466\
        );

    \I__1214\ : Span4Mux_v
    port map (
            O => \N__5509\,
            I => \N__5466\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__5506\,
            I => \N__5466\
        );

    \I__1212\ : Span4Mux_h
    port map (
            O => \N__5501\,
            I => \N__5463\
        );

    \I__1211\ : InMux
    port map (
            O => \N__5500\,
            I => \N__5456\
        );

    \I__1210\ : InMux
    port map (
            O => \N__5499\,
            I => \N__5456\
        );

    \I__1209\ : InMux
    port map (
            O => \N__5498\,
            I => \N__5456\
        );

    \I__1208\ : InMux
    port map (
            O => \N__5497\,
            I => \N__5451\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5496\,
            I => \N__5451\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__5493\,
            I => \N__5448\
        );

    \I__1205\ : Odrv4
    port map (
            O => \N__5490\,
            I => \eeprom.state_3\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__5483\,
            I => \eeprom.state_3\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__5476\,
            I => \eeprom.state_3\
        );

    \I__1202\ : Odrv12
    port map (
            O => \N__5473\,
            I => \eeprom.state_3\
        );

    \I__1201\ : Odrv4
    port map (
            O => \N__5466\,
            I => \eeprom.state_3\
        );

    \I__1200\ : Odrv4
    port map (
            O => \N__5463\,
            I => \eeprom.state_3\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__5456\,
            I => \eeprom.state_3\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__5451\,
            I => \eeprom.state_3\
        );

    \I__1197\ : Odrv4
    port map (
            O => \N__5448\,
            I => \eeprom.state_3\
        );

    \I__1196\ : InMux
    port map (
            O => \N__5429\,
            I => \N__5425\
        );

    \I__1195\ : CascadeMux
    port map (
            O => \N__5428\,
            I => \N__5416\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__5425\,
            I => \N__5411\
        );

    \I__1193\ : InMux
    port map (
            O => \N__5424\,
            I => \N__5408\
        );

    \I__1192\ : InMux
    port map (
            O => \N__5423\,
            I => \N__5405\
        );

    \I__1191\ : InMux
    port map (
            O => \N__5422\,
            I => \N__5402\
        );

    \I__1190\ : InMux
    port map (
            O => \N__5421\,
            I => \N__5392\
        );

    \I__1189\ : InMux
    port map (
            O => \N__5420\,
            I => \N__5389\
        );

    \I__1188\ : InMux
    port map (
            O => \N__5419\,
            I => \N__5384\
        );

    \I__1187\ : InMux
    port map (
            O => \N__5416\,
            I => \N__5384\
        );

    \I__1186\ : InMux
    port map (
            O => \N__5415\,
            I => \N__5381\
        );

    \I__1185\ : InMux
    port map (
            O => \N__5414\,
            I => \N__5378\
        );

    \I__1184\ : Span4Mux_v
    port map (
            O => \N__5411\,
            I => \N__5373\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__5408\,
            I => \N__5373\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__5405\,
            I => \N__5368\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__5402\,
            I => \N__5368\
        );

    \I__1180\ : CascadeMux
    port map (
            O => \N__5401\,
            I => \N__5361\
        );

    \I__1179\ : CascadeMux
    port map (
            O => \N__5400\,
            I => \N__5357\
        );

    \I__1178\ : InMux
    port map (
            O => \N__5399\,
            I => \N__5353\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5398\,
            I => \N__5350\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5397\,
            I => \N__5347\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5396\,
            I => \N__5342\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5342\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__5392\,
            I => \N__5335\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__5389\,
            I => \N__5335\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__5384\,
            I => \N__5335\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__5381\,
            I => \N__5328\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__5378\,
            I => \N__5328\
        );

    \I__1168\ : Span4Mux_h
    port map (
            O => \N__5373\,
            I => \N__5328\
        );

    \I__1167\ : Span4Mux_h
    port map (
            O => \N__5368\,
            I => \N__5325\
        );

    \I__1166\ : InMux
    port map (
            O => \N__5367\,
            I => \N__5316\
        );

    \I__1165\ : InMux
    port map (
            O => \N__5366\,
            I => \N__5316\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5365\,
            I => \N__5316\
        );

    \I__1163\ : InMux
    port map (
            O => \N__5364\,
            I => \N__5316\
        );

    \I__1162\ : InMux
    port map (
            O => \N__5361\,
            I => \N__5313\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5360\,
            I => \N__5310\
        );

    \I__1160\ : InMux
    port map (
            O => \N__5357\,
            I => \N__5305\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5356\,
            I => \N__5305\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5353\,
            I => state_0_adj_386
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__5350\,
            I => state_0_adj_386
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__5347\,
            I => state_0_adj_386
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__5342\,
            I => state_0_adj_386
        );

    \I__1154\ : Odrv4
    port map (
            O => \N__5335\,
            I => state_0_adj_386
        );

    \I__1153\ : Odrv4
    port map (
            O => \N__5328\,
            I => state_0_adj_386
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__5325\,
            I => state_0_adj_386
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__5316\,
            I => state_0_adj_386
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__5313\,
            I => state_0_adj_386
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__5310\,
            I => state_0_adj_386
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__5305\,
            I => state_0_adj_386
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__5282\,
            I => \N__5274\
        );

    \I__1146\ : CascadeMux
    port map (
            O => \N__5281\,
            I => \N__5271\
        );

    \I__1145\ : CascadeMux
    port map (
            O => \N__5280\,
            I => \N__5267\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__5279\,
            I => \N__5263\
        );

    \I__1143\ : InMux
    port map (
            O => \N__5278\,
            I => \N__5254\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5277\,
            I => \N__5249\
        );

    \I__1141\ : InMux
    port map (
            O => \N__5274\,
            I => \N__5249\
        );

    \I__1140\ : InMux
    port map (
            O => \N__5271\,
            I => \N__5246\
        );

    \I__1139\ : InMux
    port map (
            O => \N__5270\,
            I => \N__5241\
        );

    \I__1138\ : InMux
    port map (
            O => \N__5267\,
            I => \N__5241\
        );

    \I__1137\ : InMux
    port map (
            O => \N__5266\,
            I => \N__5238\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5263\,
            I => \N__5233\
        );

    \I__1135\ : CascadeMux
    port map (
            O => \N__5262\,
            I => \N__5230\
        );

    \I__1134\ : InMux
    port map (
            O => \N__5261\,
            I => \N__5227\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5260\,
            I => \N__5222\
        );

    \I__1132\ : InMux
    port map (
            O => \N__5259\,
            I => \N__5222\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5258\,
            I => \N__5217\
        );

    \I__1130\ : InMux
    port map (
            O => \N__5257\,
            I => \N__5217\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__5254\,
            I => \N__5214\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__5249\,
            I => \N__5211\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__5246\,
            I => \N__5204\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__5241\,
            I => \N__5204\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__5238\,
            I => \N__5204\
        );

    \I__1124\ : CascadeMux
    port map (
            O => \N__5237\,
            I => \N__5201\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__5236\,
            I => \N__5196\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__5233\,
            I => \N__5189\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5230\,
            I => \N__5186\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__5227\,
            I => \N__5179\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__5222\,
            I => \N__5179\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__5217\,
            I => \N__5179\
        );

    \I__1117\ : Span4Mux_v
    port map (
            O => \N__5214\,
            I => \N__5172\
        );

    \I__1116\ : Span4Mux_v
    port map (
            O => \N__5211\,
            I => \N__5172\
        );

    \I__1115\ : Span4Mux_v
    port map (
            O => \N__5204\,
            I => \N__5172\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5201\,
            I => \N__5169\
        );

    \I__1113\ : InMux
    port map (
            O => \N__5200\,
            I => \N__5162\
        );

    \I__1112\ : InMux
    port map (
            O => \N__5199\,
            I => \N__5162\
        );

    \I__1111\ : InMux
    port map (
            O => \N__5196\,
            I => \N__5162\
        );

    \I__1110\ : InMux
    port map (
            O => \N__5195\,
            I => \N__5159\
        );

    \I__1109\ : InMux
    port map (
            O => \N__5194\,
            I => \N__5152\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5193\,
            I => \N__5152\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5192\,
            I => \N__5152\
        );

    \I__1106\ : Odrv4
    port map (
            O => \N__5189\,
            I => \eeprom.state_1_adj_383\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__5186\,
            I => \eeprom.state_1_adj_383\
        );

    \I__1104\ : Odrv4
    port map (
            O => \N__5179\,
            I => \eeprom.state_1_adj_383\
        );

    \I__1103\ : Odrv4
    port map (
            O => \N__5172\,
            I => \eeprom.state_1_adj_383\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5169\,
            I => \eeprom.state_1_adj_383\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__5162\,
            I => \eeprom.state_1_adj_383\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__5159\,
            I => \eeprom.state_1_adj_383\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__5152\,
            I => \eeprom.state_1_adj_383\
        );

    \I__1098\ : InMux
    port map (
            O => \N__5135\,
            I => \N__5120\
        );

    \I__1097\ : InMux
    port map (
            O => \N__5134\,
            I => \N__5114\
        );

    \I__1096\ : InMux
    port map (
            O => \N__5133\,
            I => \N__5114\
        );

    \I__1095\ : InMux
    port map (
            O => \N__5132\,
            I => \N__5111\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5131\,
            I => \N__5108\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5130\,
            I => \N__5101\
        );

    \I__1092\ : InMux
    port map (
            O => \N__5129\,
            I => \N__5101\
        );

    \I__1091\ : InMux
    port map (
            O => \N__5128\,
            I => \N__5101\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5127\,
            I => \N__5098\
        );

    \I__1089\ : InMux
    port map (
            O => \N__5126\,
            I => \N__5094\
        );

    \I__1088\ : InMux
    port map (
            O => \N__5125\,
            I => \N__5087\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5124\,
            I => \N__5087\
        );

    \I__1086\ : InMux
    port map (
            O => \N__5123\,
            I => \N__5087\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__5120\,
            I => \N__5083\
        );

    \I__1084\ : InMux
    port map (
            O => \N__5119\,
            I => \N__5080\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__5114\,
            I => \N__5071\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__5111\,
            I => \N__5071\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__5108\,
            I => \N__5071\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__5101\,
            I => \N__5071\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__5098\,
            I => \N__5061\
        );

    \I__1078\ : InMux
    port map (
            O => \N__5097\,
            I => \N__5058\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__5094\,
            I => \N__5055\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5087\,
            I => \N__5052\
        );

    \I__1075\ : InMux
    port map (
            O => \N__5086\,
            I => \N__5049\
        );

    \I__1074\ : Span4Mux_v
    port map (
            O => \N__5083\,
            I => \N__5042\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__5080\,
            I => \N__5042\
        );

    \I__1072\ : Span4Mux_v
    port map (
            O => \N__5071\,
            I => \N__5042\
        );

    \I__1071\ : InMux
    port map (
            O => \N__5070\,
            I => \N__5035\
        );

    \I__1070\ : InMux
    port map (
            O => \N__5069\,
            I => \N__5035\
        );

    \I__1069\ : InMux
    port map (
            O => \N__5068\,
            I => \N__5035\
        );

    \I__1068\ : InMux
    port map (
            O => \N__5067\,
            I => \N__5026\
        );

    \I__1067\ : InMux
    port map (
            O => \N__5066\,
            I => \N__5026\
        );

    \I__1066\ : InMux
    port map (
            O => \N__5065\,
            I => \N__5026\
        );

    \I__1065\ : InMux
    port map (
            O => \N__5064\,
            I => \N__5026\
        );

    \I__1064\ : Odrv4
    port map (
            O => \N__5061\,
            I => \eeprom.state_2\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__5058\,
            I => \eeprom.state_2\
        );

    \I__1062\ : Odrv4
    port map (
            O => \N__5055\,
            I => \eeprom.state_2\
        );

    \I__1061\ : Odrv4
    port map (
            O => \N__5052\,
            I => \eeprom.state_2\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__5049\,
            I => \eeprom.state_2\
        );

    \I__1059\ : Odrv4
    port map (
            O => \N__5042\,
            I => \eeprom.state_2\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__5035\,
            I => \eeprom.state_2\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__5026\,
            I => \eeprom.state_2\
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__5009\,
            I => \N__5006\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5006\,
            I => \N__5003\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__5003\,
            I => \eeprom.i2c.n11_adj_382\
        );

    \I__1053\ : IoInMux
    port map (
            O => \N__5000\,
            I => \N__4997\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__4997\,
            I => \N__4994\
        );

    \I__1051\ : Span4Mux_s2_h
    port map (
            O => \N__4994\,
            I => \N__4991\
        );

    \I__1050\ : Span4Mux_v
    port map (
            O => \N__4991\,
            I => \N__4987\
        );

    \I__1049\ : InMux
    port map (
            O => \N__4990\,
            I => \N__4984\
        );

    \I__1048\ : Sp12to4
    port map (
            O => \N__4987\,
            I => \N__4979\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__4984\,
            I => \N__4979\
        );

    \I__1046\ : Odrv12
    port map (
            O => \N__4979\,
            I => scl_enable
        );

    \I__1045\ : ClkMux
    port map (
            O => \N__4976\,
            I => \N__4969\
        );

    \I__1044\ : ClkMux
    port map (
            O => \N__4975\,
            I => \N__4966\
        );

    \I__1043\ : ClkMux
    port map (
            O => \N__4974\,
            I => \N__4963\
        );

    \I__1042\ : ClkMux
    port map (
            O => \N__4973\,
            I => \N__4960\
        );

    \I__1041\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4957\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__4969\,
            I => \N__4950\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__4966\,
            I => \N__4947\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__4963\,
            I => \N__4941\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__4960\,
            I => \N__4941\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__4957\,
            I => \N__4938\
        );

    \I__1035\ : ClkMux
    port map (
            O => \N__4956\,
            I => \N__4935\
        );

    \I__1034\ : ClkMux
    port map (
            O => \N__4955\,
            I => \N__4932\
        );

    \I__1033\ : ClkMux
    port map (
            O => \N__4954\,
            I => \N__4929\
        );

    \I__1032\ : ClkMux
    port map (
            O => \N__4953\,
            I => \N__4926\
        );

    \I__1031\ : Span4Mux_h
    port map (
            O => \N__4950\,
            I => \N__4921\
        );

    \I__1030\ : Span4Mux_v
    port map (
            O => \N__4947\,
            I => \N__4921\
        );

    \I__1029\ : ClkMux
    port map (
            O => \N__4946\,
            I => \N__4918\
        );

    \I__1028\ : Span4Mux_v
    port map (
            O => \N__4941\,
            I => \N__4915\
        );

    \I__1027\ : Span4Mux_v
    port map (
            O => \N__4938\,
            I => \N__4912\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__4935\,
            I => \N__4907\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__4932\,
            I => \N__4907\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__4929\,
            I => \N__4904\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__4926\,
            I => \N__4897\
        );

    \I__1022\ : Span4Mux_h
    port map (
            O => \N__4921\,
            I => \N__4897\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__4918\,
            I => \N__4897\
        );

    \I__1020\ : Span4Mux_h
    port map (
            O => \N__4915\,
            I => \N__4891\
        );

    \I__1019\ : Span4Mux_h
    port map (
            O => \N__4912\,
            I => \N__4886\
        );

    \I__1018\ : Span4Mux_v
    port map (
            O => \N__4907\,
            I => \N__4886\
        );

    \I__1017\ : Span4Mux_v
    port map (
            O => \N__4904\,
            I => \N__4883\
        );

    \I__1016\ : Span4Mux_v
    port map (
            O => \N__4897\,
            I => \N__4880\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4896\,
            I => \N__4877\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4895\,
            I => \N__4872\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4894\,
            I => \N__4872\
        );

    \I__1012\ : Odrv4
    port map (
            O => \N__4891\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1011\ : Odrv4
    port map (
            O => \N__4886\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1010\ : Odrv4
    port map (
            O => \N__4883\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1009\ : Odrv4
    port map (
            O => \N__4880\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__4877\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__4872\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1006\ : IoInMux
    port map (
            O => \N__4859\,
            I => \N__4856\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__4856\,
            I => \N__4853\
        );

    \I__1004\ : Span4Mux_s3_h
    port map (
            O => \N__4853\,
            I => \N__4850\
        );

    \I__1003\ : Span4Mux_v
    port map (
            O => \N__4850\,
            I => \N__4847\
        );

    \I__1002\ : Odrv4
    port map (
            O => \N__4847\,
            I => scl_c
        );

    \I__1001\ : InMux
    port map (
            O => \N__4844\,
            I => \N__4841\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4841\,
            I => \N__4837\
        );

    \I__999\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4834\
        );

    \I__998\ : Odrv12
    port map (
            O => \N__4837\,
            I => \eeprom.i2c.n2654\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__4834\,
            I => \eeprom.i2c.n2654\
        );

    \I__996\ : InMux
    port map (
            O => \N__4829\,
            I => \N__4826\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__4826\,
            I => \N__4822\
        );

    \I__994\ : InMux
    port map (
            O => \N__4825\,
            I => \N__4817\
        );

    \I__993\ : Span4Mux_h
    port map (
            O => \N__4822\,
            I => \N__4814\
        );

    \I__992\ : InMux
    port map (
            O => \N__4821\,
            I => \N__4809\
        );

    \I__991\ : InMux
    port map (
            O => \N__4820\,
            I => \N__4809\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__4817\,
            I => \eeprom.i2c.counter_1\
        );

    \I__989\ : Odrv4
    port map (
            O => \N__4814\,
            I => \eeprom.i2c.counter_1\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__4809\,
            I => \eeprom.i2c.counter_1\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__4802\,
            I => \eeprom.i2c.n2063_cascade_\
        );

    \I__986\ : InMux
    port map (
            O => \N__4799\,
            I => \N__4796\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__4796\,
            I => \N__4792\
        );

    \I__984\ : InMux
    port map (
            O => \N__4795\,
            I => \N__4786\
        );

    \I__983\ : Span4Mux_h
    port map (
            O => \N__4792\,
            I => \N__4783\
        );

    \I__982\ : InMux
    port map (
            O => \N__4791\,
            I => \N__4776\
        );

    \I__981\ : InMux
    port map (
            O => \N__4790\,
            I => \N__4776\
        );

    \I__980\ : InMux
    port map (
            O => \N__4789\,
            I => \N__4776\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__4786\,
            I => \eeprom.i2c.counter_0\
        );

    \I__978\ : Odrv4
    port map (
            O => \N__4783\,
            I => \eeprom.i2c.counter_0\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__4776\,
            I => \eeprom.i2c.counter_0\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__4769\,
            I => \eeprom.i2c.n1358_cascade_\
        );

    \I__975\ : InMux
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__4763\,
            I => \N__4760\
        );

    \I__973\ : Odrv4
    port map (
            O => \N__4760\,
            I => \eeprom.i2c.n2726\
        );

    \I__972\ : CascadeMux
    port map (
            O => \N__4757\,
            I => \eeprom.i2c.n876_cascade_\
        );

    \I__971\ : SRMux
    port map (
            O => \N__4754\,
            I => \N__4751\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__4751\,
            I => \eeprom.i2c.n2078\
        );

    \I__969\ : InMux
    port map (
            O => \N__4748\,
            I => \N__4739\
        );

    \I__968\ : InMux
    port map (
            O => \N__4747\,
            I => \N__4739\
        );

    \I__967\ : InMux
    port map (
            O => \N__4746\,
            I => \N__4739\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4739\,
            I => \eeprom.i2c.n11_adj_376\
        );

    \I__965\ : InMux
    port map (
            O => \N__4736\,
            I => \N__4733\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__4733\,
            I => \eeprom.i2c.n21\
        );

    \I__963\ : InMux
    port map (
            O => \N__4730\,
            I => \N__4727\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__4727\,
            I => \N__4724\
        );

    \I__961\ : Odrv12
    port map (
            O => \N__4724\,
            I => \eeprom.i2c.n2714\
        );

    \I__960\ : CascadeMux
    port map (
            O => \N__4721\,
            I => \eeprom.i2c.n2741_cascade_\
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__4718\,
            I => \N__4715\
        );

    \I__958\ : InMux
    port map (
            O => \N__4715\,
            I => \N__4710\
        );

    \I__957\ : InMux
    port map (
            O => \N__4714\,
            I => \N__4707\
        );

    \I__956\ : InMux
    port map (
            O => \N__4713\,
            I => \N__4704\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4710\,
            I => \eeprom.i2c.n11_adj_377\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4707\,
            I => \eeprom.i2c.n11_adj_377\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4704\,
            I => \eeprom.i2c.n11_adj_377\
        );

    \I__952\ : InMux
    port map (
            O => \N__4697\,
            I => \N__4694\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__4694\,
            I => \N__4691\
        );

    \I__950\ : Odrv4
    port map (
            O => \N__4691\,
            I => \eeprom.i2c.n11_adj_378\
        );

    \I__949\ : CascadeMux
    port map (
            O => \N__4688\,
            I => \N__4684\
        );

    \I__948\ : InMux
    port map (
            O => \N__4687\,
            I => \N__4681\
        );

    \I__947\ : InMux
    port map (
            O => \N__4684\,
            I => \N__4678\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4681\,
            I => \N__4675\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4678\,
            I => \eeprom.i2c.counter_4\
        );

    \I__944\ : Odrv4
    port map (
            O => \N__4675\,
            I => \eeprom.i2c.counter_4\
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__4670\,
            I => \N__4666\
        );

    \I__942\ : InMux
    port map (
            O => \N__4669\,
            I => \N__4663\
        );

    \I__941\ : InMux
    port map (
            O => \N__4666\,
            I => \N__4660\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__4663\,
            I => \N__4657\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4660\,
            I => \eeprom.i2c.counter_6\
        );

    \I__938\ : Odrv12
    port map (
            O => \N__4657\,
            I => \eeprom.i2c.counter_6\
        );

    \I__937\ : CascadeMux
    port map (
            O => \N__4652\,
            I => \N__4649\
        );

    \I__936\ : InMux
    port map (
            O => \N__4649\,
            I => \N__4645\
        );

    \I__935\ : InMux
    port map (
            O => \N__4648\,
            I => \N__4642\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__4645\,
            I => \N__4639\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4642\,
            I => \eeprom.i2c.counter_7\
        );

    \I__932\ : Odrv4
    port map (
            O => \N__4639\,
            I => \eeprom.i2c.counter_7\
        );

    \I__931\ : InMux
    port map (
            O => \N__4634\,
            I => \N__4630\
        );

    \I__930\ : InMux
    port map (
            O => \N__4633\,
            I => \N__4627\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__4630\,
            I => \N__4624\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__4627\,
            I => \eeprom.i2c.counter_5\
        );

    \I__927\ : Odrv4
    port map (
            O => \N__4624\,
            I => \eeprom.i2c.counter_5\
        );

    \I__926\ : InMux
    port map (
            O => \N__4619\,
            I => \N__4615\
        );

    \I__925\ : InMux
    port map (
            O => \N__4618\,
            I => \N__4612\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__4615\,
            I => \N__4609\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__4612\,
            I => \eeprom.i2c.counter_3\
        );

    \I__922\ : Odrv4
    port map (
            O => \N__4609\,
            I => \eeprom.i2c.counter_3\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__4604\,
            I => \eeprom.i2c.n10_adj_380_cascade_\
        );

    \I__920\ : CascadeMux
    port map (
            O => \N__4601\,
            I => \N__4597\
        );

    \I__919\ : InMux
    port map (
            O => \N__4600\,
            I => \N__4593\
        );

    \I__918\ : InMux
    port map (
            O => \N__4597\,
            I => \N__4590\
        );

    \I__917\ : InMux
    port map (
            O => \N__4596\,
            I => \N__4587\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4593\,
            I => \N__4584\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__4590\,
            I => \eeprom.i2c.counter_2\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4587\,
            I => \eeprom.i2c.counter_2\
        );

    \I__913\ : Odrv4
    port map (
            O => \N__4584\,
            I => \eeprom.i2c.counter_2\
        );

    \I__912\ : SRMux
    port map (
            O => \N__4577\,
            I => \N__4574\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__4574\,
            I => \eeprom.i2c.n2706\
        );

    \I__910\ : CascadeMux
    port map (
            O => \N__4571\,
            I => \eeprom.i2c.n39_cascade_\
        );

    \I__909\ : CEMux
    port map (
            O => \N__4568\,
            I => \N__4565\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4565\,
            I => \N__4562\
        );

    \I__907\ : Span4Mux_h
    port map (
            O => \N__4562\,
            I => \N__4559\
        );

    \I__906\ : Odrv4
    port map (
            O => \N__4559\,
            I => \eeprom.i2c.n952\
        );

    \I__905\ : CascadeMux
    port map (
            O => \N__4556\,
            I => \eeprom.i2c.n33_cascade_\
        );

    \I__904\ : InMux
    port map (
            O => \N__4553\,
            I => \N__4550\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4550\,
            I => \eeprom.i2c.n16\
        );

    \I__902\ : CascadeMux
    port map (
            O => \N__4547\,
            I => \eeprom.i2c.n34_cascade_\
        );

    \I__901\ : CEMux
    port map (
            O => \N__4544\,
            I => \N__4541\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4541\,
            I => \N__4538\
        );

    \I__899\ : Odrv4
    port map (
            O => \N__4538\,
            I => \eeprom.i2c.n2616\
        );

    \I__898\ : InMux
    port map (
            O => \N__4535\,
            I => \N__4532\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__4532\,
            I => \N__4527\
        );

    \I__896\ : InMux
    port map (
            O => \N__4531\,
            I => \N__4522\
        );

    \I__895\ : InMux
    port map (
            O => \N__4530\,
            I => \N__4522\
        );

    \I__894\ : Odrv4
    port map (
            O => \N__4527\,
            I => \eeprom.i2c.n36\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4522\,
            I => \eeprom.i2c.n36\
        );

    \I__892\ : InMux
    port map (
            O => \N__4517\,
            I => \N__4511\
        );

    \I__891\ : InMux
    port map (
            O => \N__4516\,
            I => \N__4511\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__4511\,
            I => \eeprom.i2c.n33\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__4508\,
            I => \eeprom.i2c.n36_cascade_\
        );

    \I__888\ : SRMux
    port map (
            O => \N__4505\,
            I => \N__4502\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__4502\,
            I => \N__4499\
        );

    \I__886\ : Span4Mux_h
    port map (
            O => \N__4499\,
            I => \N__4496\
        );

    \I__885\ : Odrv4
    port map (
            O => \N__4496\,
            I => \eeprom.i2c.n1493\
        );

    \I__884\ : IoInMux
    port map (
            O => \N__4493\,
            I => \N__4490\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__4490\,
            I => \N__4487\
        );

    \I__882\ : Span12Mux_s6_h
    port map (
            O => \N__4487\,
            I => \N__4483\
        );

    \I__881\ : InMux
    port map (
            O => \N__4486\,
            I => \N__4480\
        );

    \I__880\ : Span12Mux_v
    port map (
            O => \N__4483\,
            I => \N__4476\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__4480\,
            I => \N__4473\
        );

    \I__878\ : InMux
    port map (
            O => \N__4479\,
            I => \N__4470\
        );

    \I__877\ : Odrv12
    port map (
            O => \N__4476\,
            I => \state_7_N_285_3\
        );

    \I__876\ : Odrv4
    port map (
            O => \N__4473\,
            I => \state_7_N_285_3\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4470\,
            I => \state_7_N_285_3\
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__4463\,
            I => \N__4460\
        );

    \I__873\ : InMux
    port map (
            O => \N__4460\,
            I => \N__4457\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4457\,
            I => \N__4454\
        );

    \I__871\ : Odrv12
    port map (
            O => \N__4454\,
            I => \eeprom.i2c.n11\
        );

    \I__870\ : InMux
    port map (
            O => \N__4451\,
            I => \N__4448\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4448\,
            I => \N__4445\
        );

    \I__868\ : Span4Mux_v
    port map (
            O => \N__4445\,
            I => \N__4440\
        );

    \I__867\ : InMux
    port map (
            O => \N__4444\,
            I => \N__4437\
        );

    \I__866\ : InMux
    port map (
            O => \N__4443\,
            I => \N__4434\
        );

    \I__865\ : Odrv4
    port map (
            O => \N__4440\,
            I => saved_addr_0
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4437\,
            I => saved_addr_0
        );

    \I__863\ : LocalMux
    port map (
            O => \N__4434\,
            I => saved_addr_0
        );

    \I__862\ : InMux
    port map (
            O => \N__4427\,
            I => \eeprom.i2c.n2511\
        );

    \I__861\ : InMux
    port map (
            O => \N__4424\,
            I => \eeprom.i2c.n2512\
        );

    \I__860\ : InMux
    port map (
            O => \N__4421\,
            I => \eeprom.i2c.n2513\
        );

    \I__859\ : InMux
    port map (
            O => \N__4418\,
            I => \eeprom.i2c.n2514\
        );

    \I__858\ : CascadeMux
    port map (
            O => \N__4415\,
            I => \N__4408\
        );

    \I__857\ : CascadeMux
    port map (
            O => \N__4414\,
            I => \N__4404\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__4413\,
            I => \N__4400\
        );

    \I__855\ : InMux
    port map (
            O => \N__4412\,
            I => \N__4385\
        );

    \I__854\ : InMux
    port map (
            O => \N__4411\,
            I => \N__4385\
        );

    \I__853\ : InMux
    port map (
            O => \N__4408\,
            I => \N__4385\
        );

    \I__852\ : InMux
    port map (
            O => \N__4407\,
            I => \N__4385\
        );

    \I__851\ : InMux
    port map (
            O => \N__4404\,
            I => \N__4385\
        );

    \I__850\ : InMux
    port map (
            O => \N__4403\,
            I => \N__4385\
        );

    \I__849\ : InMux
    port map (
            O => \N__4400\,
            I => \N__4385\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4385\,
            I => \CONSTANT_ONE_NET\
        );

    \I__847\ : InMux
    port map (
            O => \N__4382\,
            I => \eeprom.i2c.n2515\
        );

    \I__846\ : CEMux
    port map (
            O => \N__4379\,
            I => \N__4376\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__4376\,
            I => \N__4373\
        );

    \I__844\ : Odrv4
    port map (
            O => \N__4373\,
            I => \eeprom.i2c.n1413\
        );

    \I__843\ : SRMux
    port map (
            O => \N__4370\,
            I => \N__4367\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4367\,
            I => \N__4364\
        );

    \I__841\ : Span4Mux_h
    port map (
            O => \N__4364\,
            I => \N__4361\
        );

    \I__840\ : Odrv4
    port map (
            O => \N__4361\,
            I => \eeprom.i2c.n1495\
        );

    \I__839\ : InMux
    port map (
            O => \N__4358\,
            I => \N__4355\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__4355\,
            I => \eeprom.i2c.n2734\
        );

    \I__837\ : CascadeMux
    port map (
            O => \N__4352\,
            I => \N__4348\
        );

    \I__836\ : SRMux
    port map (
            O => \N__4351\,
            I => \N__4345\
        );

    \I__835\ : InMux
    port map (
            O => \N__4348\,
            I => \N__4342\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__4345\,
            I => \N__4338\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4342\,
            I => \N__4335\
        );

    \I__832\ : InMux
    port map (
            O => \N__4341\,
            I => \N__4332\
        );

    \I__831\ : Span4Mux_h
    port map (
            O => \N__4338\,
            I => \N__4329\
        );

    \I__830\ : Span4Mux_h
    port map (
            O => \N__4335\,
            I => \N__4324\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__4332\,
            I => \N__4324\
        );

    \I__828\ : Odrv4
    port map (
            O => \N__4329\,
            I => \eeprom.enable\
        );

    \I__827\ : Odrv4
    port map (
            O => \N__4324\,
            I => \eeprom.enable\
        );

    \I__826\ : InMux
    port map (
            O => \N__4319\,
            I => \N__4316\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__4316\,
            I => \eeprom.i2c.n2736\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__4313\,
            I => \N__4310\
        );

    \I__823\ : InMux
    port map (
            O => \N__4310\,
            I => \N__4307\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__4307\,
            I => \N__4304\
        );

    \I__821\ : Span4Mux_v
    port map (
            O => \N__4304\,
            I => \N__4301\
        );

    \I__820\ : Odrv4
    port map (
            O => \N__4301\,
            I => \eeprom.i2c.n2664\
        );

    \I__819\ : CascadeMux
    port map (
            O => \N__4298\,
            I => \n15_cascade_\
        );

    \I__818\ : InMux
    port map (
            O => \N__4295\,
            I => \N__4292\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__4292\,
            I => \N__4289\
        );

    \I__816\ : Odrv4
    port map (
            O => \N__4289\,
            I => \eeprom.i2c.n37\
        );

    \I__815\ : InMux
    port map (
            O => \N__4286\,
            I => \N__4283\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__4283\,
            I => \N__4280\
        );

    \I__813\ : Odrv12
    port map (
            O => \N__4280\,
            I => n7_adj_385
        );

    \I__812\ : InMux
    port map (
            O => \N__4277\,
            I => \bfn_21_14_0_\
        );

    \I__811\ : InMux
    port map (
            O => \N__4274\,
            I => \eeprom.i2c.n2509\
        );

    \I__810\ : InMux
    port map (
            O => \N__4271\,
            I => \eeprom.i2c.n2510\
        );

    \I__809\ : CascadeMux
    port map (
            O => \N__4268\,
            I => \eeprom.i2c.n2740_cascade_\
        );

    \I__808\ : InMux
    port map (
            O => \N__4265\,
            I => \N__4262\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__4262\,
            I => \eeprom.i2c.n970\
        );

    \I__806\ : CascadeMux
    port map (
            O => \N__4259\,
            I => \eeprom.i2c.n2747_cascade_\
        );

    \I__805\ : CascadeMux
    port map (
            O => \N__4256\,
            I => \eeprom.i2c.n15_adj_381_cascade_\
        );

    \I__804\ : InMux
    port map (
            O => \N__4253\,
            I => \N__4250\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__4250\,
            I => \eeprom.i2c.n2671\
        );

    \I__802\ : CascadeMux
    port map (
            O => \N__4247\,
            I => \eeprom.i2c.n2671_cascade_\
        );

    \I__801\ : CascadeMux
    port map (
            O => \N__4244\,
            I => \N__4241\
        );

    \I__800\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4238\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4238\,
            I => \N__4235\
        );

    \I__798\ : Span4Mux_h
    port map (
            O => \N__4235\,
            I => \N__4232\
        );

    \I__797\ : Span4Mux_v
    port map (
            O => \N__4232\,
            I => \N__4228\
        );

    \I__796\ : InMux
    port map (
            O => \N__4231\,
            I => \N__4225\
        );

    \I__795\ : Odrv4
    port map (
            O => \N__4228\,
            I => rw
        );

    \I__794\ : LocalMux
    port map (
            O => \N__4225\,
            I => rw
        );

    \I__793\ : InMux
    port map (
            O => \N__4220\,
            I => \N__4211\
        );

    \I__792\ : InMux
    port map (
            O => \N__4219\,
            I => \N__4211\
        );

    \I__791\ : InMux
    port map (
            O => \N__4218\,
            I => \N__4208\
        );

    \I__790\ : CascadeMux
    port map (
            O => \N__4217\,
            I => \N__4205\
        );

    \I__789\ : InMux
    port map (
            O => \N__4216\,
            I => \N__4202\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__4211\,
            I => \N__4197\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__4208\,
            I => \N__4197\
        );

    \I__786\ : InMux
    port map (
            O => \N__4205\,
            I => \N__4194\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__4202\,
            I => \N__4191\
        );

    \I__784\ : Span4Mux_v
    port map (
            O => \N__4197\,
            I => \N__4188\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__4194\,
            I => \N__4185\
        );

    \I__782\ : Span4Mux_v
    port map (
            O => \N__4191\,
            I => \N__4181\
        );

    \I__781\ : Sp12to4
    port map (
            O => \N__4188\,
            I => \N__4176\
        );

    \I__780\ : Span12Mux_v
    port map (
            O => \N__4185\,
            I => \N__4176\
        );

    \I__779\ : InMux
    port map (
            O => \N__4184\,
            I => \N__4173\
        );

    \I__778\ : Odrv4
    port map (
            O => \N__4181\,
            I => n15
        );

    \I__777\ : Odrv12
    port map (
            O => \N__4176\,
            I => n15
        );

    \I__776\ : LocalMux
    port map (
            O => \N__4173\,
            I => n15
        );

    \I__775\ : InMux
    port map (
            O => \N__4166\,
            I => \N__4160\
        );

    \I__774\ : InMux
    port map (
            O => \N__4165\,
            I => \N__4160\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__4160\,
            I => \state_7_N_269_0\
        );

    \I__772\ : InMux
    port map (
            O => \N__4157\,
            I => \N__4153\
        );

    \I__771\ : InMux
    port map (
            O => \N__4156\,
            I => \N__4150\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__4153\,
            I => \eeprom.i2c.counter2_0\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__4150\,
            I => \eeprom.i2c.counter2_0\
        );

    \I__768\ : InMux
    port map (
            O => \N__4145\,
            I => \bfn_19_17_0_\
        );

    \I__767\ : InMux
    port map (
            O => \N__4142\,
            I => \N__4138\
        );

    \I__766\ : InMux
    port map (
            O => \N__4141\,
            I => \N__4135\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__4138\,
            I => \eeprom.i2c.counter2_1\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__4135\,
            I => \eeprom.i2c.counter2_1\
        );

    \I__763\ : InMux
    port map (
            O => \N__4130\,
            I => \eeprom.i2c.n2531\
        );

    \I__762\ : InMux
    port map (
            O => \N__4127\,
            I => \N__4123\
        );

    \I__761\ : InMux
    port map (
            O => \N__4126\,
            I => \N__4120\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__4123\,
            I => \eeprom.i2c.counter2_2\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__4120\,
            I => \eeprom.i2c.counter2_2\
        );

    \I__758\ : InMux
    port map (
            O => \N__4115\,
            I => \eeprom.i2c.n2532\
        );

    \I__757\ : InMux
    port map (
            O => \N__4112\,
            I => \N__4108\
        );

    \I__756\ : InMux
    port map (
            O => \N__4111\,
            I => \N__4105\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__4108\,
            I => \eeprom.i2c.counter2_3\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__4105\,
            I => \eeprom.i2c.counter2_3\
        );

    \I__753\ : InMux
    port map (
            O => \N__4100\,
            I => \eeprom.i2c.n2533\
        );

    \I__752\ : InMux
    port map (
            O => \N__4097\,
            I => \eeprom.i2c.n2534\
        );

    \I__751\ : InMux
    port map (
            O => \N__4094\,
            I => \N__4090\
        );

    \I__750\ : InMux
    port map (
            O => \N__4093\,
            I => \N__4087\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__4090\,
            I => \eeprom.i2c.counter2_4\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__4087\,
            I => \eeprom.i2c.counter2_4\
        );

    \I__747\ : SRMux
    port map (
            O => \N__4082\,
            I => \N__4079\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__4079\,
            I => \N__4076\
        );

    \I__745\ : Span4Mux_h
    port map (
            O => \N__4076\,
            I => \N__4071\
        );

    \I__744\ : InMux
    port map (
            O => \N__4075\,
            I => \N__4068\
        );

    \I__743\ : InMux
    port map (
            O => \N__4074\,
            I => \N__4065\
        );

    \I__742\ : Odrv4
    port map (
            O => \N__4071\,
            I => \eeprom.i2c.counter2_7__N_256\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__4068\,
            I => \eeprom.i2c.counter2_7__N_256\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__4065\,
            I => \eeprom.i2c.counter2_7__N_256\
        );

    \I__739\ : CascadeMux
    port map (
            O => \N__4058\,
            I => \N__4053\
        );

    \I__738\ : InMux
    port map (
            O => \N__4057\,
            I => \N__4046\
        );

    \I__737\ : InMux
    port map (
            O => \N__4056\,
            I => \N__4046\
        );

    \I__736\ : InMux
    port map (
            O => \N__4053\,
            I => \N__4043\
        );

    \I__735\ : InMux
    port map (
            O => \N__4052\,
            I => \N__4040\
        );

    \I__734\ : InMux
    port map (
            O => \N__4051\,
            I => \N__4037\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__4046\,
            I => \N__4034\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__4043\,
            I => \N__4029\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4040\,
            I => \N__4029\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__4037\,
            I => \N__4026\
        );

    \I__729\ : Span4Mux_v
    port map (
            O => \N__4034\,
            I => \N__4021\
        );

    \I__728\ : Span4Mux_h
    port map (
            O => \N__4029\,
            I => \N__4021\
        );

    \I__727\ : Span12Mux_h
    port map (
            O => \N__4026\,
            I => \N__4018\
        );

    \I__726\ : Span4Mux_v
    port map (
            O => \N__4021\,
            I => \N__4015\
        );

    \I__725\ : Odrv12
    port map (
            O => \N__4018\,
            I => read
        );

    \I__724\ : Odrv4
    port map (
            O => \N__4015\,
            I => read
        );

    \I__723\ : InMux
    port map (
            O => \N__4010\,
            I => \N__4007\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4007\,
            I => \N__3995\
        );

    \I__721\ : InMux
    port map (
            O => \N__4006\,
            I => \N__3992\
        );

    \I__720\ : InMux
    port map (
            O => \N__4005\,
            I => \N__3987\
        );

    \I__719\ : InMux
    port map (
            O => \N__4004\,
            I => \N__3987\
        );

    \I__718\ : InMux
    port map (
            O => \N__4003\,
            I => \N__3978\
        );

    \I__717\ : InMux
    port map (
            O => \N__4002\,
            I => \N__3978\
        );

    \I__716\ : InMux
    port map (
            O => \N__4001\,
            I => \N__3978\
        );

    \I__715\ : InMux
    port map (
            O => \N__4000\,
            I => \N__3978\
        );

    \I__714\ : InMux
    port map (
            O => \N__3999\,
            I => \N__3973\
        );

    \I__713\ : InMux
    port map (
            O => \N__3998\,
            I => \N__3973\
        );

    \I__712\ : Odrv4
    port map (
            O => \N__3995\,
            I => state_0
        );

    \I__711\ : LocalMux
    port map (
            O => \N__3992\,
            I => state_0
        );

    \I__710\ : LocalMux
    port map (
            O => \N__3987\,
            I => state_0
        );

    \I__709\ : LocalMux
    port map (
            O => \N__3978\,
            I => state_0
        );

    \I__708\ : LocalMux
    port map (
            O => \N__3973\,
            I => state_0
        );

    \I__707\ : CascadeMux
    port map (
            O => \N__3962\,
            I => \N__3957\
        );

    \I__706\ : InMux
    port map (
            O => \N__3961\,
            I => \N__3954\
        );

    \I__705\ : InMux
    port map (
            O => \N__3960\,
            I => \N__3951\
        );

    \I__704\ : InMux
    port map (
            O => \N__3957\,
            I => \N__3948\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__3954\,
            I => \eeprom.n1338\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__3951\,
            I => \eeprom.n1338\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__3948\,
            I => \eeprom.n1338\
        );

    \I__700\ : ClkMux
    port map (
            O => \N__3941\,
            I => \N__3890\
        );

    \I__699\ : ClkMux
    port map (
            O => \N__3940\,
            I => \N__3890\
        );

    \I__698\ : ClkMux
    port map (
            O => \N__3939\,
            I => \N__3890\
        );

    \I__697\ : ClkMux
    port map (
            O => \N__3938\,
            I => \N__3890\
        );

    \I__696\ : ClkMux
    port map (
            O => \N__3937\,
            I => \N__3890\
        );

    \I__695\ : ClkMux
    port map (
            O => \N__3936\,
            I => \N__3890\
        );

    \I__694\ : ClkMux
    port map (
            O => \N__3935\,
            I => \N__3890\
        );

    \I__693\ : ClkMux
    port map (
            O => \N__3934\,
            I => \N__3890\
        );

    \I__692\ : ClkMux
    port map (
            O => \N__3933\,
            I => \N__3890\
        );

    \I__691\ : ClkMux
    port map (
            O => \N__3932\,
            I => \N__3890\
        );

    \I__690\ : ClkMux
    port map (
            O => \N__3931\,
            I => \N__3890\
        );

    \I__689\ : ClkMux
    port map (
            O => \N__3930\,
            I => \N__3890\
        );

    \I__688\ : ClkMux
    port map (
            O => \N__3929\,
            I => \N__3890\
        );

    \I__687\ : ClkMux
    port map (
            O => \N__3928\,
            I => \N__3890\
        );

    \I__686\ : ClkMux
    port map (
            O => \N__3927\,
            I => \N__3890\
        );

    \I__685\ : ClkMux
    port map (
            O => \N__3926\,
            I => \N__3890\
        );

    \I__684\ : ClkMux
    port map (
            O => \N__3925\,
            I => \N__3890\
        );

    \I__683\ : GlobalMux
    port map (
            O => \N__3890\,
            I => \N__3887\
        );

    \I__682\ : gio2CtrlBuf
    port map (
            O => \N__3887\,
            I => \CLK_c\
        );

    \I__681\ : SRMux
    port map (
            O => \N__3884\,
            I => \N__3881\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__3881\,
            I => \N__3878\
        );

    \I__679\ : Span4Mux_h
    port map (
            O => \N__3878\,
            I => \N__3870\
        );

    \I__678\ : InMux
    port map (
            O => \N__3877\,
            I => \N__3865\
        );

    \I__677\ : InMux
    port map (
            O => \N__3876\,
            I => \N__3865\
        );

    \I__676\ : InMux
    port map (
            O => \N__3875\,
            I => \N__3860\
        );

    \I__675\ : InMux
    port map (
            O => \N__3874\,
            I => \N__3860\
        );

    \I__674\ : InMux
    port map (
            O => \N__3873\,
            I => \N__3857\
        );

    \I__673\ : Odrv4
    port map (
            O => \N__3870\,
            I => state_1
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3865\,
            I => state_1
        );

    \I__671\ : LocalMux
    port map (
            O => \N__3860\,
            I => state_1
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3857\,
            I => state_1
        );

    \I__669\ : CascadeMux
    port map (
            O => \N__3848\,
            I => \n624_cascade_\
        );

    \I__668\ : CascadeMux
    port map (
            O => \N__3845\,
            I => \N__3842\
        );

    \I__667\ : InMux
    port map (
            O => \N__3842\,
            I => \N__3838\
        );

    \I__666\ : InMux
    port map (
            O => \N__3841\,
            I => \N__3835\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3838\,
            I => \eeprom.delay_counter_14\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__3835\,
            I => \eeprom.delay_counter_14\
        );

    \I__663\ : InMux
    port map (
            O => \N__3830\,
            I => \N__3826\
        );

    \I__662\ : InMux
    port map (
            O => \N__3829\,
            I => \N__3823\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__3826\,
            I => \eeprom.delay_counter_11\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3823\,
            I => \eeprom.delay_counter_11\
        );

    \I__659\ : CascadeMux
    port map (
            O => \N__3818\,
            I => \N__3814\
        );

    \I__658\ : InMux
    port map (
            O => \N__3817\,
            I => \N__3811\
        );

    \I__657\ : InMux
    port map (
            O => \N__3814\,
            I => \N__3808\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__3811\,
            I => \eeprom.delay_counter_15\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__3808\,
            I => \eeprom.delay_counter_15\
        );

    \I__654\ : InMux
    port map (
            O => \N__3803\,
            I => \N__3799\
        );

    \I__653\ : InMux
    port map (
            O => \N__3802\,
            I => \N__3796\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__3799\,
            I => \eeprom.delay_counter_9\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3796\,
            I => \eeprom.delay_counter_9\
        );

    \I__650\ : InMux
    port map (
            O => \N__3791\,
            I => \N__3787\
        );

    \I__649\ : InMux
    port map (
            O => \N__3790\,
            I => \N__3784\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__3787\,
            I => \eeprom.delay_counter_1\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3784\,
            I => \eeprom.delay_counter_1\
        );

    \I__646\ : InMux
    port map (
            O => \N__3779\,
            I => \N__3775\
        );

    \I__645\ : InMux
    port map (
            O => \N__3778\,
            I => \N__3772\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3775\,
            I => \eeprom.delay_counter_7\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__3772\,
            I => \eeprom.delay_counter_7\
        );

    \I__642\ : CascadeMux
    port map (
            O => \N__3767\,
            I => \eeprom.n2685_cascade_\
        );

    \I__641\ : InMux
    port map (
            O => \N__3764\,
            I => \N__3760\
        );

    \I__640\ : InMux
    port map (
            O => \N__3763\,
            I => \N__3757\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__3760\,
            I => \eeprom.delay_counter_3\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__3757\,
            I => \eeprom.delay_counter_3\
        );

    \I__637\ : InMux
    port map (
            O => \N__3752\,
            I => \N__3749\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__3749\,
            I => \eeprom.n22\
        );

    \I__635\ : InMux
    port map (
            O => \N__3746\,
            I => \N__3742\
        );

    \I__634\ : InMux
    port map (
            O => \N__3745\,
            I => \N__3739\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3742\,
            I => \eeprom.delay_counter_13\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__3739\,
            I => \eeprom.delay_counter_13\
        );

    \I__631\ : CascadeMux
    port map (
            O => \N__3734\,
            I => \N__3731\
        );

    \I__630\ : InMux
    port map (
            O => \N__3731\,
            I => \N__3727\
        );

    \I__629\ : InMux
    port map (
            O => \N__3730\,
            I => \N__3724\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__3727\,
            I => \eeprom.delay_counter_8\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__3724\,
            I => \eeprom.delay_counter_8\
        );

    \I__626\ : CascadeMux
    port map (
            O => \N__3719\,
            I => \N__3716\
        );

    \I__625\ : InMux
    port map (
            O => \N__3716\,
            I => \N__3712\
        );

    \I__624\ : InMux
    port map (
            O => \N__3715\,
            I => \N__3709\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3712\,
            I => \eeprom.delay_counter_4\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__3709\,
            I => \eeprom.delay_counter_4\
        );

    \I__621\ : InMux
    port map (
            O => \N__3704\,
            I => \N__3701\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__3701\,
            I => \eeprom.n20\
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__3698\,
            I => \eeprom.i2c.n6_cascade_\
        );

    \I__618\ : CascadeMux
    port map (
            O => \N__3695\,
            I => \eeprom.i2c.counter2_7__N_256_cascade_\
        );

    \I__617\ : CEMux
    port map (
            O => \N__3692\,
            I => \N__3689\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__3689\,
            I => \eeprom.i2c.n1384\
        );

    \I__615\ : CascadeMux
    port map (
            O => \N__3686\,
            I => \n6_adj_397_cascade_\
        );

    \I__614\ : CascadeMux
    port map (
            O => \N__3683\,
            I => \n2662_cascade_\
        );

    \I__613\ : InMux
    port map (
            O => \N__3680\,
            I => \N__3675\
        );

    \I__612\ : InMux
    port map (
            O => \N__3679\,
            I => \N__3670\
        );

    \I__611\ : InMux
    port map (
            O => \N__3678\,
            I => \N__3670\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__3675\,
            I => n2668
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3670\,
            I => n2668
        );

    \I__608\ : CascadeMux
    port map (
            O => \N__3665\,
            I => \N__3662\
        );

    \I__607\ : InMux
    port map (
            O => \N__3662\,
            I => \N__3658\
        );

    \I__606\ : InMux
    port map (
            O => \N__3661\,
            I => \N__3655\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3658\,
            I => \eeprom.delay_counter_0\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3655\,
            I => \eeprom.delay_counter_0\
        );

    \I__603\ : CascadeMux
    port map (
            O => \N__3650\,
            I => \N__3646\
        );

    \I__602\ : CascadeMux
    port map (
            O => \N__3649\,
            I => \N__3643\
        );

    \I__601\ : InMux
    port map (
            O => \N__3646\,
            I => \N__3640\
        );

    \I__600\ : InMux
    port map (
            O => \N__3643\,
            I => \N__3637\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3640\,
            I => \eeprom.delay_counter_2\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3637\,
            I => \eeprom.delay_counter_2\
        );

    \I__597\ : InMux
    port map (
            O => \N__3632\,
            I => \N__3628\
        );

    \I__596\ : InMux
    port map (
            O => \N__3631\,
            I => \N__3625\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3628\,
            I => \eeprom.delay_counter_5\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__3625\,
            I => \eeprom.delay_counter_5\
        );

    \I__593\ : CascadeMux
    port map (
            O => \N__3620\,
            I => \N__3617\
        );

    \I__592\ : InMux
    port map (
            O => \N__3617\,
            I => \N__3613\
        );

    \I__591\ : InMux
    port map (
            O => \N__3616\,
            I => \N__3610\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3613\,
            I => \eeprom.delay_counter_10\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3610\,
            I => \eeprom.delay_counter_10\
        );

    \I__588\ : CascadeMux
    port map (
            O => \N__3605\,
            I => \eeprom.n24_cascade_\
        );

    \I__587\ : CascadeMux
    port map (
            O => \N__3602\,
            I => \eeprom.n1338_cascade_\
        );

    \I__586\ : CascadeMux
    port map (
            O => \N__3599\,
            I => \N__3587\
        );

    \I__585\ : CascadeMux
    port map (
            O => \N__3598\,
            I => \N__3583\
        );

    \I__584\ : CascadeMux
    port map (
            O => \N__3597\,
            I => \N__3579\
        );

    \I__583\ : CascadeMux
    port map (
            O => \N__3596\,
            I => \N__3575\
        );

    \I__582\ : CascadeMux
    port map (
            O => \N__3595\,
            I => \N__3572\
        );

    \I__581\ : CascadeMux
    port map (
            O => \N__3594\,
            I => \N__3569\
        );

    \I__580\ : CascadeMux
    port map (
            O => \N__3593\,
            I => \N__3565\
        );

    \I__579\ : CascadeMux
    port map (
            O => \N__3592\,
            I => \N__3561\
        );

    \I__578\ : InMux
    port map (
            O => \N__3591\,
            I => \N__3543\
        );

    \I__577\ : InMux
    port map (
            O => \N__3590\,
            I => \N__3543\
        );

    \I__576\ : InMux
    port map (
            O => \N__3587\,
            I => \N__3543\
        );

    \I__575\ : InMux
    port map (
            O => \N__3586\,
            I => \N__3543\
        );

    \I__574\ : InMux
    port map (
            O => \N__3583\,
            I => \N__3543\
        );

    \I__573\ : InMux
    port map (
            O => \N__3582\,
            I => \N__3543\
        );

    \I__572\ : InMux
    port map (
            O => \N__3579\,
            I => \N__3543\
        );

    \I__571\ : InMux
    port map (
            O => \N__3578\,
            I => \N__3543\
        );

    \I__570\ : InMux
    port map (
            O => \N__3575\,
            I => \N__3540\
        );

    \I__569\ : InMux
    port map (
            O => \N__3572\,
            I => \N__3525\
        );

    \I__568\ : InMux
    port map (
            O => \N__3569\,
            I => \N__3525\
        );

    \I__567\ : InMux
    port map (
            O => \N__3568\,
            I => \N__3525\
        );

    \I__566\ : InMux
    port map (
            O => \N__3565\,
            I => \N__3525\
        );

    \I__565\ : InMux
    port map (
            O => \N__3564\,
            I => \N__3525\
        );

    \I__564\ : InMux
    port map (
            O => \N__3561\,
            I => \N__3525\
        );

    \I__563\ : InMux
    port map (
            O => \N__3560\,
            I => \N__3525\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3543\,
            I => \eeprom.n575\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__3540\,
            I => \eeprom.n575\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3525\,
            I => \eeprom.n575\
        );

    \I__559\ : CEMux
    port map (
            O => \N__3518\,
            I => \N__3514\
        );

    \I__558\ : CEMux
    port map (
            O => \N__3517\,
            I => \N__3511\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3514\,
            I => \eeprom.n1435\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__3511\,
            I => \eeprom.n1435\
        );

    \I__555\ : CascadeMux
    port map (
            O => \N__3506\,
            I => \eeprom.n1435_cascade_\
        );

    \I__554\ : SRMux
    port map (
            O => \N__3503\,
            I => \N__3499\
        );

    \I__553\ : SRMux
    port map (
            O => \N__3502\,
            I => \N__3496\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__3499\,
            I => \N__3493\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3496\,
            I => \eeprom.n1503\
        );

    \I__550\ : Odrv4
    port map (
            O => \N__3493\,
            I => \eeprom.n1503\
        );

    \I__549\ : InMux
    port map (
            O => \N__3488\,
            I => \N__3484\
        );

    \I__548\ : InMux
    port map (
            O => \N__3487\,
            I => \N__3481\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__3484\,
            I => \eeprom.delay_counter_6\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3481\,
            I => \eeprom.delay_counter_6\
        );

    \I__545\ : CascadeMux
    port map (
            O => \N__3476\,
            I => \N__3473\
        );

    \I__544\ : InMux
    port map (
            O => \N__3473\,
            I => \N__3469\
        );

    \I__543\ : InMux
    port map (
            O => \N__3472\,
            I => \N__3466\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__3469\,
            I => \eeprom.delay_counter_12\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3466\,
            I => \eeprom.delay_counter_12\
        );

    \I__540\ : InMux
    port map (
            O => \N__3461\,
            I => \N__3458\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3458\,
            I => \eeprom.n16\
        );

    \I__538\ : InMux
    port map (
            O => \N__3455\,
            I => \bfn_17_20_0_\
        );

    \I__537\ : InMux
    port map (
            O => \N__3452\,
            I => \eeprom.n2524\
        );

    \I__536\ : InMux
    port map (
            O => \N__3449\,
            I => \eeprom.n2525\
        );

    \I__535\ : InMux
    port map (
            O => \N__3446\,
            I => \eeprom.n2526\
        );

    \I__534\ : InMux
    port map (
            O => \N__3443\,
            I => \eeprom.n2527\
        );

    \I__533\ : InMux
    port map (
            O => \N__3440\,
            I => \eeprom.n2528\
        );

    \I__532\ : InMux
    port map (
            O => \N__3437\,
            I => \eeprom.n2529\
        );

    \I__531\ : InMux
    port map (
            O => \N__3434\,
            I => \eeprom.n2530\
        );

    \I__530\ : InMux
    port map (
            O => \N__3431\,
            I => \N__3428\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__3428\,
            I => n2077
        );

    \I__528\ : CascadeMux
    port map (
            O => \N__3425\,
            I => \n12_cascade_\
        );

    \I__527\ : InMux
    port map (
            O => \N__3422\,
            I => \eeprom.n2516\
        );

    \I__526\ : InMux
    port map (
            O => \N__3419\,
            I => \eeprom.n2517\
        );

    \I__525\ : InMux
    port map (
            O => \N__3416\,
            I => \eeprom.n2518\
        );

    \I__524\ : InMux
    port map (
            O => \N__3413\,
            I => \eeprom.n2519\
        );

    \I__523\ : InMux
    port map (
            O => \N__3410\,
            I => \eeprom.n2520\
        );

    \I__522\ : InMux
    port map (
            O => \N__3407\,
            I => \eeprom.n2521\
        );

    \I__521\ : InMux
    port map (
            O => \N__3404\,
            I => \eeprom.n2522\
        );

    \I__520\ : InMux
    port map (
            O => \N__3401\,
            I => \N__3397\
        );

    \I__519\ : InMux
    port map (
            O => \N__3400\,
            I => \N__3394\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__3397\,
            I => \N__3389\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3394\,
            I => \N__3389\
        );

    \I__516\ : Odrv4
    port map (
            O => \N__3389\,
            I => delay_counter_18
        );

    \I__515\ : InMux
    port map (
            O => \N__3386\,
            I => \N__3382\
        );

    \I__514\ : InMux
    port map (
            O => \N__3385\,
            I => \N__3379\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3382\,
            I => delay_counter_19
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3379\,
            I => delay_counter_19
        );

    \I__511\ : CascadeMux
    port map (
            O => \N__3374\,
            I => \n2721_cascade_\
        );

    \I__510\ : InMux
    port map (
            O => \N__3371\,
            I => \N__3367\
        );

    \I__509\ : InMux
    port map (
            O => \N__3370\,
            I => \N__3364\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__3367\,
            I => delay_counter_22
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3364\,
            I => delay_counter_22
        );

    \I__506\ : InMux
    port map (
            O => \N__3359\,
            I => \N__3355\
        );

    \I__505\ : InMux
    port map (
            O => \N__3358\,
            I => \N__3352\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__3355\,
            I => delay_counter_21
        );

    \I__503\ : LocalMux
    port map (
            O => \N__3352\,
            I => delay_counter_21
        );

    \I__502\ : InMux
    port map (
            O => \N__3347\,
            I => \N__3343\
        );

    \I__501\ : InMux
    port map (
            O => \N__3346\,
            I => \N__3340\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3343\,
            I => delay_counter_23
        );

    \I__499\ : LocalMux
    port map (
            O => \N__3340\,
            I => delay_counter_23
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__3335\,
            I => \n7_cascade_\
        );

    \I__497\ : InMux
    port map (
            O => \N__3332\,
            I => \N__3328\
        );

    \I__496\ : InMux
    port map (
            O => \N__3331\,
            I => \N__3325\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__3328\,
            I => \N__3322\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__3325\,
            I => delay_counter_20
        );

    \I__493\ : Odrv4
    port map (
            O => \N__3322\,
            I => delay_counter_20
        );

    \I__492\ : InMux
    port map (
            O => \N__3317\,
            I => \N__3313\
        );

    \I__491\ : InMux
    port map (
            O => \N__3316\,
            I => \N__3310\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3313\,
            I => delay_counter_29
        );

    \I__489\ : LocalMux
    port map (
            O => \N__3310\,
            I => delay_counter_29
        );

    \I__488\ : InMux
    port map (
            O => \N__3305\,
            I => \N__3301\
        );

    \I__487\ : InMux
    port map (
            O => \N__3304\,
            I => \N__3298\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3301\,
            I => delay_counter_25
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3298\,
            I => delay_counter_25
        );

    \I__484\ : CascadeMux
    port map (
            O => \N__3293\,
            I => \n2695_cascade_\
        );

    \I__483\ : InMux
    port map (
            O => \N__3290\,
            I => \N__3286\
        );

    \I__482\ : InMux
    port map (
            O => \N__3289\,
            I => \N__3283\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__3286\,
            I => delay_counter_28
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3283\,
            I => delay_counter_28
        );

    \I__479\ : CascadeMux
    port map (
            O => \N__3278\,
            I => \n13_cascade_\
        );

    \I__478\ : SRMux
    port map (
            O => \N__3275\,
            I => \N__3272\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3272\,
            I => \N__3269\
        );

    \I__476\ : Span4Mux_h
    port map (
            O => \N__3269\,
            I => \N__3263\
        );

    \I__475\ : SRMux
    port map (
            O => \N__3268\,
            I => \N__3260\
        );

    \I__474\ : SRMux
    port map (
            O => \N__3267\,
            I => \N__3257\
        );

    \I__473\ : SRMux
    port map (
            O => \N__3266\,
            I => \N__3254\
        );

    \I__472\ : Odrv4
    port map (
            O => \N__3263\,
            I => \addr_10__N_70\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__3260\,
            I => \addr_10__N_70\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3257\,
            I => \addr_10__N_70\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3254\,
            I => \addr_10__N_70\
        );

    \I__468\ : InMux
    port map (
            O => \N__3245\,
            I => \N__3240\
        );

    \I__467\ : InMux
    port map (
            O => \N__3244\,
            I => \N__3237\
        );

    \I__466\ : InMux
    port map (
            O => \N__3243\,
            I => \N__3234\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__3240\,
            I => delay_counter_31
        );

    \I__464\ : LocalMux
    port map (
            O => \N__3237\,
            I => delay_counter_31
        );

    \I__463\ : LocalMux
    port map (
            O => \N__3234\,
            I => delay_counter_31
        );

    \I__462\ : InMux
    port map (
            O => \N__3227\,
            I => \N__3224\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__3224\,
            I => n13
        );

    \I__460\ : InMux
    port map (
            O => \N__3221\,
            I => \N__3217\
        );

    \I__459\ : InMux
    port map (
            O => \N__3220\,
            I => \N__3214\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__3217\,
            I => delay_counter_26
        );

    \I__457\ : LocalMux
    port map (
            O => \N__3214\,
            I => delay_counter_26
        );

    \I__456\ : InMux
    port map (
            O => \N__3209\,
            I => \N__3205\
        );

    \I__455\ : InMux
    port map (
            O => \N__3208\,
            I => \N__3202\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__3205\,
            I => delay_counter_30
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3202\,
            I => delay_counter_30
        );

    \I__452\ : CascadeMux
    port map (
            O => \N__3197\,
            I => \N__3193\
        );

    \I__451\ : InMux
    port map (
            O => \N__3196\,
            I => \N__3190\
        );

    \I__450\ : InMux
    port map (
            O => \N__3193\,
            I => \N__3187\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__3190\,
            I => delay_counter_27
        );

    \I__448\ : LocalMux
    port map (
            O => \N__3187\,
            I => delay_counter_27
        );

    \I__447\ : InMux
    port map (
            O => \N__3182\,
            I => \N__3178\
        );

    \I__446\ : InMux
    port map (
            O => \N__3181\,
            I => \N__3175\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__3178\,
            I => delay_counter_24
        );

    \I__444\ : LocalMux
    port map (
            O => \N__3175\,
            I => delay_counter_24
        );

    \I__443\ : InMux
    port map (
            O => \N__3170\,
            I => \N__3164\
        );

    \I__442\ : InMux
    port map (
            O => \N__3169\,
            I => \N__3164\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__3164\,
            I => n14
        );

    \I__440\ : CascadeMux
    port map (
            O => \N__3161\,
            I => \n2077_cascade_\
        );

    \I__439\ : InMux
    port map (
            O => \N__3158\,
            I => n2508
        );

    \I__438\ : InMux
    port map (
            O => \N__3155\,
            I => \N__3151\
        );

    \I__437\ : InMux
    port map (
            O => \N__3154\,
            I => \N__3148\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__3151\,
            I => delay_counter_6
        );

    \I__435\ : LocalMux
    port map (
            O => \N__3148\,
            I => delay_counter_6
        );

    \I__434\ : InMux
    port map (
            O => \N__3143\,
            I => \N__3139\
        );

    \I__433\ : InMux
    port map (
            O => \N__3142\,
            I => \N__3136\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__3139\,
            I => delay_counter_0
        );

    \I__431\ : LocalMux
    port map (
            O => \N__3136\,
            I => delay_counter_0
        );

    \I__430\ : CascadeMux
    port map (
            O => \N__3131\,
            I => \N__3127\
        );

    \I__429\ : InMux
    port map (
            O => \N__3130\,
            I => \N__3124\
        );

    \I__428\ : InMux
    port map (
            O => \N__3127\,
            I => \N__3121\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3124\,
            I => delay_counter_9
        );

    \I__426\ : LocalMux
    port map (
            O => \N__3121\,
            I => delay_counter_9
        );

    \I__425\ : InMux
    port map (
            O => \N__3116\,
            I => \N__3112\
        );

    \I__424\ : InMux
    port map (
            O => \N__3115\,
            I => \N__3109\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__3112\,
            I => delay_counter_4
        );

    \I__422\ : LocalMux
    port map (
            O => \N__3109\,
            I => delay_counter_4
        );

    \I__421\ : InMux
    port map (
            O => \N__3104\,
            I => \N__3100\
        );

    \I__420\ : InMux
    port map (
            O => \N__3103\,
            I => \N__3097\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__3100\,
            I => delay_counter_2
        );

    \I__418\ : LocalMux
    port map (
            O => \N__3097\,
            I => delay_counter_2
        );

    \I__417\ : InMux
    port map (
            O => \N__3092\,
            I => \N__3088\
        );

    \I__416\ : InMux
    port map (
            O => \N__3091\,
            I => \N__3085\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__3088\,
            I => delay_counter_7
        );

    \I__414\ : LocalMux
    port map (
            O => \N__3085\,
            I => delay_counter_7
        );

    \I__413\ : CascadeMux
    port map (
            O => \N__3080\,
            I => \N__3076\
        );

    \I__412\ : InMux
    port map (
            O => \N__3079\,
            I => \N__3073\
        );

    \I__411\ : InMux
    port map (
            O => \N__3076\,
            I => \N__3070\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__3073\,
            I => delay_counter_5
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3070\,
            I => delay_counter_5
        );

    \I__408\ : InMux
    port map (
            O => \N__3065\,
            I => \N__3061\
        );

    \I__407\ : InMux
    port map (
            O => \N__3064\,
            I => \N__3058\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__3061\,
            I => delay_counter_3
        );

    \I__405\ : LocalMux
    port map (
            O => \N__3058\,
            I => delay_counter_3
        );

    \I__404\ : InMux
    port map (
            O => \N__3053\,
            I => \N__3049\
        );

    \I__403\ : InMux
    port map (
            O => \N__3052\,
            I => \N__3046\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__3049\,
            I => delay_counter_8
        );

    \I__401\ : LocalMux
    port map (
            O => \N__3046\,
            I => delay_counter_8
        );

    \I__400\ : InMux
    port map (
            O => \N__3041\,
            I => \N__3037\
        );

    \I__399\ : InMux
    port map (
            O => \N__3040\,
            I => \N__3034\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__3037\,
            I => delay_counter_1
        );

    \I__397\ : LocalMux
    port map (
            O => \N__3034\,
            I => delay_counter_1
        );

    \I__396\ : CascadeMux
    port map (
            O => \N__3029\,
            I => \N__3026\
        );

    \I__395\ : InMux
    port map (
            O => \N__3026\,
            I => \N__3023\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3023\,
            I => \N__3020\
        );

    \I__393\ : Odrv4
    port map (
            O => \N__3020\,
            I => n17
        );

    \I__392\ : InMux
    port map (
            O => \N__3017\,
            I => \N__3014\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__3014\,
            I => n16
        );

    \I__390\ : InMux
    port map (
            O => \N__3011\,
            I => \N__3007\
        );

    \I__389\ : InMux
    port map (
            O => \N__3010\,
            I => \N__3004\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__3007\,
            I => delay_counter_11
        );

    \I__387\ : LocalMux
    port map (
            O => \N__3004\,
            I => delay_counter_11
        );

    \I__386\ : InMux
    port map (
            O => \N__2999\,
            I => \N__2995\
        );

    \I__385\ : InMux
    port map (
            O => \N__2998\,
            I => \N__2992\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__2995\,
            I => delay_counter_10
        );

    \I__383\ : LocalMux
    port map (
            O => \N__2992\,
            I => delay_counter_10
        );

    \I__382\ : CascadeMux
    port map (
            O => \N__2987\,
            I => \n2722_cascade_\
        );

    \I__381\ : InMux
    port map (
            O => \N__2984\,
            I => \N__2980\
        );

    \I__380\ : InMux
    port map (
            O => \N__2983\,
            I => \N__2977\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2980\,
            I => delay_counter_12
        );

    \I__378\ : LocalMux
    port map (
            O => \N__2977\,
            I => delay_counter_12
        );

    \I__377\ : InMux
    port map (
            O => \N__2972\,
            I => \N__2968\
        );

    \I__376\ : InMux
    port map (
            O => \N__2971\,
            I => \N__2965\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__2968\,
            I => \N__2962\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__2965\,
            I => delay_counter_17
        );

    \I__373\ : Odrv4
    port map (
            O => \N__2962\,
            I => delay_counter_17
        );

    \I__372\ : InMux
    port map (
            O => \N__2957\,
            I => \N__2953\
        );

    \I__371\ : InMux
    port map (
            O => \N__2956\,
            I => \N__2950\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2953\,
            I => delay_counter_15
        );

    \I__369\ : LocalMux
    port map (
            O => \N__2950\,
            I => delay_counter_15
        );

    \I__368\ : InMux
    port map (
            O => \N__2945\,
            I => \N__2941\
        );

    \I__367\ : InMux
    port map (
            O => \N__2944\,
            I => \N__2938\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__2941\,
            I => delay_counter_14
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2938\,
            I => delay_counter_14
        );

    \I__364\ : InMux
    port map (
            O => \N__2933\,
            I => \N__2930\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__2930\,
            I => n8
        );

    \I__362\ : InMux
    port map (
            O => \N__2927\,
            I => \N__2923\
        );

    \I__361\ : InMux
    port map (
            O => \N__2926\,
            I => \N__2920\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__2923\,
            I => delay_counter_16
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2920\,
            I => delay_counter_16
        );

    \I__358\ : CascadeMux
    port map (
            O => \N__2915\,
            I => \N__2911\
        );

    \I__357\ : InMux
    port map (
            O => \N__2914\,
            I => \N__2908\
        );

    \I__356\ : InMux
    port map (
            O => \N__2911\,
            I => \N__2905\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__2908\,
            I => delay_counter_13
        );

    \I__354\ : LocalMux
    port map (
            O => \N__2905\,
            I => delay_counter_13
        );

    \I__353\ : InMux
    port map (
            O => \N__2900\,
            I => \N__2897\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__2897\,
            I => n2715
        );

    \I__351\ : InMux
    port map (
            O => \N__2894\,
            I => n2499
        );

    \I__350\ : InMux
    port map (
            O => \N__2891\,
            I => n2500
        );

    \I__349\ : InMux
    port map (
            O => \N__2888\,
            I => \bfn_14_24_0_\
        );

    \I__348\ : InMux
    port map (
            O => \N__2885\,
            I => n2502
        );

    \I__347\ : InMux
    port map (
            O => \N__2882\,
            I => n2503
        );

    \I__346\ : InMux
    port map (
            O => \N__2879\,
            I => n2504
        );

    \I__345\ : InMux
    port map (
            O => \N__2876\,
            I => n2505
        );

    \I__344\ : InMux
    port map (
            O => \N__2873\,
            I => n2506
        );

    \I__343\ : InMux
    port map (
            O => \N__2870\,
            I => n2507
        );

    \I__342\ : InMux
    port map (
            O => \N__2867\,
            I => n2490
        );

    \I__341\ : InMux
    port map (
            O => \N__2864\,
            I => n2491
        );

    \I__340\ : InMux
    port map (
            O => \N__2861\,
            I => n2492
        );

    \I__339\ : InMux
    port map (
            O => \N__2858\,
            I => \bfn_14_23_0_\
        );

    \I__338\ : InMux
    port map (
            O => \N__2855\,
            I => n2494
        );

    \I__337\ : InMux
    port map (
            O => \N__2852\,
            I => n2495
        );

    \I__336\ : InMux
    port map (
            O => \N__2849\,
            I => n2496
        );

    \I__335\ : InMux
    port map (
            O => \N__2846\,
            I => n2497
        );

    \I__334\ : InMux
    port map (
            O => \N__2843\,
            I => n2498
        );

    \I__333\ : InMux
    port map (
            O => \N__2840\,
            I => n2480
        );

    \I__332\ : InMux
    port map (
            O => \N__2837\,
            I => n2481
        );

    \I__331\ : InMux
    port map (
            O => \N__2834\,
            I => n2482
        );

    \I__330\ : InMux
    port map (
            O => \N__2831\,
            I => n2483
        );

    \I__329\ : InMux
    port map (
            O => \N__2828\,
            I => n2484
        );

    \I__328\ : InMux
    port map (
            O => \N__2825\,
            I => \bfn_14_22_0_\
        );

    \I__327\ : InMux
    port map (
            O => \N__2822\,
            I => n2486
        );

    \I__326\ : InMux
    port map (
            O => \N__2819\,
            I => n2487
        );

    \I__325\ : InMux
    port map (
            O => \N__2816\,
            I => n2488
        );

    \I__324\ : InMux
    port map (
            O => \N__2813\,
            I => n2489
        );

    \I__323\ : InMux
    port map (
            O => \N__2810\,
            I => \bfn_13_24_0_\
        );

    \I__322\ : InMux
    port map (
            O => \N__2807\,
            I => n2559
        );

    \I__321\ : InMux
    port map (
            O => \N__2804\,
            I => \N__2797\
        );

    \I__320\ : InMux
    port map (
            O => \N__2803\,
            I => \N__2797\
        );

    \I__319\ : InMux
    port map (
            O => \N__2802\,
            I => \N__2794\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__2797\,
            I => blink_counter_21
        );

    \I__317\ : LocalMux
    port map (
            O => \N__2794\,
            I => blink_counter_21
        );

    \I__316\ : InMux
    port map (
            O => \N__2789\,
            I => \N__2780\
        );

    \I__315\ : InMux
    port map (
            O => \N__2788\,
            I => \N__2780\
        );

    \I__314\ : InMux
    port map (
            O => \N__2787\,
            I => \N__2780\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__2780\,
            I => blink_counter_24
        );

    \I__312\ : CascadeMux
    port map (
            O => \N__2777\,
            I => \N__2773\
        );

    \I__311\ : CascadeMux
    port map (
            O => \N__2776\,
            I => \N__2770\
        );

    \I__310\ : InMux
    port map (
            O => \N__2773\,
            I => \N__2764\
        );

    \I__309\ : InMux
    port map (
            O => \N__2770\,
            I => \N__2764\
        );

    \I__308\ : InMux
    port map (
            O => \N__2769\,
            I => \N__2761\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2764\,
            I => blink_counter_23
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2761\,
            I => blink_counter_23
        );

    \I__305\ : InMux
    port map (
            O => \N__2756\,
            I => \N__2749\
        );

    \I__304\ : InMux
    port map (
            O => \N__2755\,
            I => \N__2749\
        );

    \I__303\ : InMux
    port map (
            O => \N__2754\,
            I => \N__2746\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2749\,
            I => blink_counter_22
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2746\,
            I => blink_counter_22
        );

    \I__300\ : InMux
    port map (
            O => \N__2741\,
            I => \N__2738\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2738\,
            I => n2730
        );

    \I__298\ : CascadeMux
    port map (
            O => \N__2735\,
            I => \n2731_cascade_\
        );

    \I__297\ : InMux
    port map (
            O => \N__2732\,
            I => \N__2726\
        );

    \I__296\ : InMux
    port map (
            O => \N__2731\,
            I => \N__2726\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2726\,
            I => blink_counter_25
        );

    \I__294\ : IoInMux
    port map (
            O => \N__2723\,
            I => \N__2720\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__2720\,
            I => \N__2717\
        );

    \I__292\ : Span4Mux_s3_v
    port map (
            O => \N__2717\,
            I => \N__2714\
        );

    \I__291\ : Sp12to4
    port map (
            O => \N__2714\,
            I => \N__2711\
        );

    \I__290\ : Span12Mux_h
    port map (
            O => \N__2711\,
            I => \N__2708\
        );

    \I__289\ : Odrv12
    port map (
            O => \N__2708\,
            I => \LED_c\
        );

    \I__288\ : InMux
    port map (
            O => \N__2705\,
            I => \bfn_14_21_0_\
        );

    \I__287\ : InMux
    port map (
            O => \N__2702\,
            I => n2478
        );

    \I__286\ : InMux
    port map (
            O => \N__2699\,
            I => n2479
        );

    \I__285\ : InMux
    port map (
            O => \N__2696\,
            I => \N__2693\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__2693\,
            I => n11
        );

    \I__283\ : InMux
    port map (
            O => \N__2690\,
            I => n2549
        );

    \I__282\ : InMux
    port map (
            O => \N__2687\,
            I => \N__2684\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2684\,
            I => n10
        );

    \I__280\ : InMux
    port map (
            O => \N__2681\,
            I => \bfn_13_23_0_\
        );

    \I__279\ : InMux
    port map (
            O => \N__2678\,
            I => \N__2675\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2675\,
            I => n9
        );

    \I__277\ : InMux
    port map (
            O => \N__2672\,
            I => n2551
        );

    \I__276\ : InMux
    port map (
            O => \N__2669\,
            I => \N__2666\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2666\,
            I => n8_adj_388
        );

    \I__274\ : InMux
    port map (
            O => \N__2663\,
            I => n2552
        );

    \I__273\ : InMux
    port map (
            O => \N__2660\,
            I => \N__2657\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__2657\,
            I => n7_adj_387
        );

    \I__271\ : InMux
    port map (
            O => \N__2654\,
            I => n2553
        );

    \I__270\ : InMux
    port map (
            O => \N__2651\,
            I => \N__2648\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__2648\,
            I => n6
        );

    \I__268\ : InMux
    port map (
            O => \N__2645\,
            I => n2554
        );

    \I__267\ : InMux
    port map (
            O => \N__2642\,
            I => n2555
        );

    \I__266\ : InMux
    port map (
            O => \N__2639\,
            I => n2556
        );

    \I__265\ : InMux
    port map (
            O => \N__2636\,
            I => n2557
        );

    \I__264\ : InMux
    port map (
            O => \N__2633\,
            I => \N__2630\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__2630\,
            I => n19
        );

    \I__262\ : InMux
    port map (
            O => \N__2627\,
            I => n2541
        );

    \I__261\ : InMux
    port map (
            O => \N__2624\,
            I => \N__2621\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__2621\,
            I => n18
        );

    \I__259\ : InMux
    port map (
            O => \N__2618\,
            I => \bfn_13_22_0_\
        );

    \I__258\ : InMux
    port map (
            O => \N__2615\,
            I => \N__2612\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__2612\,
            I => n17_adj_394
        );

    \I__256\ : InMux
    port map (
            O => \N__2609\,
            I => n2543
        );

    \I__255\ : InMux
    port map (
            O => \N__2606\,
            I => \N__2603\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__2603\,
            I => n16_adj_393
        );

    \I__253\ : InMux
    port map (
            O => \N__2600\,
            I => n2544
        );

    \I__252\ : InMux
    port map (
            O => \N__2597\,
            I => \N__2594\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__2594\,
            I => n15_adj_392
        );

    \I__250\ : InMux
    port map (
            O => \N__2591\,
            I => n2545
        );

    \I__249\ : InMux
    port map (
            O => \N__2588\,
            I => \N__2585\
        );

    \I__248\ : LocalMux
    port map (
            O => \N__2585\,
            I => n14_adj_391
        );

    \I__247\ : InMux
    port map (
            O => \N__2582\,
            I => n2546
        );

    \I__246\ : InMux
    port map (
            O => \N__2579\,
            I => \N__2576\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__2576\,
            I => n13_adj_390
        );

    \I__244\ : InMux
    port map (
            O => \N__2573\,
            I => n2547
        );

    \I__243\ : InMux
    port map (
            O => \N__2570\,
            I => \N__2567\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__2567\,
            I => n12_adj_389
        );

    \I__241\ : InMux
    port map (
            O => \N__2564\,
            I => n2548
        );

    \I__240\ : InMux
    port map (
            O => \N__2561\,
            I => \N__2558\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__2558\,
            I => n26
        );

    \I__238\ : InMux
    port map (
            O => \N__2555\,
            I => \bfn_13_21_0_\
        );

    \I__237\ : InMux
    port map (
            O => \N__2552\,
            I => \N__2549\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__2549\,
            I => n25
        );

    \I__235\ : InMux
    port map (
            O => \N__2546\,
            I => n2535
        );

    \I__234\ : InMux
    port map (
            O => \N__2543\,
            I => \N__2540\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__2540\,
            I => n24
        );

    \I__232\ : InMux
    port map (
            O => \N__2537\,
            I => n2536
        );

    \I__231\ : InMux
    port map (
            O => \N__2534\,
            I => \N__2531\
        );

    \I__230\ : LocalMux
    port map (
            O => \N__2531\,
            I => n23
        );

    \I__229\ : InMux
    port map (
            O => \N__2528\,
            I => n2537
        );

    \I__228\ : InMux
    port map (
            O => \N__2525\,
            I => \N__2522\
        );

    \I__227\ : LocalMux
    port map (
            O => \N__2522\,
            I => n22
        );

    \I__226\ : InMux
    port map (
            O => \N__2519\,
            I => n2538
        );

    \I__225\ : InMux
    port map (
            O => \N__2516\,
            I => \N__2513\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__2513\,
            I => n21
        );

    \I__223\ : InMux
    port map (
            O => \N__2510\,
            I => n2539
        );

    \I__222\ : InMux
    port map (
            O => \N__2507\,
            I => \N__2504\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__2504\,
            I => n20
        );

    \I__220\ : InMux
    port map (
            O => \N__2501\,
            I => n2540
        );

    \I__219\ : IoInMux
    port map (
            O => \N__2498\,
            I => \N__2495\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__2495\,
            I => \N__2492\
        );

    \I__217\ : IoSpan4Mux
    port map (
            O => \N__2492\,
            I => \N__2489\
        );

    \I__216\ : IoSpan4Mux
    port map (
            O => \N__2489\,
            I => \N__2486\
        );

    \I__215\ : IoSpan4Mux
    port map (
            O => \N__2486\,
            I => \N__2483\
        );

    \I__214\ : Odrv4
    port map (
            O => \N__2483\,
            I => \CLK_pad_gb_input\
        );

    \INVeeprom.i2c.i2c_scl_enable_124C\ : INV
    port map (
            O => \INVeeprom.i2c.i2c_scl_enable_124C_net\,
            I => \N__4974\
        );

    \INVeeprom.i2c.write_enable_132C\ : INV
    port map (
            O => \INVeeprom.i2c.write_enable_132C_net\,
            I => \N__4946\
        );

    \INVeeprom.i2c.sda_out_133C\ : INV
    port map (
            O => \INVeeprom.i2c.sda_out_133C_net\,
            I => \N__4975\
        );

    \IN_MUX_bfv_21_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_14_0_\
        );

    \IN_MUX_bfv_19_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_17_0_\
        );

    \IN_MUX_bfv_17_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_19_0_\
        );

    \IN_MUX_bfv_17_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n2523\,
            carryinitout => \bfn_17_20_0_\
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_21_0_\
        );

    \IN_MUX_bfv_14_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2485,
            carryinitout => \bfn_14_22_0_\
        );

    \IN_MUX_bfv_14_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2493,
            carryinitout => \bfn_14_23_0_\
        );

    \IN_MUX_bfv_14_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2501,
            carryinitout => \bfn_14_24_0_\
        );

    \IN_MUX_bfv_13_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_21_0_\
        );

    \IN_MUX_bfv_13_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2542,
            carryinitout => \bfn_13_22_0_\
        );

    \IN_MUX_bfv_13_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2550,
            carryinitout => \bfn_13_23_0_\
        );

    \IN_MUX_bfv_13_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2558,
            carryinitout => \bfn_13_24_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2498\,
            GLOBALBUFFEROUTPUT => \CLK_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \blink_counter_332__i0_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2561\,
            in2 => \_gnd_net_\,
            in3 => \N__2555\,
            lcout => n26,
            ltout => OPEN,
            carryin => \bfn_13_21_0_\,
            carryout => n2535,
            clk => \N__3925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i1_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2552\,
            in2 => \_gnd_net_\,
            in3 => \N__2546\,
            lcout => n25,
            ltout => OPEN,
            carryin => n2535,
            carryout => n2536,
            clk => \N__3925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i2_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2543\,
            in2 => \_gnd_net_\,
            in3 => \N__2537\,
            lcout => n24,
            ltout => OPEN,
            carryin => n2536,
            carryout => n2537,
            clk => \N__3925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i3_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2534\,
            in2 => \_gnd_net_\,
            in3 => \N__2528\,
            lcout => n23,
            ltout => OPEN,
            carryin => n2537,
            carryout => n2538,
            clk => \N__3925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i4_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2525\,
            in2 => \_gnd_net_\,
            in3 => \N__2519\,
            lcout => n22,
            ltout => OPEN,
            carryin => n2538,
            carryout => n2539,
            clk => \N__3925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i5_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2516\,
            in2 => \_gnd_net_\,
            in3 => \N__2510\,
            lcout => n21,
            ltout => OPEN,
            carryin => n2539,
            carryout => n2540,
            clk => \N__3925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i6_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2507\,
            in2 => \_gnd_net_\,
            in3 => \N__2501\,
            lcout => n20,
            ltout => OPEN,
            carryin => n2540,
            carryout => n2541,
            clk => \N__3925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i7_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2633\,
            in2 => \_gnd_net_\,
            in3 => \N__2627\,
            lcout => n19,
            ltout => OPEN,
            carryin => n2541,
            carryout => n2542,
            clk => \N__3925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i8_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2624\,
            in2 => \_gnd_net_\,
            in3 => \N__2618\,
            lcout => n18,
            ltout => OPEN,
            carryin => \bfn_13_22_0_\,
            carryout => n2543,
            clk => \N__3926\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i9_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2615\,
            in2 => \_gnd_net_\,
            in3 => \N__2609\,
            lcout => n17_adj_394,
            ltout => OPEN,
            carryin => n2543,
            carryout => n2544,
            clk => \N__3926\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i10_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2606\,
            in2 => \_gnd_net_\,
            in3 => \N__2600\,
            lcout => n16_adj_393,
            ltout => OPEN,
            carryin => n2544,
            carryout => n2545,
            clk => \N__3926\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i11_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2597\,
            in2 => \_gnd_net_\,
            in3 => \N__2591\,
            lcout => n15_adj_392,
            ltout => OPEN,
            carryin => n2545,
            carryout => n2546,
            clk => \N__3926\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i12_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2588\,
            in2 => \_gnd_net_\,
            in3 => \N__2582\,
            lcout => n14_adj_391,
            ltout => OPEN,
            carryin => n2546,
            carryout => n2547,
            clk => \N__3926\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i13_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2579\,
            in2 => \_gnd_net_\,
            in3 => \N__2573\,
            lcout => n13_adj_390,
            ltout => OPEN,
            carryin => n2547,
            carryout => n2548,
            clk => \N__3926\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i14_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2570\,
            in2 => \_gnd_net_\,
            in3 => \N__2564\,
            lcout => n12_adj_389,
            ltout => OPEN,
            carryin => n2548,
            carryout => n2549,
            clk => \N__3926\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i15_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2696\,
            in2 => \_gnd_net_\,
            in3 => \N__2690\,
            lcout => n11,
            ltout => OPEN,
            carryin => n2549,
            carryout => n2550,
            clk => \N__3926\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i16_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2687\,
            in2 => \_gnd_net_\,
            in3 => \N__2681\,
            lcout => n10,
            ltout => OPEN,
            carryin => \bfn_13_23_0_\,
            carryout => n2551,
            clk => \N__3930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i17_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2678\,
            in2 => \_gnd_net_\,
            in3 => \N__2672\,
            lcout => n9,
            ltout => OPEN,
            carryin => n2551,
            carryout => n2552,
            clk => \N__3930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i18_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2669\,
            in2 => \_gnd_net_\,
            in3 => \N__2663\,
            lcout => n8_adj_388,
            ltout => OPEN,
            carryin => n2552,
            carryout => n2553,
            clk => \N__3930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i19_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2660\,
            in2 => \_gnd_net_\,
            in3 => \N__2654\,
            lcout => n7_adj_387,
            ltout => OPEN,
            carryin => n2553,
            carryout => n2554,
            clk => \N__3930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i20_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2651\,
            in2 => \_gnd_net_\,
            in3 => \N__2645\,
            lcout => n6,
            ltout => OPEN,
            carryin => n2554,
            carryout => n2555,
            clk => \N__3930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i21_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2802\,
            in2 => \_gnd_net_\,
            in3 => \N__2642\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n2555,
            carryout => n2556,
            clk => \N__3930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i22_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2754\,
            in2 => \_gnd_net_\,
            in3 => \N__2639\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n2556,
            carryout => n2557,
            clk => \N__3930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i23_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2769\,
            in2 => \_gnd_net_\,
            in3 => \N__2636\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n2557,
            carryout => n2558,
            clk => \N__3930\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i24_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2787\,
            in2 => \_gnd_net_\,
            in3 => \N__2810\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_13_24_0_\,
            carryout => n2559,
            clk => \N__3933\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_332__i25_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2731\,
            in2 => \_gnd_net_\,
            in3 => \N__2807\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3933\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1846_4_lut_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000100010"
        )
    port map (
            in0 => \N__2803\,
            in1 => \N__2788\,
            in2 => \N__2776\,
            in3 => \N__2755\,
            lcout => n2730,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1847_4_lut_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011111000"
        )
    port map (
            in0 => \N__2804\,
            in1 => \N__2789\,
            in2 => \N__2777\,
            in3 => \N__2756\,
            lcout => OPEN,
            ltout => \n2731_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1848_3_lut_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__2741\,
            in1 => \_gnd_net_\,
            in2 => \N__2735\,
            in3 => \N__2732\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_counter_331__i0_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3143\,
            in2 => \_gnd_net_\,
            in3 => \N__2705\,
            lcout => delay_counter_0,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => n2478,
            clk => \N__3927\,
            ce => 'H',
            sr => \N__3275\
        );

    \delay_counter_331__i1_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3041\,
            in2 => \_gnd_net_\,
            in3 => \N__2702\,
            lcout => delay_counter_1,
            ltout => OPEN,
            carryin => n2478,
            carryout => n2479,
            clk => \N__3927\,
            ce => 'H',
            sr => \N__3275\
        );

    \delay_counter_331__i2_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3104\,
            in2 => \_gnd_net_\,
            in3 => \N__2699\,
            lcout => delay_counter_2,
            ltout => OPEN,
            carryin => n2479,
            carryout => n2480,
            clk => \N__3927\,
            ce => 'H',
            sr => \N__3275\
        );

    \delay_counter_331__i3_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3065\,
            in2 => \_gnd_net_\,
            in3 => \N__2840\,
            lcout => delay_counter_3,
            ltout => OPEN,
            carryin => n2480,
            carryout => n2481,
            clk => \N__3927\,
            ce => 'H',
            sr => \N__3275\
        );

    \delay_counter_331__i4_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3116\,
            in2 => \_gnd_net_\,
            in3 => \N__2837\,
            lcout => delay_counter_4,
            ltout => OPEN,
            carryin => n2481,
            carryout => n2482,
            clk => \N__3927\,
            ce => 'H',
            sr => \N__3275\
        );

    \delay_counter_331__i5_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3079\,
            in2 => \_gnd_net_\,
            in3 => \N__2834\,
            lcout => delay_counter_5,
            ltout => OPEN,
            carryin => n2482,
            carryout => n2483,
            clk => \N__3927\,
            ce => 'H',
            sr => \N__3275\
        );

    \delay_counter_331__i6_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3155\,
            in2 => \_gnd_net_\,
            in3 => \N__2831\,
            lcout => delay_counter_6,
            ltout => OPEN,
            carryin => n2483,
            carryout => n2484,
            clk => \N__3927\,
            ce => 'H',
            sr => \N__3275\
        );

    \delay_counter_331__i7_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3092\,
            in2 => \_gnd_net_\,
            in3 => \N__2828\,
            lcout => delay_counter_7,
            ltout => OPEN,
            carryin => n2484,
            carryout => n2485,
            clk => \N__3927\,
            ce => 'H',
            sr => \N__3275\
        );

    \delay_counter_331__i8_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3053\,
            in2 => \_gnd_net_\,
            in3 => \N__2825\,
            lcout => delay_counter_8,
            ltout => OPEN,
            carryin => \bfn_14_22_0_\,
            carryout => n2486,
            clk => \N__3931\,
            ce => 'H',
            sr => \N__3267\
        );

    \delay_counter_331__i9_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3130\,
            in2 => \_gnd_net_\,
            in3 => \N__2822\,
            lcout => delay_counter_9,
            ltout => OPEN,
            carryin => n2486,
            carryout => n2487,
            clk => \N__3931\,
            ce => 'H',
            sr => \N__3267\
        );

    \delay_counter_331__i10_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2999\,
            in2 => \_gnd_net_\,
            in3 => \N__2819\,
            lcout => delay_counter_10,
            ltout => OPEN,
            carryin => n2487,
            carryout => n2488,
            clk => \N__3931\,
            ce => 'H',
            sr => \N__3267\
        );

    \delay_counter_331__i11_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3011\,
            in2 => \_gnd_net_\,
            in3 => \N__2816\,
            lcout => delay_counter_11,
            ltout => OPEN,
            carryin => n2488,
            carryout => n2489,
            clk => \N__3931\,
            ce => 'H',
            sr => \N__3267\
        );

    \delay_counter_331__i12_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2984\,
            in2 => \_gnd_net_\,
            in3 => \N__2813\,
            lcout => delay_counter_12,
            ltout => OPEN,
            carryin => n2489,
            carryout => n2490,
            clk => \N__3931\,
            ce => 'H',
            sr => \N__3267\
        );

    \delay_counter_331__i13_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2914\,
            in2 => \_gnd_net_\,
            in3 => \N__2867\,
            lcout => delay_counter_13,
            ltout => OPEN,
            carryin => n2490,
            carryout => n2491,
            clk => \N__3931\,
            ce => 'H',
            sr => \N__3267\
        );

    \delay_counter_331__i14_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2945\,
            in2 => \_gnd_net_\,
            in3 => \N__2864\,
            lcout => delay_counter_14,
            ltout => OPEN,
            carryin => n2491,
            carryout => n2492,
            clk => \N__3931\,
            ce => 'H',
            sr => \N__3267\
        );

    \delay_counter_331__i15_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2957\,
            in2 => \_gnd_net_\,
            in3 => \N__2861\,
            lcout => delay_counter_15,
            ltout => OPEN,
            carryin => n2492,
            carryout => n2493,
            clk => \N__3931\,
            ce => 'H',
            sr => \N__3267\
        );

    \delay_counter_331__i16_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2927\,
            in2 => \_gnd_net_\,
            in3 => \N__2858\,
            lcout => delay_counter_16,
            ltout => OPEN,
            carryin => \bfn_14_23_0_\,
            carryout => n2494,
            clk => \N__3934\,
            ce => 'H',
            sr => \N__3266\
        );

    \delay_counter_331__i17_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2971\,
            in2 => \_gnd_net_\,
            in3 => \N__2855\,
            lcout => delay_counter_17,
            ltout => OPEN,
            carryin => n2494,
            carryout => n2495,
            clk => \N__3934\,
            ce => 'H',
            sr => \N__3266\
        );

    \delay_counter_331__i18_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3401\,
            in2 => \_gnd_net_\,
            in3 => \N__2852\,
            lcout => delay_counter_18,
            ltout => OPEN,
            carryin => n2495,
            carryout => n2496,
            clk => \N__3934\,
            ce => 'H',
            sr => \N__3266\
        );

    \delay_counter_331__i19_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3386\,
            in2 => \_gnd_net_\,
            in3 => \N__2849\,
            lcout => delay_counter_19,
            ltout => OPEN,
            carryin => n2496,
            carryout => n2497,
            clk => \N__3934\,
            ce => 'H',
            sr => \N__3266\
        );

    \delay_counter_331__i20_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3331\,
            in2 => \_gnd_net_\,
            in3 => \N__2846\,
            lcout => delay_counter_20,
            ltout => OPEN,
            carryin => n2497,
            carryout => n2498,
            clk => \N__3934\,
            ce => 'H',
            sr => \N__3266\
        );

    \delay_counter_331__i21_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3359\,
            in2 => \_gnd_net_\,
            in3 => \N__2843\,
            lcout => delay_counter_21,
            ltout => OPEN,
            carryin => n2498,
            carryout => n2499,
            clk => \N__3934\,
            ce => 'H',
            sr => \N__3266\
        );

    \delay_counter_331__i22_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3371\,
            in2 => \_gnd_net_\,
            in3 => \N__2894\,
            lcout => delay_counter_22,
            ltout => OPEN,
            carryin => n2499,
            carryout => n2500,
            clk => \N__3934\,
            ce => 'H',
            sr => \N__3266\
        );

    \delay_counter_331__i23_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3347\,
            in2 => \_gnd_net_\,
            in3 => \N__2891\,
            lcout => delay_counter_23,
            ltout => OPEN,
            carryin => n2500,
            carryout => n2501,
            clk => \N__3934\,
            ce => 'H',
            sr => \N__3266\
        );

    \delay_counter_331__i24_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3182\,
            in2 => \_gnd_net_\,
            in3 => \N__2888\,
            lcout => delay_counter_24,
            ltout => OPEN,
            carryin => \bfn_14_24_0_\,
            carryout => n2502,
            clk => \N__3939\,
            ce => 'H',
            sr => \N__3268\
        );

    \delay_counter_331__i25_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3305\,
            in2 => \_gnd_net_\,
            in3 => \N__2885\,
            lcout => delay_counter_25,
            ltout => OPEN,
            carryin => n2502,
            carryout => n2503,
            clk => \N__3939\,
            ce => 'H',
            sr => \N__3268\
        );

    \delay_counter_331__i26_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3221\,
            in2 => \_gnd_net_\,
            in3 => \N__2882\,
            lcout => delay_counter_26,
            ltout => OPEN,
            carryin => n2503,
            carryout => n2504,
            clk => \N__3939\,
            ce => 'H',
            sr => \N__3268\
        );

    \delay_counter_331__i27_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3196\,
            in2 => \_gnd_net_\,
            in3 => \N__2879\,
            lcout => delay_counter_27,
            ltout => OPEN,
            carryin => n2504,
            carryout => n2505,
            clk => \N__3939\,
            ce => 'H',
            sr => \N__3268\
        );

    \delay_counter_331__i28_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3290\,
            in2 => \_gnd_net_\,
            in3 => \N__2876\,
            lcout => delay_counter_28,
            ltout => OPEN,
            carryin => n2505,
            carryout => n2506,
            clk => \N__3939\,
            ce => 'H',
            sr => \N__3268\
        );

    \delay_counter_331__i29_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3317\,
            in2 => \_gnd_net_\,
            in3 => \N__2873\,
            lcout => delay_counter_29,
            ltout => OPEN,
            carryin => n2506,
            carryout => n2507,
            clk => \N__3939\,
            ce => 'H',
            sr => \N__3268\
        );

    \delay_counter_331__i30_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3209\,
            in2 => \_gnd_net_\,
            in3 => \N__2870\,
            lcout => delay_counter_30,
            ltout => OPEN,
            carryin => n2507,
            carryout => n2508,
            clk => \N__3939\,
            ce => 'H',
            sr => \N__3268\
        );

    \delay_counter_331__i31_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3245\,
            in2 => \_gnd_net_\,
            in3 => \N__3158\,
            lcout => delay_counter_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3939\,
            ce => 'H',
            sr => \N__3268\
        );

    \i6_4_lut_adj_15_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3154\,
            in1 => \N__3142\,
            in2 => \N__3131\,
            in3 => \N__3115\,
            lcout => n16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3103\,
            in1 => \N__3091\,
            in2 => \N__3080\,
            in3 => \N__3064\,
            lcout => n17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9_4_lut_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3052\,
            in1 => \N__3040\,
            in2 => \N__3029\,
            in3 => \N__3017\,
            lcout => OPEN,
            ltout => \n2722_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_17_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__3010\,
            in1 => \N__2998\,
            in2 => \N__2987\,
            in3 => \N__2983\,
            lcout => n2715,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_3_lut_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__2972\,
            in1 => \N__2956\,
            in2 => \_gnd_net_\,
            in3 => \N__2944\,
            lcout => n8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_adj_18_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__2933\,
            in1 => \N__2926\,
            in2 => \N__2915\,
            in3 => \N__2900\,
            lcout => OPEN,
            ltout => \n2721_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__3400\,
            in1 => \N__3385\,
            in2 => \N__3374\,
            in3 => \N__3370\,
            lcout => OPEN,
            ltout => \n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3358\,
            in1 => \N__3346\,
            in2 => \N__3335\,
            in3 => \N__3332\,
            lcout => OPEN,
            ltout => \n2695_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3316\,
            in1 => \N__3304\,
            in2 => \N__3293\,
            in3 => \N__3289\,
            lcout => n13,
            ltout => \n13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1200_3_lut_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3243\,
            in2 => \N__3278\,
            in3 => \N__3169\,
            lcout => \addr_10__N_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \read_15_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__3244\,
            in1 => \N__3170\,
            in2 => \_gnd_net_\,
            in3 => \N__3227\,
            lcout => read,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3220\,
            in1 => \N__3208\,
            in2 => \N__3197\,
            in3 => \N__3181\,
            lcout => n14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1275_2_lut_3_lut_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__4216\,
            in1 => \N__3876\,
            in2 => \_gnd_net_\,
            in3 => \N__4004\,
            lcout => n2077,
            ltout => \n2077_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.state__i0_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001000010000000"
        )
    port map (
            in0 => \N__4005\,
            in1 => \N__3680\,
            in2 => \N__3161\,
            in3 => \N__4057\,
            lcout => state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__4056\,
            in1 => \N__3877\,
            in2 => \_gnd_net_\,
            in3 => \N__3678\,
            lcout => OPEN,
            ltout => \n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.state__i1_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__3679\,
            in1 => \N__3431\,
            in2 => \N__3425\,
            in3 => \N__4006\,
            lcout => state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3928\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i0_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3560\,
            in2 => \N__3665\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.delay_counter_0\,
            ltout => OPEN,
            carryin => \bfn_17_19_0_\,
            carryout => \eeprom.n2516\,
            clk => \N__3932\,
            ce => \N__3517\,
            sr => \N__3503\
        );

    \eeprom.delay_counter_i0_i1_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3791\,
            in2 => \N__3592\,
            in3 => \N__3422\,
            lcout => \eeprom.delay_counter_1\,
            ltout => OPEN,
            carryin => \eeprom.n2516\,
            carryout => \eeprom.n2517\,
            clk => \N__3932\,
            ce => \N__3517\,
            sr => \N__3503\
        );

    \eeprom.delay_counter_i0_i2_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3564\,
            in2 => \N__3650\,
            in3 => \N__3419\,
            lcout => \eeprom.delay_counter_2\,
            ltout => OPEN,
            carryin => \eeprom.n2517\,
            carryout => \eeprom.n2518\,
            clk => \N__3932\,
            ce => \N__3517\,
            sr => \N__3503\
        );

    \eeprom.delay_counter_i0_i3_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3764\,
            in2 => \N__3593\,
            in3 => \N__3416\,
            lcout => \eeprom.delay_counter_3\,
            ltout => OPEN,
            carryin => \eeprom.n2518\,
            carryout => \eeprom.n2519\,
            clk => \N__3932\,
            ce => \N__3517\,
            sr => \N__3503\
        );

    \eeprom.delay_counter_i0_i4_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3568\,
            in2 => \N__3719\,
            in3 => \N__3413\,
            lcout => \eeprom.delay_counter_4\,
            ltout => OPEN,
            carryin => \eeprom.n2519\,
            carryout => \eeprom.n2520\,
            clk => \N__3932\,
            ce => \N__3517\,
            sr => \N__3503\
        );

    \eeprom.delay_counter_i0_i5_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3632\,
            in2 => \N__3594\,
            in3 => \N__3410\,
            lcout => \eeprom.delay_counter_5\,
            ltout => OPEN,
            carryin => \eeprom.n2520\,
            carryout => \eeprom.n2521\,
            clk => \N__3932\,
            ce => \N__3517\,
            sr => \N__3503\
        );

    \eeprom.delay_counter_i0_i6_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3488\,
            in2 => \N__3596\,
            in3 => \N__3407\,
            lcout => \eeprom.delay_counter_6\,
            ltout => OPEN,
            carryin => \eeprom.n2521\,
            carryout => \eeprom.n2522\,
            clk => \N__3932\,
            ce => \N__3517\,
            sr => \N__3503\
        );

    \eeprom.delay_counter_i0_i7_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3779\,
            in2 => \N__3595\,
            in3 => \N__3404\,
            lcout => \eeprom.delay_counter_7\,
            ltout => OPEN,
            carryin => \eeprom.n2522\,
            carryout => \eeprom.n2523\,
            clk => \N__3932\,
            ce => \N__3517\,
            sr => \N__3503\
        );

    \eeprom.delay_counter_i0_i8_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3578\,
            in2 => \N__3734\,
            in3 => \N__3455\,
            lcout => \eeprom.delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_17_20_0_\,
            carryout => \eeprom.n2524\,
            clk => \N__3935\,
            ce => \N__3518\,
            sr => \N__3502\
        );

    \eeprom.delay_counter_i0_i9_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3803\,
            in2 => \N__3597\,
            in3 => \N__3452\,
            lcout => \eeprom.delay_counter_9\,
            ltout => OPEN,
            carryin => \eeprom.n2524\,
            carryout => \eeprom.n2525\,
            clk => \N__3935\,
            ce => \N__3518\,
            sr => \N__3502\
        );

    \eeprom.delay_counter_i0_i10_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3582\,
            in2 => \N__3620\,
            in3 => \N__3449\,
            lcout => \eeprom.delay_counter_10\,
            ltout => OPEN,
            carryin => \eeprom.n2525\,
            carryout => \eeprom.n2526\,
            clk => \N__3935\,
            ce => \N__3518\,
            sr => \N__3502\
        );

    \eeprom.delay_counter_i0_i11_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3830\,
            in2 => \N__3598\,
            in3 => \N__3446\,
            lcout => \eeprom.delay_counter_11\,
            ltout => OPEN,
            carryin => \eeprom.n2526\,
            carryout => \eeprom.n2527\,
            clk => \N__3935\,
            ce => \N__3518\,
            sr => \N__3502\
        );

    \eeprom.delay_counter_i0_i12_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3586\,
            in2 => \N__3476\,
            in3 => \N__3443\,
            lcout => \eeprom.delay_counter_12\,
            ltout => OPEN,
            carryin => \eeprom.n2527\,
            carryout => \eeprom.n2528\,
            clk => \N__3935\,
            ce => \N__3518\,
            sr => \N__3502\
        );

    \eeprom.delay_counter_i0_i13_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3746\,
            in2 => \N__3599\,
            in3 => \N__3440\,
            lcout => \eeprom.delay_counter_13\,
            ltout => OPEN,
            carryin => \eeprom.n2528\,
            carryout => \eeprom.n2529\,
            clk => \N__3935\,
            ce => \N__3518\,
            sr => \N__3502\
        );

    \eeprom.delay_counter_i0_i14_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3590\,
            in2 => \N__3845\,
            in3 => \N__3437\,
            lcout => \eeprom.delay_counter_14\,
            ltout => OPEN,
            carryin => \eeprom.n2529\,
            carryout => \eeprom.n2530\,
            clk => \N__3935\,
            ce => \N__3518\,
            sr => \N__3502\
        );

    \eeprom.delay_counter_i0_i15_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__3591\,
            in1 => \N__3817\,
            in2 => \_gnd_net_\,
            in3 => \N__3434\,
            lcout => \eeprom.delay_counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3935\,
            ce => \N__3518\,
            sr => \N__3502\
        );

    \eeprom.i2_2_lut_adj_14_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3962\,
            in3 => \N__5579\,
            lcout => OPEN,
            ltout => \n6_adj_397_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1779_4_lut_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__3998\,
            in1 => \N__4286\,
            in2 => \N__3686\,
            in3 => \N__5429\,
            lcout => OPEN,
            ltout => \n2662_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1785_4_lut_4_lut_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__4218\,
            in1 => \N__3999\,
            in2 => \N__3683\,
            in3 => \N__3873\,
            lcout => n2668,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i11_4_lut_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3661\,
            in1 => \N__3461\,
            in2 => \N__3649\,
            in3 => \N__3752\,
            lcout => OPEN,
            ltout => \eeprom.n24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i12_4_lut_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3631\,
            in1 => \N__3616\,
            in2 => \N__3605\,
            in3 => \N__3704\,
            lcout => \eeprom.n1338\,
            ltout => \eeprom.n1338_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1902_2_lut_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3602\,
            in3 => \N__4219\,
            lcout => \eeprom.n575\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__4052\,
            in1 => \N__3874\,
            in2 => \_gnd_net_\,
            in3 => \N__4000\,
            lcout => \eeprom.n1435\,
            ltout => \eeprom.n1435_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i717_2_lut_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__4001\,
            in1 => \_gnd_net_\,
            in2 => \N__3506\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n1503\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i3_2_lut_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3487\,
            in2 => \_gnd_net_\,
            in3 => \N__3472\,
            lcout => \eeprom.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.mux_161_Mux_0_i1_4_lut_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__4002\,
            in1 => \N__4220\,
            in2 => \N__4058\,
            in3 => \N__3960\,
            lcout => OPEN,
            ltout => \n624_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rw_43_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010001010"
        )
    port map (
            in0 => \N__4231\,
            in1 => \N__3875\,
            in2 => \N__3848\,
            in3 => \N__4003\,
            lcout => rw,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3936\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i3_4_lut_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3841\,
            in1 => \N__3829\,
            in2 => \N__3818\,
            in3 => \N__3802\,
            lcout => OPEN,
            ltout => \eeprom.n2685_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i9_4_lut_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3790\,
            in1 => \N__3778\,
            in2 => \N__3767\,
            in3 => \N__3763\,
            lcout => \eeprom.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i7_3_lut_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__3745\,
            in1 => \N__3730\,
            in2 => \_gnd_net_\,
            in3 => \N__3715\,
            lcout => \eeprom.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.enable_slow_121_LC_19_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4896\,
            in2 => \_gnd_net_\,
            in3 => \N__4075\,
            lcout => \state_7_N_269_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3941\,
            ce => \N__3692\,
            sr => \N__4351\
        );

    \eeprom.i2c.i1_2_lut_LC_19_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4156\,
            in2 => \_gnd_net_\,
            in3 => \N__4093\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i4_4_lut_LC_19_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4141\,
            in1 => \N__4126\,
            in2 => \N__3698\,
            in3 => \N__4111\,
            lcout => \eeprom.i2c.counter2_7__N_256\,
            ltout => \eeprom.i2c.counter2_7__N_256_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_3_lut_LC_19_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__4894\,
            in1 => \_gnd_net_\,
            in2 => \N__3695\,
            in3 => \N__4341\,
            lcout => \eeprom.i2c.n1384\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2c_clk_122_LC_19_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__4895\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4074\,
            lcout => \eeprom.i2c.i2c_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3937\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.counter2_333_334__i1_LC_19_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4157\,
            in2 => \_gnd_net_\,
            in3 => \N__4145\,
            lcout => \eeprom.i2c.counter2_0\,
            ltout => OPEN,
            carryin => \bfn_19_17_0_\,
            carryout => \eeprom.i2c.n2531\,
            clk => \N__3929\,
            ce => 'H',
            sr => \N__4082\
        );

    \eeprom.i2c.counter2_333_334__i2_LC_19_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4142\,
            in2 => \_gnd_net_\,
            in3 => \N__4130\,
            lcout => \eeprom.i2c.counter2_1\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2531\,
            carryout => \eeprom.i2c.n2532\,
            clk => \N__3929\,
            ce => 'H',
            sr => \N__4082\
        );

    \eeprom.i2c.counter2_333_334__i3_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4127\,
            in2 => \_gnd_net_\,
            in3 => \N__4115\,
            lcout => \eeprom.i2c.counter2_2\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2532\,
            carryout => \eeprom.i2c.n2533\,
            clk => \N__3929\,
            ce => 'H',
            sr => \N__4082\
        );

    \eeprom.i2c.counter2_333_334__i4_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4112\,
            in2 => \_gnd_net_\,
            in3 => \N__4100\,
            lcout => \eeprom.i2c.counter2_3\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2533\,
            carryout => \eeprom.i2c.n2534\,
            clk => \N__3929\,
            ce => 'H',
            sr => \N__4082\
        );

    \eeprom.i2c.counter2_333_334__i5_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4094\,
            in2 => \_gnd_net_\,
            in3 => \N__4097\,
            lcout => \eeprom.i2c.counter2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3929\,
            ce => 'H',
            sr => \N__4082\
        );

    \eeprom.enable_39_LC_19_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000101110"
        )
    port map (
            in0 => \N__4051\,
            in1 => \N__4010\,
            in2 => \N__4217\,
            in3 => \N__3961\,
            lcout => \eeprom.enable\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3938\,
            ce => 'H',
            sr => \N__3884\
        );

    \eeprom.i2c.i1878_2_lut_3_lut_LC_20_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__4443\,
            in1 => \N__4820\,
            in2 => \_gnd_net_\,
            in3 => \N__4789\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n2740_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1880_4_lut_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__4790\,
            in1 => \N__4596\,
            in2 => \N__4268\,
            in3 => \N__5266\,
            lcout => \eeprom.i2c.n2734\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_3_lut_adj_11_LC_20_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__5546\,
            in1 => \N__5131\,
            in2 => \_gnd_net_\,
            in3 => \N__5424\,
            lcout => \eeprom.i2c.n970\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1881_2_lut_3_lut_LC_20_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4844\,
            in1 => \N__4821\,
            in2 => \_gnd_net_\,
            in3 => \N__4791\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n2747_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i17_4_lut_LC_20_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011101010"
        )
    port map (
            in0 => \N__4265\,
            in1 => \N__4295\,
            in2 => \N__4259\,
            in3 => \N__4253\,
            lcout => \eeprom.i2c.n1413\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_31_i11_2_lut_3_lut_4_lut_LC_20_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__5129\,
            in1 => \N__5270\,
            in2 => \N__5428\,
            in3 => \N__5566\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n15_adj_381_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1788_2_lut_3_lut_LC_20_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5706\,
            in2 => \N__4256\,
            in3 => \N__5650\,
            lcout => \eeprom.i2c.n2671\,
            ltout => \eeprom.i2c.n2671_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1787_2_lut_4_lut_LC_20_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5130\,
            in1 => \N__5420\,
            in2 => \N__4247\,
            in3 => \N__5568\,
            lcout => \eeprom.i2c.n1495\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.saved_addr__i1_LC_20_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__4166\,
            in1 => \N__4184\,
            in2 => \N__4244\,
            in3 => \N__4444\,
            lcout => saved_addr_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4954\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1844_2_lut_3_lut_4_lut_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5567\,
            in1 => \N__5419\,
            in2 => \N__5280\,
            in3 => \N__5128\,
            lcout => n15,
            ltout => \n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2_2_lut_LC_20_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__4165\,
            in1 => \_gnd_net_\,
            in2 => \N__4298\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.i2c.n2714\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_adj_9_LC_20_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5565\,
            in2 => \_gnd_net_\,
            in3 => \N__4535\,
            lcout => \eeprom.i2c.n37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i375_2_lut_LC_20_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5705\,
            in2 => \_gnd_net_\,
            in3 => \N__5649\,
            lcout => \state_7_N_285_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1781_2_lut_LC_20_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5573\,
            in2 => \_gnd_net_\,
            in3 => \N__5133\,
            lcout => \eeprom.i2c.n2664\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_145_i11_2_lut_3_lut_4_lut_LC_20_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__5574\,
            in1 => \N__5423\,
            in2 => \N__5281\,
            in3 => \N__5134\,
            lcout => \eeprom.i2c.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2_2_lut_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5278\,
            in2 => \_gnd_net_\,
            in3 => \N__5135\,
            lcout => n7_adj_385,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_21_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.counter_i0_LC_21_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4795\,
            in2 => \_gnd_net_\,
            in3 => \N__4277\,
            lcout => \eeprom.i2c.counter_0\,
            ltout => OPEN,
            carryin => \bfn_21_14_0_\,
            carryout => \eeprom.i2c.n2509\,
            clk => \N__4953\,
            ce => \N__4379\,
            sr => \N__4370\
        );

    \eeprom.i2c.counter_i1_LC_21_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4825\,
            in2 => \N__4413\,
            in3 => \N__4274\,
            lcout => \eeprom.i2c.counter_1\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2509\,
            carryout => \eeprom.i2c.n2510\,
            clk => \N__4953\,
            ce => \N__4379\,
            sr => \N__4370\
        );

    \eeprom.i2c.counter_i2_LC_21_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4403\,
            in2 => \N__4601\,
            in3 => \N__4271\,
            lcout => \eeprom.i2c.counter_2\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2510\,
            carryout => \eeprom.i2c.n2511\,
            clk => \N__4953\,
            ce => \N__4379\,
            sr => \N__4370\
        );

    \eeprom.i2c.counter_i3_LC_21_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4618\,
            in2 => \N__4414\,
            in3 => \N__4427\,
            lcout => \eeprom.i2c.counter_3\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2511\,
            carryout => \eeprom.i2c.n2512\,
            clk => \N__4953\,
            ce => \N__4379\,
            sr => \N__4370\
        );

    \eeprom.i2c.counter_i4_LC_21_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4407\,
            in2 => \N__4688\,
            in3 => \N__4424\,
            lcout => \eeprom.i2c.counter_4\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2512\,
            carryout => \eeprom.i2c.n2513\,
            clk => \N__4953\,
            ce => \N__4379\,
            sr => \N__4370\
        );

    \eeprom.i2c.counter_i5_LC_21_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4633\,
            in2 => \N__4415\,
            in3 => \N__4421\,
            lcout => \eeprom.i2c.counter_5\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2513\,
            carryout => \eeprom.i2c.n2514\,
            clk => \N__4953\,
            ce => \N__4379\,
            sr => \N__4370\
        );

    \eeprom.i2c.counter_i6_LC_21_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4411\,
            in2 => \N__4670\,
            in3 => \N__4418\,
            lcout => \eeprom.i2c.counter_6\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2514\,
            carryout => \eeprom.i2c.n2515\,
            clk => \N__4953\,
            ce => \N__4379\,
            sr => \N__4370\
        );

    \eeprom.i2c.counter_i7_LC_21_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__4412\,
            in1 => \N__4648\,
            in2 => \_gnd_net_\,
            in3 => \N__4382\,
            lcout => \eeprom.i2c.counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4953\,
            ce => \N__4379\,
            sr => \N__4370\
        );

    \eeprom.i2c.sda_out_133_LC_21_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011100"
        )
    port map (
            in0 => \N__5421\,
            in1 => \N__4358\,
            in2 => \N__4718\,
            in3 => \N__5132\,
            lcout => \eeprom.i2c.sda_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.sda_out_133C_net\,
            ce => \N__4544\,
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1865_4_lut_LC_21_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000011"
        )
    port map (
            in0 => \N__5682\,
            in1 => \N__5747\,
            in2 => \N__4352\,
            in3 => \N__4479\,
            lcout => \eeprom.i2c.n2736\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.write_enable_132_LC_21_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__4714\,
            in1 => \N__5422\,
            in2 => \_gnd_net_\,
            in3 => \N__5119\,
            lcout => sda_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.write_enable_132C_net\,
            ce => \N__4568\,
            sr => \N__4505\
        );

    \eeprom.i2c.state_i0_i3_LC_22_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100000001010"
        )
    port map (
            in0 => \N__5261\,
            in1 => \N__4319\,
            in2 => \N__4313\,
            in3 => \N__5399\,
            lcout => \eeprom.state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4956\,
            ce => \N__5631\,
            sr => \N__4577\
        );

    \eeprom.i2c.i1_2_lut_4_lut_LC_22_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100100010"
        )
    port map (
            in0 => \N__4530\,
            in1 => \N__5498\,
            in2 => \N__5236\,
            in3 => \N__4516\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1897_4_lut_4_lut_LC_22_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__4713\,
            in1 => \N__5200\,
            in2 => \N__4571\,
            in3 => \N__5067\,
            lcout => \eeprom.i2c.n952\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_4_lut_4_lut_LC_22_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001000"
        )
    port map (
            in0 => \N__5066\,
            in1 => \N__5193\,
            in2 => \N__5401\,
            in3 => \N__5499\,
            lcout => \eeprom.i2c.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i56_3_lut_LC_22_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5496\,
            in2 => \N__5400\,
            in3 => \N__5064\,
            lcout => \eeprom.i2c.n33\,
            ltout => \eeprom.i2c.n33_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_adj_13_LC_22_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4556\,
            in3 => \N__5194\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1891_4_lut_LC_22_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100110000"
        )
    port map (
            in0 => \N__5500\,
            in1 => \N__4553\,
            in2 => \N__4547\,
            in3 => \N__4531\,
            lcout => \eeprom.i2c.n2616\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i57_3_lut_3_lut_LC_22_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101100110"
        )
    port map (
            in0 => \N__5065\,
            in1 => \N__5356\,
            in2 => \_gnd_net_\,
            in3 => \N__5192\,
            lcout => \eeprom.i2c.n36\,
            ltout => \eeprom.i2c.n36_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_3_lut_4_lut_LC_22_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111010"
        )
    port map (
            in0 => \N__4517\,
            in1 => \N__5497\,
            in2 => \N__4508\,
            in3 => \N__5199\,
            lcout => \eeprom.i2c.n1493\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_i0_i1_LC_22_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001111100001111"
        )
    port map (
            in0 => \N__4697\,
            in1 => \N__4486\,
            in2 => \N__4463\,
            in3 => \N__4451\,
            lcout => \eeprom.state_1_adj_383\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4955\,
            ce => \N__5632\,
            sr => \N__4754\
        );

    \eeprom.i2c.i22_3_lut_3_lut_LC_22_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101000100"
        )
    port map (
            in0 => \N__5195\,
            in1 => \N__5535\,
            in2 => \_gnd_net_\,
            in3 => \N__5360\,
            lcout => \eeprom.i2c.n11_adj_377\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_25_i10_2_lut_LC_22_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5086\,
            in2 => \_gnd_net_\,
            in3 => \N__5562\,
            lcout => \eeprom.i2c.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_140_i11_2_lut_4_lut_LC_22_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__5415\,
            in1 => \N__5578\,
            in2 => \N__5279\,
            in3 => \N__5127\,
            lcout => \eeprom.i2c.n11_adj_378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1221_2_lut_LC_23_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5257\,
            in2 => \_gnd_net_\,
            in3 => \N__5364\,
            lcout => \eeprom.i2c.n2018\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i4_4_lut_adj_12_LC_23_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4687\,
            in1 => \N__4669\,
            in2 => \N__4652\,
            in3 => \N__4634\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n10_adj_380_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i5_3_lut_LC_23_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__4619\,
            in1 => \_gnd_net_\,
            in2 => \N__4604\,
            in3 => \N__4600\,
            lcout => \eeprom.i2c.n2654\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_3_lut_2_lut_LC_23_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__5365\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5260\,
            lcout => \eeprom.i2c.n2726\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1900_3_lut_4_lut_LC_23_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5125\,
            in1 => \N__5258\,
            in2 => \N__5633\,
            in3 => \N__5531\,
            lcout => \eeprom.i2c.n2706\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2_3_lut_4_lut_LC_23_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__5366\,
            in1 => \N__5259\,
            in2 => \N__5563\,
            in3 => \N__5123\,
            lcout => \eeprom.i2c.n11_adj_376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_4_lut_2_lut_4_lut_LC_23_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__5124\,
            in1 => \N__5530\,
            in2 => \_gnd_net_\,
            in3 => \N__5367\,
            lcout => \eeprom.i2c.n21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1904_4_lut_LC_23_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000000"
        )
    port map (
            in0 => \N__5746\,
            in1 => \N__4747\,
            in2 => \N__5588\,
            in3 => \N__5625\,
            lcout => \eeprom.i2c.n2008\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1264_3_lut_4_lut_LC_23_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101011"
        )
    port map (
            in0 => \N__5524\,
            in1 => \N__5068\,
            in2 => \N__5237\,
            in3 => \N__5395\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n2063_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_4_lut_LC_23_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__4840\,
            in1 => \N__4829\,
            in2 => \N__4802\,
            in3 => \N__4799\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n1358_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1888_4_lut_LC_23_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000111"
        )
    port map (
            in0 => \N__5526\,
            in1 => \N__5070\,
            in2 => \N__4769\,
            in3 => \N__5731\,
            lcout => \eeprom.i2c.n876\,
            ltout => \eeprom.i2c.n876_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1913_4_lut_LC_23_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011110000"
        )
    port map (
            in0 => \N__4766\,
            in1 => \N__5683\,
            in2 => \N__4757\,
            in3 => \N__4748\,
            lcout => \eeprom.i2c.n2078\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1874_4_lut_LC_23_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__4746\,
            in1 => \N__4736\,
            in2 => \N__5009\,
            in3 => \N__4730\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n2741_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_i0_i0_LC_23_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__5396\,
            in1 => \_gnd_net_\,
            in2 => \N__4721\,
            in3 => \N__5626\,
            lcout => state_0_adj_386,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4973\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_141_i10_2_lut_LC_23_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111011"
        )
    port map (
            in0 => \N__5525\,
            in1 => \N__5069\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.i2c.n10_adj_379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_i0_i2_LC_23_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000001000001010"
        )
    port map (
            in0 => \N__5732\,
            in1 => \N__5713\,
            in2 => \N__5684\,
            in3 => \N__5657\,
            lcout => \eeprom.state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4976\,
            ce => \N__5630\,
            sr => \N__5597\
        );

    \eeprom.i2c.i2c_scl_enable_124_LC_23_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__5569\,
            in1 => \N__5414\,
            in2 => \N__5262\,
            in3 => \N__5097\,
            lcout => scl_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.i2c_scl_enable_124C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_139_i9_2_lut_LC_24_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5397\,
            in2 => \_gnd_net_\,
            in3 => \N__5277\,
            lcout => \eeprom.i2c.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_139_i11_2_lut_4_lut_LC_24_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__5564\,
            in1 => \N__5398\,
            in2 => \N__5282\,
            in3 => \N__5126\,
            lcout => \eeprom.i2c.n11_adj_382\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1198_2_lut_LC_26_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4990\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4972\,
            lcout => scl_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
