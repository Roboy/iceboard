-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Feb 24 2020 16:35:42

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : inout std_logic;
    TX : inout std_logic;
    SDA : inout std_logic;
    SCL : inout std_logic;
    RX : inout std_logic;
    NEOPXL : out std_logic;
    LED : out std_logic;
    INLC : inout std_logic;
    INLB : inout std_logic;
    INLA : inout std_logic;
    INHC : inout std_logic;
    INHB : inout std_logic;
    INHA : inout std_logic;
    HALL3 : inout std_logic;
    HALL2 : inout std_logic;
    HALL1 : inout std_logic;
    FAULT_N : inout std_logic;
    ENCODER1_B : inout std_logic;
    ENCODER1_A : inout std_logic;
    ENCODER0_B : inout std_logic;
    ENCODER0_A : inout std_logic;
    DE : inout std_logic;
    CS_MISO : inout std_logic;
    CS_CLK : inout std_logic;
    CS : inout std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__51103\ : std_logic;
signal \N__51102\ : std_logic;
signal \N__51101\ : std_logic;
signal \N__51094\ : std_logic;
signal \N__51093\ : std_logic;
signal \N__51092\ : std_logic;
signal \N__51085\ : std_logic;
signal \N__51084\ : std_logic;
signal \N__51083\ : std_logic;
signal \N__51076\ : std_logic;
signal \N__51075\ : std_logic;
signal \N__51074\ : std_logic;
signal \N__51067\ : std_logic;
signal \N__51066\ : std_logic;
signal \N__51065\ : std_logic;
signal \N__51058\ : std_logic;
signal \N__51057\ : std_logic;
signal \N__51056\ : std_logic;
signal \N__51049\ : std_logic;
signal \N__51048\ : std_logic;
signal \N__51047\ : std_logic;
signal \N__51040\ : std_logic;
signal \N__51039\ : std_logic;
signal \N__51038\ : std_logic;
signal \N__51031\ : std_logic;
signal \N__51030\ : std_logic;
signal \N__51029\ : std_logic;
signal \N__51022\ : std_logic;
signal \N__51021\ : std_logic;
signal \N__51020\ : std_logic;
signal \N__51013\ : std_logic;
signal \N__51012\ : std_logic;
signal \N__51011\ : std_logic;
signal \N__51004\ : std_logic;
signal \N__51003\ : std_logic;
signal \N__51002\ : std_logic;
signal \N__50995\ : std_logic;
signal \N__50994\ : std_logic;
signal \N__50993\ : std_logic;
signal \N__50986\ : std_logic;
signal \N__50985\ : std_logic;
signal \N__50984\ : std_logic;
signal \N__50977\ : std_logic;
signal \N__50976\ : std_logic;
signal \N__50975\ : std_logic;
signal \N__50968\ : std_logic;
signal \N__50967\ : std_logic;
signal \N__50966\ : std_logic;
signal \N__50959\ : std_logic;
signal \N__50958\ : std_logic;
signal \N__50957\ : std_logic;
signal \N__50950\ : std_logic;
signal \N__50949\ : std_logic;
signal \N__50948\ : std_logic;
signal \N__50941\ : std_logic;
signal \N__50940\ : std_logic;
signal \N__50939\ : std_logic;
signal \N__50932\ : std_logic;
signal \N__50931\ : std_logic;
signal \N__50930\ : std_logic;
signal \N__50923\ : std_logic;
signal \N__50922\ : std_logic;
signal \N__50921\ : std_logic;
signal \N__50914\ : std_logic;
signal \N__50913\ : std_logic;
signal \N__50912\ : std_logic;
signal \N__50905\ : std_logic;
signal \N__50904\ : std_logic;
signal \N__50903\ : std_logic;
signal \N__50896\ : std_logic;
signal \N__50895\ : std_logic;
signal \N__50894\ : std_logic;
signal \N__50887\ : std_logic;
signal \N__50886\ : std_logic;
signal \N__50885\ : std_logic;
signal \N__50878\ : std_logic;
signal \N__50877\ : std_logic;
signal \N__50876\ : std_logic;
signal \N__50859\ : std_logic;
signal \N__50856\ : std_logic;
signal \N__50853\ : std_logic;
signal \N__50850\ : std_logic;
signal \N__50847\ : std_logic;
signal \N__50844\ : std_logic;
signal \N__50841\ : std_logic;
signal \N__50838\ : std_logic;
signal \N__50835\ : std_logic;
signal \N__50832\ : std_logic;
signal \N__50829\ : std_logic;
signal \N__50826\ : std_logic;
signal \N__50823\ : std_logic;
signal \N__50820\ : std_logic;
signal \N__50817\ : std_logic;
signal \N__50816\ : std_logic;
signal \N__50815\ : std_logic;
signal \N__50812\ : std_logic;
signal \N__50809\ : std_logic;
signal \N__50806\ : std_logic;
signal \N__50803\ : std_logic;
signal \N__50800\ : std_logic;
signal \N__50797\ : std_logic;
signal \N__50790\ : std_logic;
signal \N__50787\ : std_logic;
signal \N__50784\ : std_logic;
signal \N__50781\ : std_logic;
signal \N__50778\ : std_logic;
signal \N__50777\ : std_logic;
signal \N__50774\ : std_logic;
signal \N__50773\ : std_logic;
signal \N__50772\ : std_logic;
signal \N__50771\ : std_logic;
signal \N__50770\ : std_logic;
signal \N__50767\ : std_logic;
signal \N__50762\ : std_logic;
signal \N__50761\ : std_logic;
signal \N__50760\ : std_logic;
signal \N__50759\ : std_logic;
signal \N__50758\ : std_logic;
signal \N__50757\ : std_logic;
signal \N__50756\ : std_logic;
signal \N__50755\ : std_logic;
signal \N__50754\ : std_logic;
signal \N__50753\ : std_logic;
signal \N__50752\ : std_logic;
signal \N__50749\ : std_logic;
signal \N__50744\ : std_logic;
signal \N__50739\ : std_logic;
signal \N__50734\ : std_logic;
signal \N__50731\ : std_logic;
signal \N__50730\ : std_logic;
signal \N__50727\ : std_logic;
signal \N__50726\ : std_logic;
signal \N__50723\ : std_logic;
signal \N__50722\ : std_logic;
signal \N__50721\ : std_logic;
signal \N__50718\ : std_logic;
signal \N__50715\ : std_logic;
signal \N__50714\ : std_logic;
signal \N__50713\ : std_logic;
signal \N__50712\ : std_logic;
signal \N__50709\ : std_logic;
signal \N__50706\ : std_logic;
signal \N__50703\ : std_logic;
signal \N__50696\ : std_logic;
signal \N__50691\ : std_logic;
signal \N__50688\ : std_logic;
signal \N__50687\ : std_logic;
signal \N__50684\ : std_logic;
signal \N__50675\ : std_logic;
signal \N__50670\ : std_logic;
signal \N__50665\ : std_logic;
signal \N__50662\ : std_logic;
signal \N__50659\ : std_logic;
signal \N__50656\ : std_logic;
signal \N__50653\ : std_logic;
signal \N__50648\ : std_logic;
signal \N__50645\ : std_logic;
signal \N__50642\ : std_logic;
signal \N__50633\ : std_logic;
signal \N__50616\ : std_logic;
signal \N__50615\ : std_logic;
signal \N__50612\ : std_logic;
signal \N__50611\ : std_logic;
signal \N__50608\ : std_logic;
signal \N__50607\ : std_logic;
signal \N__50604\ : std_logic;
signal \N__50599\ : std_logic;
signal \N__50596\ : std_logic;
signal \N__50595\ : std_logic;
signal \N__50590\ : std_logic;
signal \N__50587\ : std_logic;
signal \N__50584\ : std_logic;
signal \N__50579\ : std_logic;
signal \N__50574\ : std_logic;
signal \N__50573\ : std_logic;
signal \N__50570\ : std_logic;
signal \N__50569\ : std_logic;
signal \N__50568\ : std_logic;
signal \N__50567\ : std_logic;
signal \N__50566\ : std_logic;
signal \N__50565\ : std_logic;
signal \N__50564\ : std_logic;
signal \N__50563\ : std_logic;
signal \N__50562\ : std_logic;
signal \N__50559\ : std_logic;
signal \N__50558\ : std_logic;
signal \N__50557\ : std_logic;
signal \N__50556\ : std_logic;
signal \N__50555\ : std_logic;
signal \N__50554\ : std_logic;
signal \N__50551\ : std_logic;
signal \N__50548\ : std_logic;
signal \N__50545\ : std_logic;
signal \N__50544\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50537\ : std_logic;
signal \N__50536\ : std_logic;
signal \N__50535\ : std_logic;
signal \N__50534\ : std_logic;
signal \N__50533\ : std_logic;
signal \N__50532\ : std_logic;
signal \N__50531\ : std_logic;
signal \N__50528\ : std_logic;
signal \N__50525\ : std_logic;
signal \N__50520\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50512\ : std_logic;
signal \N__50509\ : std_logic;
signal \N__50506\ : std_logic;
signal \N__50503\ : std_logic;
signal \N__50500\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50496\ : std_logic;
signal \N__50493\ : std_logic;
signal \N__50492\ : std_logic;
signal \N__50491\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50487\ : std_logic;
signal \N__50482\ : std_logic;
signal \N__50479\ : std_logic;
signal \N__50476\ : std_logic;
signal \N__50473\ : std_logic;
signal \N__50470\ : std_logic;
signal \N__50467\ : std_logic;
signal \N__50462\ : std_logic;
signal \N__50459\ : std_logic;
signal \N__50454\ : std_logic;
signal \N__50449\ : std_logic;
signal \N__50446\ : std_logic;
signal \N__50445\ : std_logic;
signal \N__50444\ : std_logic;
signal \N__50437\ : std_logic;
signal \N__50434\ : std_logic;
signal \N__50429\ : std_logic;
signal \N__50424\ : std_logic;
signal \N__50421\ : std_logic;
signal \N__50418\ : std_logic;
signal \N__50411\ : std_logic;
signal \N__50398\ : std_logic;
signal \N__50393\ : std_logic;
signal \N__50388\ : std_logic;
signal \N__50385\ : std_logic;
signal \N__50378\ : std_logic;
signal \N__50369\ : std_logic;
signal \N__50358\ : std_logic;
signal \N__50357\ : std_logic;
signal \N__50356\ : std_logic;
signal \N__50355\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50353\ : std_logic;
signal \N__50352\ : std_logic;
signal \N__50349\ : std_logic;
signal \N__50348\ : std_logic;
signal \N__50347\ : std_logic;
signal \N__50346\ : std_logic;
signal \N__50345\ : std_logic;
signal \N__50344\ : std_logic;
signal \N__50343\ : std_logic;
signal \N__50342\ : std_logic;
signal \N__50339\ : std_logic;
signal \N__50338\ : std_logic;
signal \N__50337\ : std_logic;
signal \N__50336\ : std_logic;
signal \N__50335\ : std_logic;
signal \N__50334\ : std_logic;
signal \N__50333\ : std_logic;
signal \N__50332\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50328\ : std_logic;
signal \N__50327\ : std_logic;
signal \N__50322\ : std_logic;
signal \N__50317\ : std_logic;
signal \N__50316\ : std_logic;
signal \N__50315\ : std_logic;
signal \N__50310\ : std_logic;
signal \N__50305\ : std_logic;
signal \N__50298\ : std_logic;
signal \N__50295\ : std_logic;
signal \N__50292\ : std_logic;
signal \N__50289\ : std_logic;
signal \N__50288\ : std_logic;
signal \N__50287\ : std_logic;
signal \N__50286\ : std_logic;
signal \N__50285\ : std_logic;
signal \N__50284\ : std_logic;
signal \N__50281\ : std_logic;
signal \N__50272\ : std_logic;
signal \N__50269\ : std_logic;
signal \N__50266\ : std_logic;
signal \N__50265\ : std_logic;
signal \N__50264\ : std_logic;
signal \N__50263\ : std_logic;
signal \N__50262\ : std_logic;
signal \N__50257\ : std_logic;
signal \N__50256\ : std_logic;
signal \N__50253\ : std_logic;
signal \N__50250\ : std_logic;
signal \N__50247\ : std_logic;
signal \N__50244\ : std_logic;
signal \N__50241\ : std_logic;
signal \N__50236\ : std_logic;
signal \N__50231\ : std_logic;
signal \N__50224\ : std_logic;
signal \N__50217\ : std_logic;
signal \N__50212\ : std_logic;
signal \N__50209\ : std_logic;
signal \N__50206\ : std_logic;
signal \N__50205\ : std_logic;
signal \N__50204\ : std_logic;
signal \N__50197\ : std_logic;
signal \N__50194\ : std_logic;
signal \N__50191\ : std_logic;
signal \N__50188\ : std_logic;
signal \N__50185\ : std_logic;
signal \N__50182\ : std_logic;
signal \N__50173\ : std_logic;
signal \N__50164\ : std_logic;
signal \N__50159\ : std_logic;
signal \N__50154\ : std_logic;
signal \N__50147\ : std_logic;
signal \N__50130\ : std_logic;
signal \N__50129\ : std_logic;
signal \N__50128\ : std_logic;
signal \N__50127\ : std_logic;
signal \N__50126\ : std_logic;
signal \N__50125\ : std_logic;
signal \N__50122\ : std_logic;
signal \N__50119\ : std_logic;
signal \N__50116\ : std_logic;
signal \N__50113\ : std_logic;
signal \N__50110\ : std_logic;
signal \N__50107\ : std_logic;
signal \N__50104\ : std_logic;
signal \N__50099\ : std_logic;
signal \N__50094\ : std_logic;
signal \N__50089\ : std_logic;
signal \N__50086\ : std_logic;
signal \N__50079\ : std_logic;
signal \N__50078\ : std_logic;
signal \N__50077\ : std_logic;
signal \N__50076\ : std_logic;
signal \N__50075\ : std_logic;
signal \N__50072\ : std_logic;
signal \N__50069\ : std_logic;
signal \N__50068\ : std_logic;
signal \N__50067\ : std_logic;
signal \N__50066\ : std_logic;
signal \N__50063\ : std_logic;
signal \N__50060\ : std_logic;
signal \N__50057\ : std_logic;
signal \N__50054\ : std_logic;
signal \N__50051\ : std_logic;
signal \N__50048\ : std_logic;
signal \N__50045\ : std_logic;
signal \N__50044\ : std_logic;
signal \N__50041\ : std_logic;
signal \N__50038\ : std_logic;
signal \N__50035\ : std_logic;
signal \N__50034\ : std_logic;
signal \N__50031\ : std_logic;
signal \N__50028\ : std_logic;
signal \N__50023\ : std_logic;
signal \N__50020\ : std_logic;
signal \N__50017\ : std_logic;
signal \N__50016\ : std_logic;
signal \N__50015\ : std_logic;
signal \N__50014\ : std_logic;
signal \N__50011\ : std_logic;
signal \N__50008\ : std_logic;
signal \N__50007\ : std_logic;
signal \N__50006\ : std_logic;
signal \N__50005\ : std_logic;
signal \N__50002\ : std_logic;
signal \N__50001\ : std_logic;
signal \N__50000\ : std_logic;
signal \N__49999\ : std_logic;
signal \N__49996\ : std_logic;
signal \N__49993\ : std_logic;
signal \N__49990\ : std_logic;
signal \N__49987\ : std_logic;
signal \N__49986\ : std_logic;
signal \N__49985\ : std_logic;
signal \N__49984\ : std_logic;
signal \N__49979\ : std_logic;
signal \N__49974\ : std_logic;
signal \N__49971\ : std_logic;
signal \N__49968\ : std_logic;
signal \N__49965\ : std_logic;
signal \N__49962\ : std_logic;
signal \N__49957\ : std_logic;
signal \N__49956\ : std_logic;
signal \N__49955\ : std_logic;
signal \N__49954\ : std_logic;
signal \N__49951\ : std_logic;
signal \N__49948\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49942\ : std_logic;
signal \N__49941\ : std_logic;
signal \N__49934\ : std_logic;
signal \N__49931\ : std_logic;
signal \N__49924\ : std_logic;
signal \N__49923\ : std_logic;
signal \N__49920\ : std_logic;
signal \N__49915\ : std_logic;
signal \N__49906\ : std_logic;
signal \N__49903\ : std_logic;
signal \N__49898\ : std_logic;
signal \N__49893\ : std_logic;
signal \N__49890\ : std_logic;
signal \N__49885\ : std_logic;
signal \N__49878\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49868\ : std_logic;
signal \N__49851\ : std_logic;
signal \N__49850\ : std_logic;
signal \N__49847\ : std_logic;
signal \N__49844\ : std_logic;
signal \N__49843\ : std_logic;
signal \N__49842\ : std_logic;
signal \N__49839\ : std_logic;
signal \N__49838\ : std_logic;
signal \N__49835\ : std_logic;
signal \N__49834\ : std_logic;
signal \N__49831\ : std_logic;
signal \N__49830\ : std_logic;
signal \N__49829\ : std_logic;
signal \N__49828\ : std_logic;
signal \N__49825\ : std_logic;
signal \N__49822\ : std_logic;
signal \N__49819\ : std_logic;
signal \N__49818\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49812\ : std_logic;
signal \N__49811\ : std_logic;
signal \N__49808\ : std_logic;
signal \N__49807\ : std_logic;
signal \N__49804\ : std_logic;
signal \N__49803\ : std_logic;
signal \N__49800\ : std_logic;
signal \N__49797\ : std_logic;
signal \N__49796\ : std_logic;
signal \N__49793\ : std_logic;
signal \N__49790\ : std_logic;
signal \N__49787\ : std_logic;
signal \N__49784\ : std_logic;
signal \N__49779\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49775\ : std_logic;
signal \N__49774\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49772\ : std_logic;
signal \N__49771\ : std_logic;
signal \N__49768\ : std_logic;
signal \N__49765\ : std_logic;
signal \N__49762\ : std_logic;
signal \N__49759\ : std_logic;
signal \N__49758\ : std_logic;
signal \N__49757\ : std_logic;
signal \N__49754\ : std_logic;
signal \N__49753\ : std_logic;
signal \N__49752\ : std_logic;
signal \N__49751\ : std_logic;
signal \N__49750\ : std_logic;
signal \N__49749\ : std_logic;
signal \N__49746\ : std_logic;
signal \N__49743\ : std_logic;
signal \N__49738\ : std_logic;
signal \N__49735\ : std_logic;
signal \N__49730\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49722\ : std_logic;
signal \N__49719\ : std_logic;
signal \N__49716\ : std_logic;
signal \N__49713\ : std_logic;
signal \N__49704\ : std_logic;
signal \N__49701\ : std_logic;
signal \N__49698\ : std_logic;
signal \N__49697\ : std_logic;
signal \N__49694\ : std_logic;
signal \N__49691\ : std_logic;
signal \N__49688\ : std_logic;
signal \N__49685\ : std_logic;
signal \N__49680\ : std_logic;
signal \N__49677\ : std_logic;
signal \N__49674\ : std_logic;
signal \N__49665\ : std_logic;
signal \N__49662\ : std_logic;
signal \N__49659\ : std_logic;
signal \N__49656\ : std_logic;
signal \N__49649\ : std_logic;
signal \N__49646\ : std_logic;
signal \N__49643\ : std_logic;
signal \N__49638\ : std_logic;
signal \N__49633\ : std_logic;
signal \N__49620\ : std_logic;
signal \N__49615\ : std_logic;
signal \N__49602\ : std_logic;
signal \N__49601\ : std_logic;
signal \N__49600\ : std_logic;
signal \N__49597\ : std_logic;
signal \N__49594\ : std_logic;
signal \N__49593\ : std_logic;
signal \N__49590\ : std_logic;
signal \N__49589\ : std_logic;
signal \N__49588\ : std_logic;
signal \N__49585\ : std_logic;
signal \N__49582\ : std_logic;
signal \N__49581\ : std_logic;
signal \N__49580\ : std_logic;
signal \N__49577\ : std_logic;
signal \N__49574\ : std_logic;
signal \N__49571\ : std_logic;
signal \N__49570\ : std_logic;
signal \N__49567\ : std_logic;
signal \N__49564\ : std_logic;
signal \N__49561\ : std_logic;
signal \N__49558\ : std_logic;
signal \N__49555\ : std_logic;
signal \N__49554\ : std_logic;
signal \N__49553\ : std_logic;
signal \N__49548\ : std_logic;
signal \N__49545\ : std_logic;
signal \N__49542\ : std_logic;
signal \N__49539\ : std_logic;
signal \N__49536\ : std_logic;
signal \N__49533\ : std_logic;
signal \N__49528\ : std_logic;
signal \N__49527\ : std_logic;
signal \N__49526\ : std_logic;
signal \N__49525\ : std_logic;
signal \N__49524\ : std_logic;
signal \N__49521\ : std_logic;
signal \N__49518\ : std_logic;
signal \N__49517\ : std_logic;
signal \N__49516\ : std_logic;
signal \N__49511\ : std_logic;
signal \N__49510\ : std_logic;
signal \N__49509\ : std_logic;
signal \N__49508\ : std_logic;
signal \N__49503\ : std_logic;
signal \N__49498\ : std_logic;
signal \N__49495\ : std_logic;
signal \N__49490\ : std_logic;
signal \N__49489\ : std_logic;
signal \N__49484\ : std_logic;
signal \N__49481\ : std_logic;
signal \N__49478\ : std_logic;
signal \N__49475\ : std_logic;
signal \N__49472\ : std_logic;
signal \N__49469\ : std_logic;
signal \N__49466\ : std_logic;
signal \N__49463\ : std_logic;
signal \N__49460\ : std_logic;
signal \N__49455\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49447\ : std_logic;
signal \N__49444\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49426\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49412\ : std_logic;
signal \N__49411\ : std_logic;
signal \N__49410\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49406\ : std_logic;
signal \N__49403\ : std_logic;
signal \N__49396\ : std_logic;
signal \N__49393\ : std_logic;
signal \N__49390\ : std_logic;
signal \N__49387\ : std_logic;
signal \N__49384\ : std_logic;
signal \N__49381\ : std_logic;
signal \N__49378\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49368\ : std_logic;
signal \N__49365\ : std_logic;
signal \N__49362\ : std_logic;
signal \N__49359\ : std_logic;
signal \N__49356\ : std_logic;
signal \N__49353\ : std_logic;
signal \N__49350\ : std_logic;
signal \N__49349\ : std_logic;
signal \N__49346\ : std_logic;
signal \N__49343\ : std_logic;
signal \N__49340\ : std_logic;
signal \N__49337\ : std_logic;
signal \N__49334\ : std_logic;
signal \N__49331\ : std_logic;
signal \N__49326\ : std_logic;
signal \N__49323\ : std_logic;
signal \N__49320\ : std_logic;
signal \N__49317\ : std_logic;
signal \N__49314\ : std_logic;
signal \N__49311\ : std_logic;
signal \N__49308\ : std_logic;
signal \N__49305\ : std_logic;
signal \N__49302\ : std_logic;
signal \N__49299\ : std_logic;
signal \N__49296\ : std_logic;
signal \N__49293\ : std_logic;
signal \N__49290\ : std_logic;
signal \N__49287\ : std_logic;
signal \N__49284\ : std_logic;
signal \N__49283\ : std_logic;
signal \N__49280\ : std_logic;
signal \N__49277\ : std_logic;
signal \N__49272\ : std_logic;
signal \N__49269\ : std_logic;
signal \N__49266\ : std_logic;
signal \N__49263\ : std_logic;
signal \N__49260\ : std_logic;
signal \N__49259\ : std_logic;
signal \N__49256\ : std_logic;
signal \N__49253\ : std_logic;
signal \N__49250\ : std_logic;
signal \N__49247\ : std_logic;
signal \N__49242\ : std_logic;
signal \N__49239\ : std_logic;
signal \N__49236\ : std_logic;
signal \N__49233\ : std_logic;
signal \N__49230\ : std_logic;
signal \N__49227\ : std_logic;
signal \N__49226\ : std_logic;
signal \N__49223\ : std_logic;
signal \N__49220\ : std_logic;
signal \N__49217\ : std_logic;
signal \N__49214\ : std_logic;
signal \N__49211\ : std_logic;
signal \N__49208\ : std_logic;
signal \N__49203\ : std_logic;
signal \N__49200\ : std_logic;
signal \N__49197\ : std_logic;
signal \N__49194\ : std_logic;
signal \N__49191\ : std_logic;
signal \N__49188\ : std_logic;
signal \N__49187\ : std_logic;
signal \N__49184\ : std_logic;
signal \N__49181\ : std_logic;
signal \N__49178\ : std_logic;
signal \N__49175\ : std_logic;
signal \N__49172\ : std_logic;
signal \N__49169\ : std_logic;
signal \N__49166\ : std_logic;
signal \N__49163\ : std_logic;
signal \N__49160\ : std_logic;
signal \N__49157\ : std_logic;
signal \N__49152\ : std_logic;
signal \N__49149\ : std_logic;
signal \N__49146\ : std_logic;
signal \N__49145\ : std_logic;
signal \N__49144\ : std_logic;
signal \N__49143\ : std_logic;
signal \N__49142\ : std_logic;
signal \N__49141\ : std_logic;
signal \N__49138\ : std_logic;
signal \N__49133\ : std_logic;
signal \N__49130\ : std_logic;
signal \N__49127\ : std_logic;
signal \N__49124\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49095\ : std_logic;
signal \N__49092\ : std_logic;
signal \N__49091\ : std_logic;
signal \N__49088\ : std_logic;
signal \N__49085\ : std_logic;
signal \N__49082\ : std_logic;
signal \N__49079\ : std_logic;
signal \N__49076\ : std_logic;
signal \N__49073\ : std_logic;
signal \N__49068\ : std_logic;
signal \N__49065\ : std_logic;
signal \N__49062\ : std_logic;
signal \N__49059\ : std_logic;
signal \N__49056\ : std_logic;
signal \N__49053\ : std_logic;
signal \N__49050\ : std_logic;
signal \N__49049\ : std_logic;
signal \N__49048\ : std_logic;
signal \N__49045\ : std_logic;
signal \N__49044\ : std_logic;
signal \N__49043\ : std_logic;
signal \N__49042\ : std_logic;
signal \N__49041\ : std_logic;
signal \N__49040\ : std_logic;
signal \N__49037\ : std_logic;
signal \N__49034\ : std_logic;
signal \N__49033\ : std_logic;
signal \N__49032\ : std_logic;
signal \N__49031\ : std_logic;
signal \N__49030\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49018\ : std_logic;
signal \N__49017\ : std_logic;
signal \N__49016\ : std_logic;
signal \N__49015\ : std_logic;
signal \N__49014\ : std_logic;
signal \N__49011\ : std_logic;
signal \N__49008\ : std_logic;
signal \N__49005\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__49003\ : std_logic;
signal \N__49002\ : std_logic;
signal \N__49001\ : std_logic;
signal \N__49000\ : std_logic;
signal \N__48999\ : std_logic;
signal \N__48998\ : std_logic;
signal \N__48997\ : std_logic;
signal \N__48996\ : std_logic;
signal \N__48995\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48993\ : std_logic;
signal \N__48992\ : std_logic;
signal \N__48989\ : std_logic;
signal \N__48986\ : std_logic;
signal \N__48985\ : std_logic;
signal \N__48984\ : std_logic;
signal \N__48979\ : std_logic;
signal \N__48976\ : std_logic;
signal \N__48973\ : std_logic;
signal \N__48970\ : std_logic;
signal \N__48969\ : std_logic;
signal \N__48968\ : std_logic;
signal \N__48967\ : std_logic;
signal \N__48964\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48956\ : std_logic;
signal \N__48955\ : std_logic;
signal \N__48950\ : std_logic;
signal \N__48947\ : std_logic;
signal \N__48940\ : std_logic;
signal \N__48937\ : std_logic;
signal \N__48928\ : std_logic;
signal \N__48925\ : std_logic;
signal \N__48922\ : std_logic;
signal \N__48921\ : std_logic;
signal \N__48920\ : std_logic;
signal \N__48919\ : std_logic;
signal \N__48914\ : std_logic;
signal \N__48913\ : std_logic;
signal \N__48910\ : std_logic;
signal \N__48907\ : std_logic;
signal \N__48902\ : std_logic;
signal \N__48895\ : std_logic;
signal \N__48894\ : std_logic;
signal \N__48891\ : std_logic;
signal \N__48884\ : std_logic;
signal \N__48877\ : std_logic;
signal \N__48874\ : std_logic;
signal \N__48869\ : std_logic;
signal \N__48862\ : std_logic;
signal \N__48859\ : std_logic;
signal \N__48854\ : std_logic;
signal \N__48849\ : std_logic;
signal \N__48846\ : std_logic;
signal \N__48845\ : std_logic;
signal \N__48844\ : std_logic;
signal \N__48843\ : std_logic;
signal \N__48842\ : std_logic;
signal \N__48839\ : std_logic;
signal \N__48836\ : std_logic;
signal \N__48829\ : std_logic;
signal \N__48826\ : std_logic;
signal \N__48819\ : std_logic;
signal \N__48810\ : std_logic;
signal \N__48803\ : std_logic;
signal \N__48794\ : std_logic;
signal \N__48787\ : std_logic;
signal \N__48774\ : std_logic;
signal \N__48773\ : std_logic;
signal \N__48770\ : std_logic;
signal \N__48767\ : std_logic;
signal \N__48764\ : std_logic;
signal \N__48761\ : std_logic;
signal \N__48756\ : std_logic;
signal \N__48753\ : std_logic;
signal \N__48750\ : std_logic;
signal \N__48747\ : std_logic;
signal \N__48746\ : std_logic;
signal \N__48743\ : std_logic;
signal \N__48740\ : std_logic;
signal \N__48737\ : std_logic;
signal \N__48734\ : std_logic;
signal \N__48731\ : std_logic;
signal \N__48728\ : std_logic;
signal \N__48723\ : std_logic;
signal \N__48720\ : std_logic;
signal \N__48717\ : std_logic;
signal \N__48714\ : std_logic;
signal \N__48711\ : std_logic;
signal \N__48708\ : std_logic;
signal \N__48705\ : std_logic;
signal \N__48702\ : std_logic;
signal \N__48701\ : std_logic;
signal \N__48700\ : std_logic;
signal \N__48699\ : std_logic;
signal \N__48698\ : std_logic;
signal \N__48697\ : std_logic;
signal \N__48696\ : std_logic;
signal \N__48695\ : std_logic;
signal \N__48692\ : std_logic;
signal \N__48691\ : std_logic;
signal \N__48686\ : std_logic;
signal \N__48683\ : std_logic;
signal \N__48682\ : std_logic;
signal \N__48681\ : std_logic;
signal \N__48680\ : std_logic;
signal \N__48677\ : std_logic;
signal \N__48672\ : std_logic;
signal \N__48671\ : std_logic;
signal \N__48670\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48666\ : std_logic;
signal \N__48663\ : std_logic;
signal \N__48660\ : std_logic;
signal \N__48657\ : std_logic;
signal \N__48654\ : std_logic;
signal \N__48651\ : std_logic;
signal \N__48648\ : std_logic;
signal \N__48647\ : std_logic;
signal \N__48646\ : std_logic;
signal \N__48645\ : std_logic;
signal \N__48642\ : std_logic;
signal \N__48637\ : std_logic;
signal \N__48628\ : std_logic;
signal \N__48625\ : std_logic;
signal \N__48620\ : std_logic;
signal \N__48613\ : std_logic;
signal \N__48610\ : std_logic;
signal \N__48607\ : std_logic;
signal \N__48604\ : std_logic;
signal \N__48597\ : std_logic;
signal \N__48594\ : std_logic;
signal \N__48589\ : std_logic;
signal \N__48576\ : std_logic;
signal \N__48573\ : std_logic;
signal \N__48572\ : std_logic;
signal \N__48569\ : std_logic;
signal \N__48566\ : std_logic;
signal \N__48563\ : std_logic;
signal \N__48560\ : std_logic;
signal \N__48559\ : std_logic;
signal \N__48554\ : std_logic;
signal \N__48553\ : std_logic;
signal \N__48550\ : std_logic;
signal \N__48547\ : std_logic;
signal \N__48544\ : std_logic;
signal \N__48537\ : std_logic;
signal \N__48534\ : std_logic;
signal \N__48531\ : std_logic;
signal \N__48528\ : std_logic;
signal \N__48527\ : std_logic;
signal \N__48526\ : std_logic;
signal \N__48523\ : std_logic;
signal \N__48520\ : std_logic;
signal \N__48519\ : std_logic;
signal \N__48516\ : std_logic;
signal \N__48513\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48498\ : std_logic;
signal \N__48495\ : std_logic;
signal \N__48492\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48483\ : std_logic;
signal \N__48482\ : std_logic;
signal \N__48481\ : std_logic;
signal \N__48478\ : std_logic;
signal \N__48475\ : std_logic;
signal \N__48474\ : std_logic;
signal \N__48471\ : std_logic;
signal \N__48468\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48462\ : std_logic;
signal \N__48453\ : std_logic;
signal \N__48452\ : std_logic;
signal \N__48451\ : std_logic;
signal \N__48450\ : std_logic;
signal \N__48449\ : std_logic;
signal \N__48448\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48446\ : std_logic;
signal \N__48445\ : std_logic;
signal \N__48444\ : std_logic;
signal \N__48443\ : std_logic;
signal \N__48442\ : std_logic;
signal \N__48441\ : std_logic;
signal \N__48440\ : std_logic;
signal \N__48439\ : std_logic;
signal \N__48438\ : std_logic;
signal \N__48437\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48435\ : std_logic;
signal \N__48434\ : std_logic;
signal \N__48433\ : std_logic;
signal \N__48432\ : std_logic;
signal \N__48431\ : std_logic;
signal \N__48430\ : std_logic;
signal \N__48429\ : std_logic;
signal \N__48428\ : std_logic;
signal \N__48427\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48425\ : std_logic;
signal \N__48424\ : std_logic;
signal \N__48423\ : std_logic;
signal \N__48422\ : std_logic;
signal \N__48421\ : std_logic;
signal \N__48420\ : std_logic;
signal \N__48419\ : std_logic;
signal \N__48418\ : std_logic;
signal \N__48417\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48415\ : std_logic;
signal \N__48414\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48411\ : std_logic;
signal \N__48410\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48408\ : std_logic;
signal \N__48407\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48405\ : std_logic;
signal \N__48404\ : std_logic;
signal \N__48403\ : std_logic;
signal \N__48402\ : std_logic;
signal \N__48401\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48399\ : std_logic;
signal \N__48398\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48395\ : std_logic;
signal \N__48394\ : std_logic;
signal \N__48393\ : std_logic;
signal \N__48392\ : std_logic;
signal \N__48391\ : std_logic;
signal \N__48390\ : std_logic;
signal \N__48389\ : std_logic;
signal \N__48388\ : std_logic;
signal \N__48387\ : std_logic;
signal \N__48386\ : std_logic;
signal \N__48385\ : std_logic;
signal \N__48384\ : std_logic;
signal \N__48383\ : std_logic;
signal \N__48240\ : std_logic;
signal \N__48237\ : std_logic;
signal \N__48234\ : std_logic;
signal \N__48233\ : std_logic;
signal \N__48230\ : std_logic;
signal \N__48227\ : std_logic;
signal \N__48222\ : std_logic;
signal \N__48219\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48207\ : std_logic;
signal \N__48204\ : std_logic;
signal \N__48201\ : std_logic;
signal \N__48198\ : std_logic;
signal \N__48197\ : std_logic;
signal \N__48194\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48176\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48170\ : std_logic;
signal \N__48165\ : std_logic;
signal \N__48162\ : std_logic;
signal \N__48161\ : std_logic;
signal \N__48158\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48150\ : std_logic;
signal \N__48149\ : std_logic;
signal \N__48148\ : std_logic;
signal \N__48147\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48138\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48133\ : std_logic;
signal \N__48132\ : std_logic;
signal \N__48129\ : std_logic;
signal \N__48124\ : std_logic;
signal \N__48121\ : std_logic;
signal \N__48116\ : std_logic;
signal \N__48113\ : std_logic;
signal \N__48108\ : std_logic;
signal \N__48103\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48087\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48078\ : std_logic;
signal \N__48077\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48073\ : std_logic;
signal \N__48070\ : std_logic;
signal \N__48067\ : std_logic;
signal \N__48064\ : std_logic;
signal \N__48061\ : std_logic;
signal \N__48058\ : std_logic;
signal \N__48055\ : std_logic;
signal \N__48052\ : std_logic;
signal \N__48045\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48039\ : std_logic;
signal \N__48038\ : std_logic;
signal \N__48035\ : std_logic;
signal \N__48032\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48028\ : std_logic;
signal \N__48025\ : std_logic;
signal \N__48022\ : std_logic;
signal \N__48019\ : std_logic;
signal \N__48016\ : std_logic;
signal \N__48009\ : std_logic;
signal \N__48006\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__48000\ : std_logic;
signal \N__47997\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47995\ : std_logic;
signal \N__47994\ : std_logic;
signal \N__47993\ : std_logic;
signal \N__47992\ : std_logic;
signal \N__47991\ : std_logic;
signal \N__47988\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47981\ : std_logic;
signal \N__47978\ : std_logic;
signal \N__47975\ : std_logic;
signal \N__47970\ : std_logic;
signal \N__47967\ : std_logic;
signal \N__47964\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47958\ : std_logic;
signal \N__47955\ : std_logic;
signal \N__47950\ : std_logic;
signal \N__47945\ : std_logic;
signal \N__47940\ : std_logic;
signal \N__47935\ : std_logic;
signal \N__47928\ : std_logic;
signal \N__47927\ : std_logic;
signal \N__47924\ : std_logic;
signal \N__47921\ : std_logic;
signal \N__47918\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47912\ : std_logic;
signal \N__47909\ : std_logic;
signal \N__47906\ : std_logic;
signal \N__47903\ : std_logic;
signal \N__47900\ : std_logic;
signal \N__47897\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47883\ : std_logic;
signal \N__47882\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47869\ : std_logic;
signal \N__47866\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47857\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47843\ : std_logic;
signal \N__47840\ : std_logic;
signal \N__47839\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47820\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47808\ : std_logic;
signal \N__47805\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47798\ : std_logic;
signal \N__47797\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47792\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47780\ : std_logic;
signal \N__47779\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47770\ : std_logic;
signal \N__47767\ : std_logic;
signal \N__47760\ : std_logic;
signal \N__47757\ : std_logic;
signal \N__47754\ : std_logic;
signal \N__47749\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47738\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47727\ : std_logic;
signal \N__47724\ : std_logic;
signal \N__47721\ : std_logic;
signal \N__47718\ : std_logic;
signal \N__47715\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47711\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47707\ : std_logic;
signal \N__47704\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47698\ : std_logic;
signal \N__47695\ : std_logic;
signal \N__47692\ : std_logic;
signal \N__47685\ : std_logic;
signal \N__47682\ : std_logic;
signal \N__47679\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47675\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47658\ : std_logic;
signal \N__47655\ : std_logic;
signal \N__47654\ : std_logic;
signal \N__47651\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47643\ : std_logic;
signal \N__47640\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47630\ : std_logic;
signal \N__47627\ : std_logic;
signal \N__47624\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47617\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47609\ : std_logic;
signal \N__47604\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47597\ : std_logic;
signal \N__47594\ : std_logic;
signal \N__47591\ : std_logic;
signal \N__47586\ : std_logic;
signal \N__47583\ : std_logic;
signal \N__47582\ : std_logic;
signal \N__47579\ : std_logic;
signal \N__47576\ : std_logic;
signal \N__47571\ : std_logic;
signal \N__47570\ : std_logic;
signal \N__47567\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47561\ : std_logic;
signal \N__47556\ : std_logic;
signal \N__47553\ : std_logic;
signal \N__47550\ : std_logic;
signal \N__47549\ : std_logic;
signal \N__47546\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47538\ : std_logic;
signal \N__47535\ : std_logic;
signal \N__47534\ : std_logic;
signal \N__47531\ : std_logic;
signal \N__47530\ : std_logic;
signal \N__47529\ : std_logic;
signal \N__47528\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47526\ : std_logic;
signal \N__47525\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47523\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47519\ : std_logic;
signal \N__47518\ : std_logic;
signal \N__47515\ : std_logic;
signal \N__47512\ : std_logic;
signal \N__47507\ : std_logic;
signal \N__47506\ : std_logic;
signal \N__47505\ : std_logic;
signal \N__47504\ : std_logic;
signal \N__47503\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47501\ : std_logic;
signal \N__47498\ : std_logic;
signal \N__47497\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47495\ : std_logic;
signal \N__47494\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47487\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47476\ : std_logic;
signal \N__47473\ : std_logic;
signal \N__47468\ : std_logic;
signal \N__47465\ : std_logic;
signal \N__47462\ : std_logic;
signal \N__47459\ : std_logic;
signal \N__47458\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47445\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47432\ : std_logic;
signal \N__47423\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47416\ : std_logic;
signal \N__47409\ : std_logic;
signal \N__47406\ : std_logic;
signal \N__47403\ : std_logic;
signal \N__47398\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47390\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47382\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47374\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47359\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47331\ : std_logic;
signal \N__47328\ : std_logic;
signal \N__47325\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47317\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47305\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47294\ : std_logic;
signal \N__47291\ : std_logic;
signal \N__47290\ : std_logic;
signal \N__47287\ : std_logic;
signal \N__47284\ : std_logic;
signal \N__47281\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47265\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47263\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47252\ : std_logic;
signal \N__47249\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47238\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47236\ : std_logic;
signal \N__47235\ : std_logic;
signal \N__47232\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47230\ : std_logic;
signal \N__47229\ : std_logic;
signal \N__47226\ : std_logic;
signal \N__47225\ : std_logic;
signal \N__47220\ : std_logic;
signal \N__47217\ : std_logic;
signal \N__47212\ : std_logic;
signal \N__47209\ : std_logic;
signal \N__47206\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47200\ : std_logic;
signal \N__47197\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47181\ : std_logic;
signal \N__47180\ : std_logic;
signal \N__47177\ : std_logic;
signal \N__47176\ : std_logic;
signal \N__47173\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47169\ : std_logic;
signal \N__47168\ : std_logic;
signal \N__47165\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47157\ : std_logic;
signal \N__47156\ : std_logic;
signal \N__47153\ : std_logic;
signal \N__47148\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47129\ : std_logic;
signal \N__47126\ : std_logic;
signal \N__47115\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47109\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47105\ : std_logic;
signal \N__47102\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47096\ : std_logic;
signal \N__47093\ : std_logic;
signal \N__47088\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47084\ : std_logic;
signal \N__47081\ : std_logic;
signal \N__47078\ : std_logic;
signal \N__47075\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47066\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47060\ : std_logic;
signal \N__47057\ : std_logic;
signal \N__47054\ : std_logic;
signal \N__47051\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47043\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47031\ : std_logic;
signal \N__47028\ : std_logic;
signal \N__47025\ : std_logic;
signal \N__47022\ : std_logic;
signal \N__47019\ : std_logic;
signal \N__47016\ : std_logic;
signal \N__47015\ : std_logic;
signal \N__47012\ : std_logic;
signal \N__47009\ : std_logic;
signal \N__47006\ : std_logic;
signal \N__47003\ : std_logic;
signal \N__46998\ : std_logic;
signal \N__46995\ : std_logic;
signal \N__46992\ : std_logic;
signal \N__46989\ : std_logic;
signal \N__46986\ : std_logic;
signal \N__46983\ : std_logic;
signal \N__46980\ : std_logic;
signal \N__46979\ : std_logic;
signal \N__46978\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46965\ : std_logic;
signal \N__46964\ : std_logic;
signal \N__46963\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46958\ : std_logic;
signal \N__46955\ : std_logic;
signal \N__46950\ : std_logic;
signal \N__46945\ : std_logic;
signal \N__46944\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46941\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46932\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46930\ : std_logic;
signal \N__46929\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46927\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46895\ : std_logic;
signal \N__46890\ : std_logic;
signal \N__46887\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46883\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46872\ : std_logic;
signal \N__46871\ : std_logic;
signal \N__46868\ : std_logic;
signal \N__46865\ : std_logic;
signal \N__46862\ : std_logic;
signal \N__46859\ : std_logic;
signal \N__46856\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46841\ : std_logic;
signal \N__46826\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46801\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46787\ : std_logic;
signal \N__46786\ : std_logic;
signal \N__46783\ : std_logic;
signal \N__46778\ : std_logic;
signal \N__46777\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46775\ : std_logic;
signal \N__46774\ : std_logic;
signal \N__46769\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46763\ : std_logic;
signal \N__46758\ : std_logic;
signal \N__46755\ : std_logic;
signal \N__46746\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46744\ : std_logic;
signal \N__46743\ : std_logic;
signal \N__46740\ : std_logic;
signal \N__46737\ : std_logic;
signal \N__46734\ : std_logic;
signal \N__46729\ : std_logic;
signal \N__46726\ : std_logic;
signal \N__46723\ : std_logic;
signal \N__46722\ : std_logic;
signal \N__46719\ : std_logic;
signal \N__46716\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46710\ : std_logic;
signal \N__46705\ : std_logic;
signal \N__46702\ : std_logic;
signal \N__46695\ : std_logic;
signal \N__46692\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46688\ : std_logic;
signal \N__46687\ : std_logic;
signal \N__46684\ : std_logic;
signal \N__46683\ : std_logic;
signal \N__46680\ : std_logic;
signal \N__46679\ : std_logic;
signal \N__46678\ : std_logic;
signal \N__46677\ : std_logic;
signal \N__46674\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46670\ : std_logic;
signal \N__46669\ : std_logic;
signal \N__46666\ : std_logic;
signal \N__46663\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46657\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46642\ : std_logic;
signal \N__46639\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46631\ : std_logic;
signal \N__46626\ : std_logic;
signal \N__46621\ : std_logic;
signal \N__46618\ : std_logic;
signal \N__46613\ : std_logic;
signal \N__46602\ : std_logic;
signal \N__46599\ : std_logic;
signal \N__46596\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46592\ : std_logic;
signal \N__46589\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46581\ : std_logic;
signal \N__46580\ : std_logic;
signal \N__46579\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46571\ : std_logic;
signal \N__46570\ : std_logic;
signal \N__46569\ : std_logic;
signal \N__46568\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46561\ : std_logic;
signal \N__46552\ : std_logic;
signal \N__46549\ : std_logic;
signal \N__46542\ : std_logic;
signal \N__46539\ : std_logic;
signal \N__46536\ : std_logic;
signal \N__46535\ : std_logic;
signal \N__46534\ : std_logic;
signal \N__46531\ : std_logic;
signal \N__46530\ : std_logic;
signal \N__46529\ : std_logic;
signal \N__46528\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46524\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46519\ : std_logic;
signal \N__46518\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46516\ : std_logic;
signal \N__46515\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46506\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46495\ : std_logic;
signal \N__46492\ : std_logic;
signal \N__46489\ : std_logic;
signal \N__46488\ : std_logic;
signal \N__46487\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46483\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46481\ : std_logic;
signal \N__46476\ : std_logic;
signal \N__46475\ : std_logic;
signal \N__46472\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46464\ : std_logic;
signal \N__46457\ : std_logic;
signal \N__46452\ : std_logic;
signal \N__46451\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46449\ : std_logic;
signal \N__46448\ : std_logic;
signal \N__46445\ : std_logic;
signal \N__46442\ : std_logic;
signal \N__46439\ : std_logic;
signal \N__46436\ : std_logic;
signal \N__46431\ : std_logic;
signal \N__46428\ : std_logic;
signal \N__46425\ : std_logic;
signal \N__46422\ : std_logic;
signal \N__46417\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46411\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46401\ : std_logic;
signal \N__46396\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46381\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46371\ : std_logic;
signal \N__46356\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46346\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46338\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46326\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46317\ : std_logic;
signal \N__46314\ : std_logic;
signal \N__46311\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46305\ : std_logic;
signal \N__46302\ : std_logic;
signal \N__46299\ : std_logic;
signal \N__46296\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46290\ : std_logic;
signal \N__46287\ : std_logic;
signal \N__46284\ : std_logic;
signal \N__46281\ : std_logic;
signal \N__46278\ : std_logic;
signal \N__46275\ : std_logic;
signal \N__46274\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46268\ : std_logic;
signal \N__46265\ : std_logic;
signal \N__46260\ : std_logic;
signal \N__46257\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46250\ : std_logic;
signal \N__46247\ : std_logic;
signal \N__46242\ : std_logic;
signal \N__46239\ : std_logic;
signal \N__46238\ : std_logic;
signal \N__46235\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46229\ : std_logic;
signal \N__46226\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46218\ : std_logic;
signal \N__46217\ : std_logic;
signal \N__46216\ : std_logic;
signal \N__46211\ : std_logic;
signal \N__46208\ : std_logic;
signal \N__46203\ : std_logic;
signal \N__46200\ : std_logic;
signal \N__46197\ : std_logic;
signal \N__46194\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46188\ : std_logic;
signal \N__46185\ : std_logic;
signal \N__46182\ : std_logic;
signal \N__46179\ : std_logic;
signal \N__46176\ : std_logic;
signal \N__46173\ : std_logic;
signal \N__46170\ : std_logic;
signal \N__46167\ : std_logic;
signal \N__46164\ : std_logic;
signal \N__46161\ : std_logic;
signal \N__46158\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46137\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46131\ : std_logic;
signal \N__46128\ : std_logic;
signal \N__46125\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46110\ : std_logic;
signal \N__46107\ : std_logic;
signal \N__46104\ : std_logic;
signal \N__46101\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46092\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46068\ : std_logic;
signal \N__46065\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46046\ : std_logic;
signal \N__46043\ : std_logic;
signal \N__46040\ : std_logic;
signal \N__46039\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46033\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__46001\ : std_logic;
signal \N__45998\ : std_logic;
signal \N__45995\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45984\ : std_logic;
signal \N__45981\ : std_logic;
signal \N__45978\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45972\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45960\ : std_logic;
signal \N__45957\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45951\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45939\ : std_logic;
signal \N__45938\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45934\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45928\ : std_logic;
signal \N__45925\ : std_logic;
signal \N__45918\ : std_logic;
signal \N__45915\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45909\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45894\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45890\ : std_logic;
signal \N__45887\ : std_logic;
signal \N__45886\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45880\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45867\ : std_logic;
signal \N__45864\ : std_logic;
signal \N__45861\ : std_logic;
signal \N__45858\ : std_logic;
signal \N__45855\ : std_logic;
signal \N__45852\ : std_logic;
signal \N__45849\ : std_logic;
signal \N__45848\ : std_logic;
signal \N__45845\ : std_logic;
signal \N__45842\ : std_logic;
signal \N__45839\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45828\ : std_logic;
signal \N__45825\ : std_logic;
signal \N__45822\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45816\ : std_logic;
signal \N__45813\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45806\ : std_logic;
signal \N__45805\ : std_logic;
signal \N__45802\ : std_logic;
signal \N__45799\ : std_logic;
signal \N__45796\ : std_logic;
signal \N__45793\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45784\ : std_logic;
signal \N__45777\ : std_logic;
signal \N__45774\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45764\ : std_logic;
signal \N__45763\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45761\ : std_logic;
signal \N__45760\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45758\ : std_logic;
signal \N__45757\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45755\ : std_logic;
signal \N__45754\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45751\ : std_logic;
signal \N__45750\ : std_logic;
signal \N__45749\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45747\ : std_logic;
signal \N__45746\ : std_logic;
signal \N__45745\ : std_logic;
signal \N__45744\ : std_logic;
signal \N__45743\ : std_logic;
signal \N__45742\ : std_logic;
signal \N__45741\ : std_logic;
signal \N__45740\ : std_logic;
signal \N__45739\ : std_logic;
signal \N__45738\ : std_logic;
signal \N__45737\ : std_logic;
signal \N__45734\ : std_logic;
signal \N__45733\ : std_logic;
signal \N__45732\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45730\ : std_logic;
signal \N__45729\ : std_logic;
signal \N__45728\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45721\ : std_logic;
signal \N__45720\ : std_logic;
signal \N__45717\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45704\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45700\ : std_logic;
signal \N__45699\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45697\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45694\ : std_logic;
signal \N__45693\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45691\ : std_logic;
signal \N__45690\ : std_logic;
signal \N__45689\ : std_logic;
signal \N__45688\ : std_logic;
signal \N__45687\ : std_logic;
signal \N__45686\ : std_logic;
signal \N__45685\ : std_logic;
signal \N__45684\ : std_logic;
signal \N__45681\ : std_logic;
signal \N__45680\ : std_logic;
signal \N__45679\ : std_logic;
signal \N__45678\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45676\ : std_logic;
signal \N__45673\ : std_logic;
signal \N__45672\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45670\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45666\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45661\ : std_logic;
signal \N__45660\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45658\ : std_logic;
signal \N__45657\ : std_logic;
signal \N__45656\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45649\ : std_logic;
signal \N__45648\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45646\ : std_logic;
signal \N__45645\ : std_logic;
signal \N__45644\ : std_logic;
signal \N__45643\ : std_logic;
signal \N__45642\ : std_logic;
signal \N__45639\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45635\ : std_logic;
signal \N__45634\ : std_logic;
signal \N__45633\ : std_logic;
signal \N__45632\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45630\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45628\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45625\ : std_logic;
signal \N__45616\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45589\ : std_logic;
signal \N__45588\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45586\ : std_logic;
signal \N__45585\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45581\ : std_logic;
signal \N__45580\ : std_logic;
signal \N__45579\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45576\ : std_logic;
signal \N__45573\ : std_logic;
signal \N__45572\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45569\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45566\ : std_logic;
signal \N__45565\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45563\ : std_logic;
signal \N__45562\ : std_logic;
signal \N__45559\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45556\ : std_logic;
signal \N__45555\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45553\ : std_logic;
signal \N__45552\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45550\ : std_logic;
signal \N__45549\ : std_logic;
signal \N__45548\ : std_logic;
signal \N__45547\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45542\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45539\ : std_logic;
signal \N__45536\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45532\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45506\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45503\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45497\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45486\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45470\ : std_logic;
signal \N__45463\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45452\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45450\ : std_logic;
signal \N__45449\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45447\ : std_logic;
signal \N__45446\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45442\ : std_logic;
signal \N__45441\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45438\ : std_logic;
signal \N__45437\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45435\ : std_logic;
signal \N__45434\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45432\ : std_logic;
signal \N__45423\ : std_logic;
signal \N__45418\ : std_logic;
signal \N__45417\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45413\ : std_logic;
signal \N__45412\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45402\ : std_logic;
signal \N__45401\ : std_logic;
signal \N__45400\ : std_logic;
signal \N__45399\ : std_logic;
signal \N__45396\ : std_logic;
signal \N__45395\ : std_logic;
signal \N__45394\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45392\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45386\ : std_logic;
signal \N__45375\ : std_logic;
signal \N__45368\ : std_logic;
signal \N__45357\ : std_logic;
signal \N__45348\ : std_logic;
signal \N__45339\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45326\ : std_logic;
signal \N__45325\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45323\ : std_logic;
signal \N__45322\ : std_logic;
signal \N__45319\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45317\ : std_logic;
signal \N__45314\ : std_logic;
signal \N__45313\ : std_logic;
signal \N__45312\ : std_logic;
signal \N__45311\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45309\ : std_logic;
signal \N__45308\ : std_logic;
signal \N__45307\ : std_logic;
signal \N__45304\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45298\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45296\ : std_logic;
signal \N__45293\ : std_logic;
signal \N__45292\ : std_logic;
signal \N__45289\ : std_logic;
signal \N__45286\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45283\ : std_logic;
signal \N__45282\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45276\ : std_logic;
signal \N__45269\ : std_logic;
signal \N__45262\ : std_logic;
signal \N__45251\ : std_logic;
signal \N__45244\ : std_logic;
signal \N__45239\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45227\ : std_logic;
signal \N__45224\ : std_logic;
signal \N__45223\ : std_logic;
signal \N__45220\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45218\ : std_logic;
signal \N__45211\ : std_logic;
signal \N__45206\ : std_logic;
signal \N__45197\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45183\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45163\ : std_logic;
signal \N__45152\ : std_logic;
signal \N__45145\ : std_logic;
signal \N__45142\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45140\ : std_logic;
signal \N__45139\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45137\ : std_logic;
signal \N__45136\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45105\ : std_logic;
signal \N__45104\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45100\ : std_logic;
signal \N__45099\ : std_logic;
signal \N__45098\ : std_logic;
signal \N__45097\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45095\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45093\ : std_logic;
signal \N__45092\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45082\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45074\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45053\ : std_logic;
signal \N__45046\ : std_logic;
signal \N__45037\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45030\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45027\ : std_logic;
signal \N__45026\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45024\ : std_logic;
signal \N__45023\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45018\ : std_logic;
signal \N__45017\ : std_logic;
signal \N__45016\ : std_logic;
signal \N__45007\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__44999\ : std_logic;
signal \N__44990\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44962\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44958\ : std_logic;
signal \N__44957\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44955\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44941\ : std_logic;
signal \N__44938\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44936\ : std_logic;
signal \N__44935\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44933\ : std_logic;
signal \N__44932\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44930\ : std_logic;
signal \N__44929\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44927\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44924\ : std_logic;
signal \N__44923\ : std_logic;
signal \N__44918\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44900\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44872\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44870\ : std_logic;
signal \N__44869\ : std_logic;
signal \N__44864\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44861\ : std_logic;
signal \N__44860\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44856\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44844\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44833\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44829\ : std_logic;
signal \N__44828\ : std_logic;
signal \N__44823\ : std_logic;
signal \N__44812\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44794\ : std_logic;
signal \N__44791\ : std_logic;
signal \N__44774\ : std_logic;
signal \N__44771\ : std_logic;
signal \N__44762\ : std_logic;
signal \N__44753\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44743\ : std_logic;
signal \N__44740\ : std_logic;
signal \N__44737\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44723\ : std_logic;
signal \N__44722\ : std_logic;
signal \N__44719\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44717\ : std_logic;
signal \N__44716\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44714\ : std_logic;
signal \N__44711\ : std_logic;
signal \N__44710\ : std_logic;
signal \N__44707\ : std_logic;
signal \N__44706\ : std_logic;
signal \N__44699\ : std_logic;
signal \N__44692\ : std_logic;
signal \N__44685\ : std_logic;
signal \N__44678\ : std_logic;
signal \N__44671\ : std_logic;
signal \N__44670\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44666\ : std_logic;
signal \N__44665\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44645\ : std_logic;
signal \N__44644\ : std_logic;
signal \N__44637\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44635\ : std_logic;
signal \N__44634\ : std_logic;
signal \N__44633\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44631\ : std_logic;
signal \N__44630\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44618\ : std_logic;
signal \N__44611\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44601\ : std_logic;
signal \N__44600\ : std_logic;
signal \N__44597\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44589\ : std_logic;
signal \N__44582\ : std_logic;
signal \N__44575\ : std_logic;
signal \N__44568\ : std_logic;
signal \N__44561\ : std_logic;
signal \N__44554\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44538\ : std_logic;
signal \N__44531\ : std_logic;
signal \N__44528\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44522\ : std_logic;
signal \N__44521\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44519\ : std_logic;
signal \N__44518\ : std_logic;
signal \N__44513\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44507\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44487\ : std_logic;
signal \N__44486\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44484\ : std_logic;
signal \N__44483\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44463\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44441\ : std_logic;
signal \N__44440\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44436\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44434\ : std_logic;
signal \N__44433\ : std_logic;
signal \N__44426\ : std_logic;
signal \N__44419\ : std_logic;
signal \N__44416\ : std_logic;
signal \N__44407\ : std_logic;
signal \N__44398\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44386\ : std_logic;
signal \N__44385\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44360\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44332\ : std_logic;
signal \N__44325\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44313\ : std_logic;
signal \N__44308\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44281\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44265\ : std_logic;
signal \N__44258\ : std_logic;
signal \N__44251\ : std_logic;
signal \N__44248\ : std_logic;
signal \N__44245\ : std_logic;
signal \N__44240\ : std_logic;
signal \N__44237\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44221\ : std_logic;
signal \N__44208\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44186\ : std_logic;
signal \N__44183\ : std_logic;
signal \N__44176\ : std_logic;
signal \N__44173\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44147\ : std_logic;
signal \N__44144\ : std_logic;
signal \N__44141\ : std_logic;
signal \N__44138\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44130\ : std_logic;
signal \N__44129\ : std_logic;
signal \N__44128\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44122\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44117\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44114\ : std_logic;
signal \N__44113\ : std_logic;
signal \N__44110\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44106\ : std_logic;
signal \N__44103\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44098\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44090\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44070\ : std_logic;
signal \N__44067\ : std_logic;
signal \N__44064\ : std_logic;
signal \N__44061\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44038\ : std_logic;
signal \N__44035\ : std_logic;
signal \N__44026\ : std_logic;
signal \N__44013\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44006\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43992\ : std_logic;
signal \N__43989\ : std_logic;
signal \N__43986\ : std_logic;
signal \N__43985\ : std_logic;
signal \N__43982\ : std_logic;
signal \N__43979\ : std_logic;
signal \N__43976\ : std_logic;
signal \N__43975\ : std_logic;
signal \N__43972\ : std_logic;
signal \N__43969\ : std_logic;
signal \N__43966\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43950\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43941\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43937\ : std_logic;
signal \N__43936\ : std_logic;
signal \N__43933\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43917\ : std_logic;
signal \N__43914\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43905\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43895\ : std_logic;
signal \N__43894\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43885\ : std_logic;
signal \N__43882\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43860\ : std_logic;
signal \N__43857\ : std_logic;
signal \N__43854\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43849\ : std_logic;
signal \N__43846\ : std_logic;
signal \N__43843\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43830\ : std_logic;
signal \N__43827\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43812\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43810\ : std_logic;
signal \N__43807\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43798\ : std_logic;
signal \N__43795\ : std_logic;
signal \N__43792\ : std_logic;
signal \N__43785\ : std_logic;
signal \N__43782\ : std_logic;
signal \N__43779\ : std_logic;
signal \N__43776\ : std_logic;
signal \N__43773\ : std_logic;
signal \N__43770\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43766\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43760\ : std_logic;
signal \N__43757\ : std_logic;
signal \N__43752\ : std_logic;
signal \N__43749\ : std_logic;
signal \N__43746\ : std_logic;
signal \N__43743\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43737\ : std_logic;
signal \N__43734\ : std_logic;
signal \N__43733\ : std_logic;
signal \N__43730\ : std_logic;
signal \N__43727\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43698\ : std_logic;
signal \N__43695\ : std_logic;
signal \N__43692\ : std_logic;
signal \N__43689\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43685\ : std_logic;
signal \N__43682\ : std_logic;
signal \N__43679\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43671\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43667\ : std_logic;
signal \N__43664\ : std_logic;
signal \N__43663\ : std_logic;
signal \N__43660\ : std_logic;
signal \N__43657\ : std_logic;
signal \N__43654\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43641\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43632\ : std_logic;
signal \N__43629\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43623\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43615\ : std_logic;
signal \N__43612\ : std_logic;
signal \N__43609\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43599\ : std_logic;
signal \N__43596\ : std_logic;
signal \N__43595\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43568\ : std_logic;
signal \N__43567\ : std_logic;
signal \N__43564\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43558\ : std_logic;
signal \N__43555\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43548\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43540\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43530\ : std_logic;
signal \N__43527\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43509\ : std_logic;
signal \N__43506\ : std_logic;
signal \N__43503\ : std_logic;
signal \N__43500\ : std_logic;
signal \N__43497\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43490\ : std_logic;
signal \N__43487\ : std_logic;
signal \N__43486\ : std_logic;
signal \N__43483\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43477\ : std_logic;
signal \N__43470\ : std_logic;
signal \N__43467\ : std_logic;
signal \N__43464\ : std_logic;
signal \N__43461\ : std_logic;
signal \N__43458\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43451\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43447\ : std_logic;
signal \N__43444\ : std_logic;
signal \N__43441\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43432\ : std_logic;
signal \N__43425\ : std_logic;
signal \N__43422\ : std_logic;
signal \N__43419\ : std_logic;
signal \N__43416\ : std_logic;
signal \N__43413\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43400\ : std_logic;
signal \N__43399\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43393\ : std_logic;
signal \N__43390\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43380\ : std_logic;
signal \N__43377\ : std_logic;
signal \N__43374\ : std_logic;
signal \N__43371\ : std_logic;
signal \N__43370\ : std_logic;
signal \N__43369\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43361\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43353\ : std_logic;
signal \N__43350\ : std_logic;
signal \N__43347\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43338\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43332\ : std_logic;
signal \N__43329\ : std_logic;
signal \N__43326\ : std_logic;
signal \N__43323\ : std_logic;
signal \N__43320\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43315\ : std_logic;
signal \N__43312\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43304\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43295\ : std_logic;
signal \N__43294\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43289\ : std_logic;
signal \N__43286\ : std_logic;
signal \N__43283\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43269\ : std_logic;
signal \N__43266\ : std_logic;
signal \N__43259\ : std_logic;
signal \N__43256\ : std_logic;
signal \N__43251\ : std_logic;
signal \N__43250\ : std_logic;
signal \N__43245\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43232\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43228\ : std_logic;
signal \N__43225\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43213\ : std_logic;
signal \N__43210\ : std_logic;
signal \N__43207\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43198\ : std_logic;
signal \N__43195\ : std_logic;
signal \N__43192\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43175\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43167\ : std_logic;
signal \N__43164\ : std_logic;
signal \N__43161\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43159\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43137\ : std_logic;
signal \N__43132\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43116\ : std_logic;
signal \N__43113\ : std_logic;
signal \N__43110\ : std_logic;
signal \N__43107\ : std_logic;
signal \N__43104\ : std_logic;
signal \N__43101\ : std_logic;
signal \N__43098\ : std_logic;
signal \N__43095\ : std_logic;
signal \N__43092\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43086\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43084\ : std_logic;
signal \N__43081\ : std_logic;
signal \N__43078\ : std_logic;
signal \N__43075\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43065\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43052\ : std_logic;
signal \N__43049\ : std_logic;
signal \N__43048\ : std_logic;
signal \N__43045\ : std_logic;
signal \N__43042\ : std_logic;
signal \N__43039\ : std_logic;
signal \N__43036\ : std_logic;
signal \N__43029\ : std_logic;
signal \N__43026\ : std_logic;
signal \N__43023\ : std_logic;
signal \N__43020\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43014\ : std_logic;
signal \N__43011\ : std_logic;
signal \N__43008\ : std_logic;
signal \N__43005\ : std_logic;
signal \N__43002\ : std_logic;
signal \N__42999\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42991\ : std_logic;
signal \N__42988\ : std_logic;
signal \N__42983\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42975\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42973\ : std_logic;
signal \N__42972\ : std_logic;
signal \N__42969\ : std_logic;
signal \N__42966\ : std_logic;
signal \N__42963\ : std_logic;
signal \N__42960\ : std_logic;
signal \N__42955\ : std_logic;
signal \N__42948\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42942\ : std_logic;
signal \N__42939\ : std_logic;
signal \N__42936\ : std_logic;
signal \N__42933\ : std_logic;
signal \N__42930\ : std_logic;
signal \N__42927\ : std_logic;
signal \N__42924\ : std_logic;
signal \N__42921\ : std_logic;
signal \N__42918\ : std_logic;
signal \N__42915\ : std_logic;
signal \N__42912\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42903\ : std_logic;
signal \N__42900\ : std_logic;
signal \N__42899\ : std_logic;
signal \N__42898\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42883\ : std_logic;
signal \N__42880\ : std_logic;
signal \N__42877\ : std_logic;
signal \N__42872\ : std_logic;
signal \N__42867\ : std_logic;
signal \N__42864\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42857\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42847\ : std_logic;
signal \N__42844\ : std_logic;
signal \N__42841\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42831\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42824\ : std_logic;
signal \N__42821\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42801\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42776\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42767\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42756\ : std_logic;
signal \N__42753\ : std_logic;
signal \N__42750\ : std_logic;
signal \N__42747\ : std_logic;
signal \N__42742\ : std_logic;
signal \N__42735\ : std_logic;
signal \N__42732\ : std_logic;
signal \N__42729\ : std_logic;
signal \N__42726\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42722\ : std_logic;
signal \N__42719\ : std_logic;
signal \N__42716\ : std_logic;
signal \N__42715\ : std_logic;
signal \N__42712\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42703\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42701\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42693\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42676\ : std_logic;
signal \N__42673\ : std_logic;
signal \N__42666\ : std_logic;
signal \N__42665\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42651\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42642\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42634\ : std_logic;
signal \N__42633\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42626\ : std_logic;
signal \N__42625\ : std_logic;
signal \N__42622\ : std_logic;
signal \N__42619\ : std_logic;
signal \N__42614\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42609\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42597\ : std_logic;
signal \N__42594\ : std_logic;
signal \N__42589\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42572\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42542\ : std_logic;
signal \N__42539\ : std_logic;
signal \N__42538\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42532\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42501\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42494\ : std_logic;
signal \N__42491\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42455\ : std_logic;
signal \N__42454\ : std_logic;
signal \N__42451\ : std_logic;
signal \N__42448\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42425\ : std_logic;
signal \N__42422\ : std_logic;
signal \N__42419\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42411\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42401\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42397\ : std_logic;
signal \N__42392\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42386\ : std_logic;
signal \N__42383\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42348\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42326\ : std_logic;
signal \N__42325\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42321\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42303\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42278\ : std_logic;
signal \N__42275\ : std_logic;
signal \N__42270\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42264\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42261\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42257\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42246\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42210\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42208\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42202\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42186\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42173\ : std_logic;
signal \N__42170\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42164\ : std_logic;
signal \N__42161\ : std_logic;
signal \N__42156\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42150\ : std_logic;
signal \N__42147\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42141\ : std_logic;
signal \N__42138\ : std_logic;
signal \N__42135\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42124\ : std_logic;
signal \N__42121\ : std_logic;
signal \N__42118\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42110\ : std_logic;
signal \N__42107\ : std_logic;
signal \N__42104\ : std_logic;
signal \N__42099\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42080\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42071\ : std_logic;
signal \N__42068\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42056\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42052\ : std_logic;
signal \N__42049\ : std_logic;
signal \N__42046\ : std_logic;
signal \N__42043\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42035\ : std_logic;
signal \N__42030\ : std_logic;
signal \N__42027\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42020\ : std_logic;
signal \N__42017\ : std_logic;
signal \N__42014\ : std_logic;
signal \N__42013\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41996\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41988\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41981\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41977\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41974\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41969\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41957\ : std_logic;
signal \N__41954\ : std_logic;
signal \N__41953\ : std_logic;
signal \N__41950\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41948\ : std_logic;
signal \N__41945\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41933\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41929\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41923\ : std_logic;
signal \N__41920\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41882\ : std_logic;
signal \N__41881\ : std_logic;
signal \N__41878\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41860\ : std_logic;
signal \N__41857\ : std_logic;
signal \N__41852\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41843\ : std_logic;
signal \N__41840\ : std_logic;
signal \N__41837\ : std_logic;
signal \N__41834\ : std_logic;
signal \N__41829\ : std_logic;
signal \N__41826\ : std_logic;
signal \N__41823\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41814\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41804\ : std_logic;
signal \N__41801\ : std_logic;
signal \N__41798\ : std_logic;
signal \N__41795\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41787\ : std_logic;
signal \N__41784\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41769\ : std_logic;
signal \N__41766\ : std_logic;
signal \N__41765\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41761\ : std_logic;
signal \N__41756\ : std_logic;
signal \N__41753\ : std_logic;
signal \N__41748\ : std_logic;
signal \N__41745\ : std_logic;
signal \N__41742\ : std_logic;
signal \N__41739\ : std_logic;
signal \N__41736\ : std_logic;
signal \N__41733\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41724\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41719\ : std_logic;
signal \N__41714\ : std_logic;
signal \N__41711\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41703\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41694\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41676\ : std_logic;
signal \N__41673\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41669\ : std_logic;
signal \N__41666\ : std_logic;
signal \N__41665\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41663\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41660\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41654\ : std_logic;
signal \N__41653\ : std_logic;
signal \N__41650\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41644\ : std_logic;
signal \N__41641\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41637\ : std_logic;
signal \N__41636\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41632\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41626\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41612\ : std_logic;
signal \N__41611\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41600\ : std_logic;
signal \N__41599\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41594\ : std_logic;
signal \N__41593\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41585\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41577\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41561\ : std_logic;
signal \N__41558\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41534\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41528\ : std_logic;
signal \N__41525\ : std_logic;
signal \N__41522\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41513\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41507\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41492\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41478\ : std_logic;
signal \N__41477\ : std_logic;
signal \N__41474\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41468\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41459\ : std_logic;
signal \N__41456\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41442\ : std_logic;
signal \N__41439\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41424\ : std_logic;
signal \N__41423\ : std_logic;
signal \N__41422\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41416\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41404\ : std_logic;
signal \N__41401\ : std_logic;
signal \N__41394\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41388\ : std_logic;
signal \N__41385\ : std_logic;
signal \N__41382\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41362\ : std_logic;
signal \N__41359\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41346\ : std_logic;
signal \N__41343\ : std_logic;
signal \N__41340\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41334\ : std_logic;
signal \N__41331\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41325\ : std_logic;
signal \N__41322\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41316\ : std_logic;
signal \N__41313\ : std_logic;
signal \N__41310\ : std_logic;
signal \N__41307\ : std_logic;
signal \N__41304\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41295\ : std_logic;
signal \N__41292\ : std_logic;
signal \N__41289\ : std_logic;
signal \N__41286\ : std_logic;
signal \N__41283\ : std_logic;
signal \N__41280\ : std_logic;
signal \N__41279\ : std_logic;
signal \N__41276\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41255\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41238\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41226\ : std_logic;
signal \N__41223\ : std_logic;
signal \N__41220\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41200\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41194\ : std_logic;
signal \N__41191\ : std_logic;
signal \N__41188\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41179\ : std_logic;
signal \N__41176\ : std_logic;
signal \N__41173\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41154\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41147\ : std_logic;
signal \N__41146\ : std_logic;
signal \N__41143\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41137\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41118\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41109\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41092\ : std_logic;
signal \N__41085\ : std_logic;
signal \N__41082\ : std_logic;
signal \N__41079\ : std_logic;
signal \N__41076\ : std_logic;
signal \N__41073\ : std_logic;
signal \N__41070\ : std_logic;
signal \N__41067\ : std_logic;
signal \N__41064\ : std_logic;
signal \N__41061\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41059\ : std_logic;
signal \N__41056\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41047\ : std_logic;
signal \N__41044\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41036\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41016\ : std_logic;
signal \N__41013\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41006\ : std_logic;
signal \N__41003\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40989\ : std_logic;
signal \N__40986\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40976\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40968\ : std_logic;
signal \N__40965\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40953\ : std_logic;
signal \N__40952\ : std_logic;
signal \N__40947\ : std_logic;
signal \N__40944\ : std_logic;
signal \N__40941\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40932\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40923\ : std_logic;
signal \N__40920\ : std_logic;
signal \N__40917\ : std_logic;
signal \N__40914\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40908\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40896\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40890\ : std_logic;
signal \N__40889\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40887\ : std_logic;
signal \N__40880\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40874\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40858\ : std_logic;
signal \N__40855\ : std_logic;
signal \N__40852\ : std_logic;
signal \N__40849\ : std_logic;
signal \N__40842\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40833\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40820\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40813\ : std_logic;
signal \N__40812\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40797\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40773\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40767\ : std_logic;
signal \N__40764\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40757\ : std_logic;
signal \N__40756\ : std_logic;
signal \N__40755\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40743\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40737\ : std_logic;
signal \N__40734\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40719\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40713\ : std_logic;
signal \N__40710\ : std_logic;
signal \N__40707\ : std_logic;
signal \N__40704\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40688\ : std_logic;
signal \N__40685\ : std_logic;
signal \N__40680\ : std_logic;
signal \N__40677\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40668\ : std_logic;
signal \N__40665\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40661\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40657\ : std_logic;
signal \N__40656\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40652\ : std_logic;
signal \N__40649\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40642\ : std_logic;
signal \N__40639\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40593\ : std_logic;
signal \N__40590\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40584\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40580\ : std_logic;
signal \N__40577\ : std_logic;
signal \N__40572\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40566\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40560\ : std_logic;
signal \N__40557\ : std_logic;
signal \N__40554\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40548\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40544\ : std_logic;
signal \N__40541\ : std_logic;
signal \N__40538\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40529\ : std_logic;
signal \N__40526\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40517\ : std_logic;
signal \N__40514\ : std_logic;
signal \N__40511\ : std_logic;
signal \N__40508\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40499\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40491\ : std_logic;
signal \N__40488\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40478\ : std_logic;
signal \N__40475\ : std_logic;
signal \N__40472\ : std_logic;
signal \N__40469\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40460\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40449\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40444\ : std_logic;
signal \N__40443\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40441\ : std_logic;
signal \N__40438\ : std_logic;
signal \N__40435\ : std_logic;
signal \N__40432\ : std_logic;
signal \N__40429\ : std_logic;
signal \N__40426\ : std_logic;
signal \N__40423\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40417\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40398\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40383\ : std_logic;
signal \N__40380\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40376\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40370\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40361\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40354\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40351\ : std_logic;
signal \N__40348\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40346\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40338\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40331\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40311\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40290\ : std_logic;
signal \N__40287\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40277\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40273\ : std_logic;
signal \N__40270\ : std_logic;
signal \N__40267\ : std_logic;
signal \N__40264\ : std_logic;
signal \N__40261\ : std_logic;
signal \N__40254\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40245\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40236\ : std_logic;
signal \N__40233\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40228\ : std_logic;
signal \N__40225\ : std_logic;
signal \N__40222\ : std_logic;
signal \N__40217\ : std_logic;
signal \N__40214\ : std_logic;
signal \N__40211\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40191\ : std_logic;
signal \N__40190\ : std_logic;
signal \N__40189\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40183\ : std_logic;
signal \N__40180\ : std_logic;
signal \N__40177\ : std_logic;
signal \N__40172\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40158\ : std_logic;
signal \N__40155\ : std_logic;
signal \N__40152\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40106\ : std_logic;
signal \N__40103\ : std_logic;
signal \N__40100\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40091\ : std_logic;
signal \N__40090\ : std_logic;
signal \N__40085\ : std_logic;
signal \N__40082\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40074\ : std_logic;
signal \N__40071\ : std_logic;
signal \N__40068\ : std_logic;
signal \N__40065\ : std_logic;
signal \N__40062\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40058\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40054\ : std_logic;
signal \N__40051\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40042\ : std_logic;
signal \N__40035\ : std_logic;
signal \N__40032\ : std_logic;
signal \N__40029\ : std_logic;
signal \N__40026\ : std_logic;
signal \N__40023\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40019\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40004\ : std_logic;
signal \N__39999\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39983\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39979\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39970\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39950\ : std_logic;
signal \N__39949\ : std_logic;
signal \N__39946\ : std_logic;
signal \N__39941\ : std_logic;
signal \N__39938\ : std_logic;
signal \N__39933\ : std_logic;
signal \N__39930\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39911\ : std_logic;
signal \N__39910\ : std_logic;
signal \N__39907\ : std_logic;
signal \N__39904\ : std_logic;
signal \N__39901\ : std_logic;
signal \N__39896\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39885\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39858\ : std_logic;
signal \N__39857\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39850\ : std_logic;
signal \N__39847\ : std_logic;
signal \N__39846\ : std_logic;
signal \N__39843\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39829\ : std_logic;
signal \N__39828\ : std_logic;
signal \N__39825\ : std_logic;
signal \N__39820\ : std_logic;
signal \N__39817\ : std_logic;
signal \N__39814\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39798\ : std_logic;
signal \N__39795\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39790\ : std_logic;
signal \N__39787\ : std_logic;
signal \N__39784\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39778\ : std_logic;
signal \N__39777\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39749\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39741\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39729\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39718\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39705\ : std_logic;
signal \N__39702\ : std_logic;
signal \N__39699\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39693\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39686\ : std_logic;
signal \N__39685\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39676\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39663\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39653\ : std_logic;
signal \N__39650\ : std_logic;
signal \N__39647\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39639\ : std_logic;
signal \N__39638\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39622\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39616\ : std_logic;
signal \N__39613\ : std_logic;
signal \N__39606\ : std_logic;
signal \N__39603\ : std_logic;
signal \N__39600\ : std_logic;
signal \N__39597\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39587\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39583\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39570\ : std_logic;
signal \N__39567\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39544\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39533\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39519\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39503\ : std_logic;
signal \N__39500\ : std_logic;
signal \N__39499\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39491\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39460\ : std_logic;
signal \N__39457\ : std_logic;
signal \N__39448\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39412\ : std_logic;
signal \N__39409\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39373\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39367\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39347\ : std_logic;
signal \N__39344\ : std_logic;
signal \N__39341\ : std_logic;
signal \N__39338\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39320\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39268\ : std_logic;
signal \N__39265\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39259\ : std_logic;
signal \N__39256\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39221\ : std_logic;
signal \N__39218\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39212\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39194\ : std_logic;
signal \N__39191\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39185\ : std_logic;
signal \N__39182\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39170\ : std_logic;
signal \N__39167\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39149\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39125\ : std_logic;
signal \N__39122\ : std_logic;
signal \N__39119\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39093\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39075\ : std_logic;
signal \N__39072\ : std_logic;
signal \N__39069\ : std_logic;
signal \N__39066\ : std_logic;
signal \N__39063\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39054\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39050\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39042\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39015\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39011\ : std_logic;
signal \N__39008\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39000\ : std_logic;
signal \N__38997\ : std_logic;
signal \N__38994\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38990\ : std_logic;
signal \N__38989\ : std_logic;
signal \N__38986\ : std_logic;
signal \N__38983\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38964\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38949\ : std_logic;
signal \N__38946\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38907\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38889\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38885\ : std_logic;
signal \N__38882\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38864\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38841\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38837\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38831\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38819\ : std_logic;
signal \N__38816\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38807\ : std_logic;
signal \N__38804\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38792\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38781\ : std_logic;
signal \N__38778\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38741\ : std_logic;
signal \N__38738\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38718\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38705\ : std_logic;
signal \N__38702\ : std_logic;
signal \N__38699\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38669\ : std_logic;
signal \N__38666\ : std_logic;
signal \N__38663\ : std_logic;
signal \N__38660\ : std_logic;
signal \N__38655\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38648\ : std_logic;
signal \N__38645\ : std_logic;
signal \N__38642\ : std_logic;
signal \N__38639\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38612\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38549\ : std_logic;
signal \N__38546\ : std_logic;
signal \N__38541\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38537\ : std_logic;
signal \N__38534\ : std_logic;
signal \N__38531\ : std_logic;
signal \N__38526\ : std_logic;
signal \N__38523\ : std_logic;
signal \N__38522\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38516\ : std_logic;
signal \N__38513\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38483\ : std_logic;
signal \N__38478\ : std_logic;
signal \N__38475\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38450\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38439\ : std_logic;
signal \N__38434\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38424\ : std_logic;
signal \N__38421\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38400\ : std_logic;
signal \N__38397\ : std_logic;
signal \N__38396\ : std_logic;
signal \N__38393\ : std_logic;
signal \N__38390\ : std_logic;
signal \N__38387\ : std_logic;
signal \N__38382\ : std_logic;
signal \N__38379\ : std_logic;
signal \N__38378\ : std_logic;
signal \N__38375\ : std_logic;
signal \N__38372\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38363\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38357\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38349\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38334\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38304\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38284\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38252\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38232\ : std_logic;
signal \N__38229\ : std_logic;
signal \N__38226\ : std_logic;
signal \N__38223\ : std_logic;
signal \N__38220\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38210\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38199\ : std_logic;
signal \N__38196\ : std_logic;
signal \N__38193\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38187\ : std_logic;
signal \N__38184\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38172\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38168\ : std_logic;
signal \N__38165\ : std_logic;
signal \N__38162\ : std_logic;
signal \N__38159\ : std_logic;
signal \N__38156\ : std_logic;
signal \N__38153\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38145\ : std_logic;
signal \N__38142\ : std_logic;
signal \N__38139\ : std_logic;
signal \N__38136\ : std_logic;
signal \N__38133\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38121\ : std_logic;
signal \N__38120\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38111\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38102\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38066\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38016\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38003\ : std_logic;
signal \N__38000\ : std_logic;
signal \N__37997\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37973\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37928\ : std_logic;
signal \N__37925\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37902\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37893\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37872\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37863\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37854\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37846\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37755\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37744\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37646\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37638\ : std_logic;
signal \N__37635\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37592\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37569\ : std_logic;
signal \N__37566\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37458\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37420\ : std_logic;
signal \N__37417\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37402\ : std_logic;
signal \N__37399\ : std_logic;
signal \N__37396\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37390\ : std_logic;
signal \N__37387\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37378\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37338\ : std_logic;
signal \N__37335\ : std_logic;
signal \N__37332\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37305\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37271\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37248\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37239\ : std_logic;
signal \N__37236\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37230\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37155\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37131\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37098\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37057\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37051\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37041\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37011\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36976\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36876\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36839\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36806\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36771\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36676\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36600\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36592\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36583\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36528\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36499\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36471\ : std_logic;
signal \N__36468\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36457\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36427\ : std_logic;
signal \N__36424\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36411\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36400\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36387\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36289\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36276\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36264\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36240\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36210\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36192\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36144\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36094\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36048\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35958\ : std_logic;
signal \N__35955\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35918\ : std_logic;
signal \N__35915\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35835\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35790\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35773\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35670\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35650\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35644\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35580\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35535\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35475\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35394\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35373\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35343\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35249\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35126\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35007\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34912\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34815\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34788\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34735\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34248\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34233\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34225\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34051\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34039\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33256\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33200\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32710\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32682\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32527\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32511\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32449\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31874\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31822\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31561\ : std_logic;
signal \N__31558\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31354\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31138\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30977\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30941\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30252\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29161\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29076\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28359\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27963\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27039\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25342\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24817\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18354\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \NEOPXL_c\ : std_logic;
signal \nx.n13325_cascade_\ : std_logic;
signal \nx.n11535_cascade_\ : std_logic;
signal \nx.n11672_cascade_\ : std_logic;
signal \nx.n13326\ : std_logic;
signal \nx.n11692\ : std_logic;
signal \nx.n12204\ : std_logic;
signal \nx.n11696_cascade_\ : std_logic;
signal \nx.n7131_cascade_\ : std_logic;
signal \nx.n13263_cascade_\ : std_logic;
signal \nx.n7120_cascade_\ : std_logic;
signal \nx.n13262_cascade_\ : std_logic;
signal \nx.n3739\ : std_logic;
signal \nx.n3739_cascade_\ : std_logic;
signal \nx.n7120\ : std_logic;
signal \nx.n9700_cascade_\ : std_logic;
signal \nx.n7131\ : std_logic;
signal \nx.n12117_cascade_\ : std_logic;
signal \n7239_cascade_\ : std_logic;
signal \nx.n9700\ : std_logic;
signal \nx.n9702\ : std_logic;
signal \nx.n11606\ : std_logic;
signal update_color : std_logic;
signal \nx.n10_adj_653\ : std_logic;
signal \nx.n13271\ : std_logic;
signal \nx.n12369_cascade_\ : std_logic;
signal neo_pixel_transmitter_t0_15 : std_logic;
signal neo_pixel_transmitter_t0_8 : std_logic;
signal \nx.n2908_cascade_\ : std_logic;
signal \nx.n3007_cascade_\ : std_logic;
signal \nx.n3106_cascade_\ : std_logic;
signal \nx.n19_adj_698\ : std_logic;
signal \nx.n3105_cascade_\ : std_logic;
signal \nx.n3100_cascade_\ : std_logic;
signal \nx.n29_adj_697_cascade_\ : std_logic;
signal \nx.n12331_cascade_\ : std_logic;
signal \nx.n12335\ : std_logic;
signal \nx.n37_adj_695_cascade_\ : std_logic;
signal \nx.n12333\ : std_logic;
signal \nx.n31_adj_691_cascade_\ : std_logic;
signal \nx.n49_adj_693_cascade_\ : std_logic;
signal \nx.n48_adj_692\ : std_logic;
signal \nx.n3116_cascade_\ : std_logic;
signal \bfn_1_26_0_\ : std_logic;
signal \nx.n3176\ : std_logic;
signal \nx.n10888\ : std_logic;
signal \nx.n10889\ : std_logic;
signal \nx.n10890\ : std_logic;
signal \nx.n3106\ : std_logic;
signal \nx.n3173\ : std_logic;
signal \nx.n10891\ : std_logic;
signal \nx.n3105\ : std_logic;
signal \nx.n3172\ : std_logic;
signal \nx.n10892\ : std_logic;
signal \nx.n10893\ : std_logic;
signal \nx.n3170\ : std_logic;
signal \nx.n10894\ : std_logic;
signal \nx.n10895\ : std_logic;
signal \nx.n3102\ : std_logic;
signal \nx.n3169\ : std_logic;
signal \bfn_1_27_0_\ : std_logic;
signal \nx.n10896\ : std_logic;
signal \nx.n3100\ : std_logic;
signal \nx.n3167\ : std_logic;
signal \nx.n10897\ : std_logic;
signal \nx.n10898\ : std_logic;
signal \nx.n10899\ : std_logic;
signal \nx.n10900\ : std_logic;
signal \nx.n3163\ : std_logic;
signal \nx.n10901\ : std_logic;
signal \nx.n10902\ : std_logic;
signal \nx.n10903\ : std_logic;
signal \bfn_1_28_0_\ : std_logic;
signal \nx.n10904\ : std_logic;
signal \nx.n10905\ : std_logic;
signal \nx.n10906\ : std_logic;
signal \nx.n10907\ : std_logic;
signal \nx.n10908\ : std_logic;
signal \nx.n10909\ : std_logic;
signal \nx.n3154\ : std_logic;
signal \nx.n10910\ : std_logic;
signal \nx.n10911\ : std_logic;
signal \nx.n3153\ : std_logic;
signal \bfn_1_29_0_\ : std_logic;
signal \nx.n3152\ : std_logic;
signal \nx.n10912\ : std_logic;
signal \nx.n10913\ : std_logic;
signal \nx.n10914\ : std_logic;
signal \nx.n10_adj_619_cascade_\ : std_logic;
signal \nx.n12_adj_621_cascade_\ : std_logic;
signal \nx.n1136_cascade_\ : std_logic;
signal \nx.n1203_cascade_\ : std_logic;
signal \nx.n1208_cascade_\ : std_logic;
signal \bfn_1_31_0_\ : std_logic;
signal \nx.n10453\ : std_logic;
signal \nx.n10454\ : std_logic;
signal \nx.n10455\ : std_logic;
signal \nx.n10456\ : std_logic;
signal \nx.n10457\ : std_logic;
signal \nx.n10458\ : std_logic;
signal \nx.n10459\ : std_logic;
signal \nx.n10460\ : std_logic;
signal \bfn_1_32_0_\ : std_logic;
signal \nx.n1203\ : std_logic;
signal \nx.n1270\ : std_logic;
signal \nx.n1302_cascade_\ : std_logic;
signal \nx.n1276\ : std_logic;
signal \nx.n1209\ : std_logic;
signal \nx.n1206_cascade_\ : std_logic;
signal \nx.n1273\ : std_logic;
signal \nx.n7\ : std_logic;
signal neo_pixel_transmitter_t0_23 : std_logic;
signal neo_pixel_transmitter_t0_24 : std_logic;
signal \nx.n7_adj_713_cascade_\ : std_logic;
signal \nx.n13491\ : std_logic;
signal \nx.n12933_cascade_\ : std_logic;
signal \nx.n12939\ : std_logic;
signal \nx.n10918\ : std_logic;
signal \nx.start\ : std_logic;
signal \nx.n18_adj_711_cascade_\ : std_logic;
signal \nx.n20_adj_712\ : std_logic;
signal neo_pixel_transmitter_t0_6 : std_logic;
signal neo_pixel_transmitter_t0_14 : std_logic;
signal neo_pixel_transmitter_t0_5 : std_logic;
signal neopxl_color_prev_5 : std_logic;
signal n10_adj_776 : std_logic;
signal neo_pixel_transmitter_t0_3 : std_logic;
signal n12_adj_774 : std_logic;
signal neo_pixel_transmitter_t0_12 : std_logic;
signal \nx.neo_pixel_transmitter_done\ : std_logic;
signal \nx.n11487_cascade_\ : std_logic;
signal \nx.n103\ : std_logic;
signal n9_adj_777 : std_logic;
signal neopxl_color_prev_4 : std_logic;
signal state_0_adj_727 : std_logic;
signal state_1_adj_726 : std_logic;
signal n7239 : std_logic;
signal \nx.n7392\ : std_logic;
signal \nx.n13155\ : std_logic;
signal \nx.n13456_cascade_\ : std_logic;
signal \nx.n13156\ : std_logic;
signal \nx.n13459\ : std_logic;
signal \nx.n4_adj_642\ : std_logic;
signal neo_pixel_transmitter_t0_26 : std_logic;
signal neo_pixel_transmitter_t0_16 : std_logic;
signal \nx.color_bit_N_571_4\ : std_logic;
signal \nx.n13158\ : std_logic;
signal \nx.n59\ : std_logic;
signal \nx.n12371\ : std_logic;
signal \nx.n13042\ : std_logic;
signal \nx.n10947\ : std_logic;
signal \nx.n10947_cascade_\ : std_logic;
signal \nx.n10975\ : std_logic;
signal \nx.n3008_cascade_\ : std_logic;
signal \nx.n3096\ : std_logic;
signal \nx.n3096_cascade_\ : std_logic;
signal \nx.n47_adj_694\ : std_logic;
signal \nx.n45\ : std_logic;
signal \nx.n49_cascade_\ : std_logic;
signal \nx.n3017_cascade_\ : std_logic;
signal \nx.n3086\ : std_logic;
signal \nx.n3087\ : std_logic;
signal \nx.n3086_cascade_\ : std_logic;
signal \nx.n3085\ : std_logic;
signal \nx.n42_adj_689\ : std_logic;
signal \nx.n3103\ : std_logic;
signal \nx.n3097\ : std_logic;
signal \nx.n3164\ : std_logic;
signal \nx.n3097_cascade_\ : std_logic;
signal \nx.n3168\ : std_logic;
signal \nx.n35_adj_699_cascade_\ : std_logic;
signal \nx.n3101\ : std_logic;
signal \nx.n12337\ : std_logic;
signal \nx.n3109\ : std_logic;
signal \nx.n12349\ : std_logic;
signal \nx.n3174\ : std_logic;
signal \nx.n23_adj_700\ : std_logic;
signal \nx.n3107\ : std_logic;
signal \nx.n3162\ : std_logic;
signal \nx.n12327_cascade_\ : std_logic;
signal \nx.n3095\ : std_logic;
signal \nx.n3166\ : std_logic;
signal \nx.n3177\ : std_logic;
signal \nx.n3209\ : std_logic;
signal \nx.n3171\ : std_logic;
signal \nx.n3175\ : std_logic;
signal \nx.n3108\ : std_logic;
signal \nx.n3165\ : std_logic;
signal \nx.n3098\ : std_logic;
signal \nx.n13_adj_696_cascade_\ : std_logic;
signal \nx.n31_adj_702\ : std_logic;
signal \nx.n21_adj_701\ : std_logic;
signal \nx.n12325_cascade_\ : std_logic;
signal \nx.n12339\ : std_logic;
signal \nx.n12347\ : std_logic;
signal \nx.n3151\ : std_logic;
signal \nx.n61\ : std_logic;
signal \nx.n3099\ : std_logic;
signal neopxl_color_prev_7 : std_logic;
signal \nx.n54\ : std_logic;
signal \nx.n43_adj_709_cascade_\ : std_logic;
signal \nx.n49_adj_710\ : std_logic;
signal \state_3_N_377_1\ : std_logic;
signal \nx.n3084\ : std_logic;
signal \nx.n1177\ : std_logic;
signal \bfn_2_29_0_\ : std_logic;
signal \nx.n1109\ : std_logic;
signal \nx.n1176\ : std_logic;
signal \nx.n10461\ : std_logic;
signal \nx.n10462\ : std_logic;
signal \nx.n1174\ : std_logic;
signal \nx.n10463\ : std_logic;
signal \nx.n10464\ : std_logic;
signal \nx.n10465\ : std_logic;
signal \nx.n1171\ : std_logic;
signal \nx.n10466\ : std_logic;
signal \nx.n10467\ : std_logic;
signal \nx.n1202\ : std_logic;
signal \nx.n1173\ : std_logic;
signal \nx.n1172\ : std_logic;
signal \nx.n1204\ : std_logic;
signal \nx.n1271\ : std_logic;
signal \nx.n1204_cascade_\ : std_logic;
signal \nx.n11_adj_624\ : std_logic;
signal \nx.n13\ : std_logic;
signal \nx.n1206\ : std_logic;
signal \nx.n1275\ : std_logic;
signal \nx.n1235_cascade_\ : std_logic;
signal \nx.n1208\ : std_logic;
signal \nx.n1175\ : std_logic;
signal \nx.n1136\ : std_logic;
signal \nx.n1207\ : std_logic;
signal \nx.n1274\ : std_logic;
signal \nx.n1207_cascade_\ : std_logic;
signal \nx.n1306_cascade_\ : std_logic;
signal \nx.n10_adj_626\ : std_logic;
signal \bfn_2_31_0_\ : std_logic;
signal \nx.n10573\ : std_logic;
signal \nx.n10574\ : std_logic;
signal \nx.n10575\ : std_logic;
signal \nx.n10576\ : std_logic;
signal \nx.n10577\ : std_logic;
signal \nx.n10578\ : std_logic;
signal \nx.n10579\ : std_logic;
signal \nx.n10580\ : std_logic;
signal \bfn_2_32_0_\ : std_logic;
signal \nx.n1301\ : std_logic;
signal \nx.n10581\ : std_logic;
signal \nx.n1302\ : std_logic;
signal \nx.n1369\ : std_logic;
signal neo_pixel_transmitter_t0_1 : std_logic;
signal neo_pixel_transmitter_t0_31 : std_logic;
signal neo_pixel_transmitter_t0_4 : std_logic;
signal \bfn_3_17_0_\ : std_logic;
signal \nx.n10479\ : std_logic;
signal \nx.n10480\ : std_logic;
signal \nx.n10481\ : std_logic;
signal \nx.n10482\ : std_logic;
signal \nx.n10483\ : std_logic;
signal \nx.n10484\ : std_logic;
signal \nx.n10485\ : std_logic;
signal \nx.n10486\ : std_logic;
signal \bfn_3_18_0_\ : std_logic;
signal \nx.n10487\ : std_logic;
signal \nx.n10488\ : std_logic;
signal \nx.n10489\ : std_logic;
signal \nx.n10490\ : std_logic;
signal \nx.n10491\ : std_logic;
signal \nx.n10492\ : std_logic;
signal \nx.n10493\ : std_logic;
signal \nx.n10494\ : std_logic;
signal \bfn_3_19_0_\ : std_logic;
signal \nx.n10495\ : std_logic;
signal \nx.n10496\ : std_logic;
signal \nx.n10497\ : std_logic;
signal \nx.n10498\ : std_logic;
signal \nx.n10499\ : std_logic;
signal \nx.n10500\ : std_logic;
signal \nx.n10501\ : std_logic;
signal \nx.n10502\ : std_logic;
signal \bfn_3_20_0_\ : std_logic;
signal \nx.n10503\ : std_logic;
signal \nx.n10504\ : std_logic;
signal \nx.n10505\ : std_logic;
signal \nx.n10506\ : std_logic;
signal \nx.n10507\ : std_logic;
signal \nx.n10508\ : std_logic;
signal \nx.n10509\ : std_logic;
signal \bfn_3_21_0_\ : std_logic;
signal \nx.n32_adj_651\ : std_logic;
signal timer_1 : std_logic;
signal \nx.n11533\ : std_logic;
signal \nx.n10422\ : std_logic;
signal \nx.one_wire_N_528_2\ : std_logic;
signal \nx.n10423\ : std_logic;
signal \nx.n30_adj_598\ : std_logic;
signal timer_3 : std_logic;
signal \nx.one_wire_N_528_3\ : std_logic;
signal \nx.n10424\ : std_logic;
signal \nx.n29\ : std_logic;
signal timer_4 : std_logic;
signal \nx.one_wire_N_528_4\ : std_logic;
signal \nx.n10425\ : std_logic;
signal timer_5 : std_logic;
signal \nx.n28\ : std_logic;
signal \nx.one_wire_N_528_5\ : std_logic;
signal \nx.n10426\ : std_logic;
signal timer_6 : std_logic;
signal \nx.n27\ : std_logic;
signal \nx.one_wire_N_528_6\ : std_logic;
signal \nx.n10427\ : std_logic;
signal \nx.one_wire_N_528_7\ : std_logic;
signal \nx.n10428\ : std_logic;
signal \nx.n10429\ : std_logic;
signal \nx.n25\ : std_logic;
signal timer_8 : std_logic;
signal \nx.one_wire_N_528_8\ : std_logic;
signal \bfn_3_22_0_\ : std_logic;
signal \nx.one_wire_N_528_9\ : std_logic;
signal \nx.n10430\ : std_logic;
signal timer_10 : std_logic;
signal \nx.one_wire_N_528_10\ : std_logic;
signal \nx.n10431\ : std_logic;
signal \nx.n10432\ : std_logic;
signal \nx.one_wire_N_528_11\ : std_logic;
signal timer_12 : std_logic;
signal \nx.n21_adj_620\ : std_logic;
signal \nx.n10433\ : std_logic;
signal \nx.n12945\ : std_logic;
signal \nx.n10434\ : std_logic;
signal \nx.n12947\ : std_logic;
signal \nx.n19_adj_622\ : std_logic;
signal timer_14 : std_logic;
signal \nx.n10435\ : std_logic;
signal \nx.n10436\ : std_logic;
signal \nx.n10436_THRU_CRY_0_THRU_CO\ : std_logic;
signal \nx.n12949\ : std_logic;
signal \nx.n18_adj_623\ : std_logic;
signal timer_15 : std_logic;
signal \bfn_3_23_0_\ : std_logic;
signal \nx.n12951\ : std_logic;
signal \nx.n17\ : std_logic;
signal timer_16 : std_logic;
signal \nx.n10437\ : std_logic;
signal \nx.n12953\ : std_logic;
signal \nx.n10438\ : std_logic;
signal \nx.n12955\ : std_logic;
signal \nx.n10439\ : std_logic;
signal \nx.n12957\ : std_logic;
signal \nx.n10440\ : std_logic;
signal \nx.n12959\ : std_logic;
signal \nx.n10441\ : std_logic;
signal \nx.n10442\ : std_logic;
signal \nx.n10442_THRU_CRY_0_THRU_CO\ : std_logic;
signal \nx.n10442_THRU_CRY_1_THRU_CO\ : std_logic;
signal \nx.n12961\ : std_logic;
signal \bfn_3_24_0_\ : std_logic;
signal \nx.n12963\ : std_logic;
signal \nx.n10443\ : std_logic;
signal \nx.n12965\ : std_logic;
signal \nx.n10\ : std_logic;
signal timer_23 : std_logic;
signal \nx.n10444\ : std_logic;
signal \nx.n12967\ : std_logic;
signal \nx.n9\ : std_logic;
signal timer_24 : std_logic;
signal \nx.n10445\ : std_logic;
signal \nx.n12969\ : std_logic;
signal \nx.n10446\ : std_logic;
signal \nx.n12971\ : std_logic;
signal \nx.n7_adj_597\ : std_logic;
signal timer_26 : std_logic;
signal \nx.n10447\ : std_logic;
signal \nx.n10448\ : std_logic;
signal \GNDG0\ : std_logic;
signal \nx.n10448_THRU_CRY_0_THRU_CO\ : std_logic;
signal \nx.n10448_THRU_CRY_1_THRU_CO\ : std_logic;
signal \nx.n12973\ : std_logic;
signal \bfn_3_25_0_\ : std_logic;
signal \nx.n12975\ : std_logic;
signal \nx.n10449\ : std_logic;
signal \nx.n12977\ : std_logic;
signal \nx.n10450\ : std_logic;
signal \nx.n12979\ : std_logic;
signal \nx.n10451\ : std_logic;
signal timer_31 : std_logic;
signal \nx.n2\ : std_logic;
signal \nx.n12981\ : std_logic;
signal \nx.n10452\ : std_logic;
signal \nx.n7181\ : std_logic;
signal timer_27 : std_logic;
signal neo_pixel_transmitter_t0_27 : std_logic;
signal \nx.n6\ : std_logic;
signal \nx.n3077\ : std_logic;
signal \bfn_3_26_0_\ : std_logic;
signal \nx.n3076\ : std_logic;
signal \nx.n10862\ : std_logic;
signal \nx.n3008\ : std_logic;
signal \nx.n3075\ : std_logic;
signal \nx.n10863\ : std_logic;
signal \nx.n3007\ : std_logic;
signal \nx.n3074\ : std_logic;
signal \nx.n10864\ : std_logic;
signal \nx.n3073\ : std_logic;
signal \nx.n10865\ : std_logic;
signal \nx.n3072\ : std_logic;
signal \nx.n10866\ : std_logic;
signal \nx.n3071\ : std_logic;
signal \nx.n10867\ : std_logic;
signal \nx.n3070\ : std_logic;
signal \nx.n10868\ : std_logic;
signal \nx.n10869\ : std_logic;
signal \nx.n3069\ : std_logic;
signal \bfn_3_27_0_\ : std_logic;
signal \nx.n3001\ : std_logic;
signal \nx.n3068\ : std_logic;
signal \nx.n10870\ : std_logic;
signal \nx.n3067\ : std_logic;
signal \nx.n10871\ : std_logic;
signal \nx.n2999\ : std_logic;
signal \nx.n3066\ : std_logic;
signal \nx.n10872\ : std_logic;
signal \nx.n3065\ : std_logic;
signal \nx.n10873\ : std_logic;
signal \nx.n3064\ : std_logic;
signal \nx.n10874\ : std_logic;
signal \nx.n3063\ : std_logic;
signal \nx.n10875\ : std_logic;
signal \nx.n10876\ : std_logic;
signal \nx.n10877\ : std_logic;
signal \bfn_3_28_0_\ : std_logic;
signal \nx.n10878\ : std_logic;
signal \nx.n3059\ : std_logic;
signal \nx.n10879\ : std_logic;
signal \nx.n10880\ : std_logic;
signal \nx.n10881\ : std_logic;
signal \nx.n10882\ : std_logic;
signal \nx.n3055\ : std_logic;
signal \nx.n10883\ : std_logic;
signal \nx.n3054\ : std_logic;
signal \nx.n10884\ : std_logic;
signal \nx.n10885\ : std_logic;
signal \nx.n3053\ : std_logic;
signal \bfn_3_29_0_\ : std_logic;
signal \nx.n3052\ : std_logic;
signal \nx.n10886\ : std_logic;
signal \nx.n10887\ : std_logic;
signal \nx.n3083\ : std_logic;
signal \nx.n45_adj_707\ : std_logic;
signal \nx.n11_adj_628_cascade_\ : std_logic;
signal \nx.n16_adj_627\ : std_logic;
signal \nx.n1307\ : std_logic;
signal \nx.n1334_cascade_\ : std_logic;
signal \nx.n1374\ : std_logic;
signal \nx.n1277\ : std_logic;
signal \nx.n1309\ : std_logic;
signal \nx.n1376\ : std_logic;
signal \nx.n1309_cascade_\ : std_logic;
signal \nx.n1272\ : std_logic;
signal \nx.n1205\ : std_logic;
signal \nx.n1235\ : std_logic;
signal \nx.n1377\ : std_logic;
signal \bfn_3_31_0_\ : std_logic;
signal \nx.n10582\ : std_logic;
signal \nx.n10583\ : std_logic;
signal \nx.n10584\ : std_logic;
signal \nx.n10585\ : std_logic;
signal \nx.n10586\ : std_logic;
signal \nx.n10587\ : std_logic;
signal \nx.n10588\ : std_logic;
signal \nx.n10589\ : std_logic;
signal \bfn_3_32_0_\ : std_logic;
signal \nx.n10590\ : std_logic;
signal \nx.n10591\ : std_logic;
signal \nx.n1303\ : std_logic;
signal \nx.n1370\ : std_logic;
signal \nx.n1400\ : std_logic;
signal \nx.n3\ : std_logic;
signal timer_30 : std_logic;
signal neo_pixel_transmitter_t0_30 : std_logic;
signal \nx.n31_adj_650\ : std_logic;
signal \nx.n16_adj_661\ : std_logic;
signal timer_17 : std_logic;
signal neo_pixel_transmitter_t0_17 : std_logic;
signal timer_2 : std_logic;
signal neo_pixel_transmitter_t0_2 : std_logic;
signal timer_29 : std_logic;
signal timer_9 : std_logic;
signal neo_pixel_transmitter_t0_10 : std_logic;
signal \nx.n23_adj_617\ : std_logic;
signal neo_pixel_transmitter_t0_29 : std_logic;
signal \nx.n4\ : std_logic;
signal timer_11 : std_logic;
signal timer_21 : std_logic;
signal timer_13 : std_logic;
signal neo_pixel_transmitter_t0_11 : std_logic;
signal \nx.n22_adj_618\ : std_logic;
signal neo_pixel_transmitter_t0_13 : std_logic;
signal \nx.n20\ : std_logic;
signal timer_7 : std_logic;
signal \nx.n13159\ : std_logic;
signal neo_pixel_transmitter_t0_21 : std_logic;
signal \nx.n12\ : std_logic;
signal timer_25 : std_logic;
signal timer_18 : std_logic;
signal \nx.n5\ : std_logic;
signal neo_pixel_transmitter_t0_25 : std_logic;
signal \nx.n8\ : std_logic;
signal neo_pixel_transmitter_t0_18 : std_logic;
signal \nx.n15\ : std_logic;
signal timer_28 : std_logic;
signal neo_pixel_transmitter_t0_28 : std_logic;
signal \nx.n2995_cascade_\ : std_logic;
signal \nx.n44_adj_681\ : std_logic;
signal \nx.n33_adj_682_cascade_\ : std_logic;
signal \nx.n48\ : std_logic;
signal \nx.n3005\ : std_logic;
signal neo_pixel_transmitter_t0_7 : std_logic;
signal \nx.n26\ : std_logic;
signal \nx.n3006\ : std_logic;
signal \nx.n2899_cascade_\ : std_logic;
signal \nx.n2998\ : std_logic;
signal \nx.n2894_cascade_\ : std_logic;
signal \nx.n2985\ : std_logic;
signal \nx.n2985_cascade_\ : std_logic;
signal \nx.n2986\ : std_logic;
signal \nx.n40_adj_683\ : std_logic;
signal \nx.n43_adj_677\ : std_logic;
signal \nx.n40_adj_678\ : std_logic;
signal \nx.n47_cascade_\ : std_logic;
signal \nx.n2918_cascade_\ : std_logic;
signal \nx.n3000\ : std_logic;
signal \nx.n38_adj_676\ : std_logic;
signal \nx.n2996\ : std_logic;
signal \nx.n2997\ : std_logic;
signal \nx.n2987\ : std_logic;
signal \nx.n3004\ : std_logic;
signal \nx.n2988\ : std_logic;
signal \nx.n2988_cascade_\ : std_logic;
signal \nx.n41_adj_686\ : std_logic;
signal \nx.n2994_cascade_\ : std_logic;
signal \nx.n3002\ : std_logic;
signal \nx.n42_adj_684\ : std_logic;
signal \nx.n3009\ : std_logic;
signal \nx.n2992\ : std_logic;
signal \nx.n2989\ : std_logic;
signal \nx.n3056\ : std_logic;
signal \nx.n3104\ : std_logic;
signal \nx.n3088_cascade_\ : std_logic;
signal \nx.n44_adj_690\ : std_logic;
signal \nx.n3061\ : std_logic;
signal \nx.n2994\ : std_logic;
signal \nx.n2991\ : std_logic;
signal \nx.n3058\ : std_logic;
signal \nx.n3161\ : std_logic;
signal \nx.n12353\ : std_logic;
signal \nx.n3160\ : std_logic;
signal \nx.n12355\ : std_logic;
signal \nx.n12357_cascade_\ : std_logic;
signal \nx.n3159\ : std_logic;
signal \nx.n3158\ : std_logic;
signal \nx.n12359_cascade_\ : std_logic;
signal \nx.n3157\ : std_logic;
signal \nx.n12361_cascade_\ : std_logic;
signal \nx.n3090\ : std_logic;
signal \nx.n3156\ : std_logic;
signal \nx.n12363_cascade_\ : std_logic;
signal \nx.n3116\ : std_logic;
signal \nx.n3088\ : std_logic;
signal \nx.n12365_cascade_\ : std_logic;
signal \nx.n3155\ : std_logic;
signal \nx.n12367\ : std_logic;
signal \nx.n2990\ : std_logic;
signal \nx.n3057\ : std_logic;
signal \nx.n3089\ : std_logic;
signal \nx.bit_ctr_0\ : std_logic;
signal \bfn_4_27_0_\ : std_logic;
signal \nx.bit_ctr_1\ : std_logic;
signal \nx.n10391\ : std_logic;
signal \nx.bit_ctr_2\ : std_logic;
signal \nx.n10392\ : std_logic;
signal \nx.bit_ctr_3\ : std_logic;
signal \nx.n10393\ : std_logic;
signal \nx.bit_ctr_4\ : std_logic;
signal \nx.n10394\ : std_logic;
signal \nx.n10395\ : std_logic;
signal \nx.n10396\ : std_logic;
signal \nx.n10397\ : std_logic;
signal \nx.n10398\ : std_logic;
signal \bfn_4_28_0_\ : std_logic;
signal \nx.n10399\ : std_logic;
signal \nx.n10400\ : std_logic;
signal \nx.n10401\ : std_logic;
signal \nx.n10402\ : std_logic;
signal \nx.n10403\ : std_logic;
signal \nx.n10404\ : std_logic;
signal \nx.n10405\ : std_logic;
signal \nx.n10406\ : std_logic;
signal \bfn_4_29_0_\ : std_logic;
signal \nx.n10407\ : std_logic;
signal \nx.n10408\ : std_logic;
signal \nx.n10409\ : std_logic;
signal \nx.n10410\ : std_logic;
signal \nx.n10411\ : std_logic;
signal \nx.n10412\ : std_logic;
signal \nx.n10413\ : std_logic;
signal \nx.n10414\ : std_logic;
signal \nx.bit_ctr_24\ : std_logic;
signal \bfn_4_30_0_\ : std_logic;
signal \nx.n10415\ : std_logic;
signal \nx.n10416\ : std_logic;
signal \nx.n10417\ : std_logic;
signal \nx.n10418\ : std_logic;
signal \nx.n10419\ : std_logic;
signal \nx.n10420\ : std_logic;
signal \nx.n10421\ : std_logic;
signal \nx.n7230\ : std_logic;
signal \nx.n7411\ : std_logic;
signal \nx.n1308\ : std_logic;
signal \nx.n1375\ : std_logic;
signal \nx.n1373\ : std_logic;
signal \nx.n1306\ : std_logic;
signal \nx.n1371\ : std_logic;
signal \nx.n1304\ : std_logic;
signal \nx.n1305\ : std_logic;
signal \nx.n1372\ : std_logic;
signal \nx.n1334\ : std_logic;
signal \nx.n1404_cascade_\ : std_logic;
signal \nx.bit_ctr_23\ : std_logic;
signal \nx.n47_adj_706\ : std_logic;
signal \nx.n1404\ : std_logic;
signal \nx.n1471\ : std_logic;
signal \nx.bit_ctr_21\ : std_logic;
signal \nx.n1477\ : std_logic;
signal \nx.n1509_cascade_\ : std_logic;
signal \nx.n16_adj_629\ : std_logic;
signal \nx.n18_adj_630_cascade_\ : std_logic;
signal \nx.n13_adj_631\ : std_logic;
signal \nx.n1469\ : std_logic;
signal \nx.n1433_cascade_\ : std_logic;
signal \nx.n1402\ : std_logic;
signal \nx.n1501_cascade_\ : std_logic;
signal \nx.n9672\ : std_logic;
signal timer_22 : std_logic;
signal timer_19 : std_logic;
signal n13171 : std_logic;
signal n13170 : std_logic;
signal neo_pixel_transmitter_t0_9 : std_logic;
signal \nx.n24\ : std_logic;
signal neo_pixel_transmitter_t0_19 : std_logic;
signal \nx.n14\ : std_logic;
signal neopxl_color_prev_6 : std_logic;
signal neopxl_color_prev_15 : std_logic;
signal n11_adj_775 : std_logic;
signal neopxl_color_prev_13 : std_logic;
signal \nx.n13_adj_649\ : std_logic;
signal timer_20 : std_logic;
signal neo_pixel_transmitter_t0_20 : std_logic;
signal \nx.n2809_cascade_\ : std_logic;
signal \nx.n31_adj_613_cascade_\ : std_logic;
signal \nx.n39_adj_614\ : std_logic;
signal \nx.n2896_cascade_\ : std_logic;
signal \nx.n2898_cascade_\ : std_logic;
signal \nx.n42_adj_675_cascade_\ : std_logic;
signal \nx.n32_adj_674\ : std_logic;
signal \nx.n46\ : std_logic;
signal \nx.n2977\ : std_logic;
signal \bfn_5_22_0_\ : std_logic;
signal \nx.n2976\ : std_logic;
signal \nx.n10837\ : std_logic;
signal \nx.n2908\ : std_logic;
signal \nx.n2975\ : std_logic;
signal \nx.n10838\ : std_logic;
signal \nx.n2907\ : std_logic;
signal \nx.n2974\ : std_logic;
signal \nx.n10839\ : std_logic;
signal \nx.n2906\ : std_logic;
signal \nx.n2973\ : std_logic;
signal \nx.n10840\ : std_logic;
signal \nx.n2972\ : std_logic;
signal \nx.n10841\ : std_logic;
signal \nx.n10842\ : std_logic;
signal \nx.n2970\ : std_logic;
signal \nx.n10843\ : std_logic;
signal \nx.n10844\ : std_logic;
signal \nx.n2969\ : std_logic;
signal \bfn_5_23_0_\ : std_logic;
signal \nx.n2901\ : std_logic;
signal \nx.n2968\ : std_logic;
signal \nx.n10845\ : std_logic;
signal \nx.n2967\ : std_logic;
signal \nx.n10846\ : std_logic;
signal \nx.n2899\ : std_logic;
signal \nx.n2966\ : std_logic;
signal \nx.n10847\ : std_logic;
signal \nx.n2898\ : std_logic;
signal \nx.n2965\ : std_logic;
signal \nx.n10848\ : std_logic;
signal \nx.n2897\ : std_logic;
signal \nx.n2964\ : std_logic;
signal \nx.n10849\ : std_logic;
signal \nx.n2896\ : std_logic;
signal \nx.n2963\ : std_logic;
signal \nx.n10850\ : std_logic;
signal \nx.n2962\ : std_logic;
signal \nx.n10851\ : std_logic;
signal \nx.n10852\ : std_logic;
signal \bfn_5_24_0_\ : std_logic;
signal \nx.n2960\ : std_logic;
signal \nx.n10853\ : std_logic;
signal \nx.n2959\ : std_logic;
signal \nx.n10854\ : std_logic;
signal \nx.n2958\ : std_logic;
signal \nx.n10855\ : std_logic;
signal \nx.n2957\ : std_logic;
signal \nx.n10856\ : std_logic;
signal \nx.n2956\ : std_logic;
signal \nx.n10857\ : std_logic;
signal \nx.n2955\ : std_logic;
signal \nx.n10858\ : std_logic;
signal \nx.n2954\ : std_logic;
signal \nx.n10859\ : std_logic;
signal \nx.n10860\ : std_logic;
signal \nx.n2953\ : std_logic;
signal \bfn_5_25_0_\ : std_logic;
signal \nx.n10861\ : std_logic;
signal \nx.n2984\ : std_logic;
signal \nx.n2961\ : std_logic;
signal \nx.n2894\ : std_logic;
signal \nx.n2993\ : std_logic;
signal \nx.n3060\ : std_logic;
signal \nx.n2993_cascade_\ : std_logic;
signal \nx.n3092\ : std_logic;
signal \nx.n3091\ : std_logic;
signal \nx.n3092_cascade_\ : std_logic;
signal \nx.n46_adj_688\ : std_logic;
signal \nx.n50\ : std_logic;
signal \nx.n3093\ : std_logic;
signal \nx.n36_adj_687\ : std_logic;
signal \nx.n1077\ : std_logic;
signal \bfn_5_26_0_\ : std_logic;
signal \nx.n10468\ : std_logic;
signal \nx.n10469\ : std_logic;
signal \nx.n10470\ : std_logic;
signal \nx.n10471\ : std_logic;
signal \nx.n10472\ : std_logic;
signal \nx.n10473\ : std_logic;
signal \nx.n1103\ : std_logic;
signal \nx.n46_adj_705\ : std_logic;
signal \nx.n1075\ : std_logic;
signal \nx.n1107\ : std_logic;
signal \nx.n1073\ : std_logic;
signal \nx.n1105\ : std_logic;
signal \nx.n11617_cascade_\ : std_logic;
signal \nx.n1076\ : std_logic;
signal \nx.n1037_cascade_\ : std_logic;
signal \nx.n1108\ : std_logic;
signal \nx.n1007\ : std_logic;
signal \nx.n1074\ : std_logic;
signal \nx.n1106\ : std_logic;
signal \nx.n1009\ : std_logic;
signal \nx.bit_ctr_25\ : std_logic;
signal \nx.n1009_cascade_\ : std_logic;
signal \nx.n7_adj_616\ : std_logic;
signal \nx.bit_ctr_5\ : std_logic;
signal \nx.bit_ctr_6\ : std_logic;
signal \nx.n44_adj_708\ : std_logic;
signal \nx.n1005\ : std_logic;
signal \nx.n1072\ : std_logic;
signal \nx.n1005_cascade_\ : std_logic;
signal \nx.n1037\ : std_logic;
signal \nx.n1104\ : std_logic;
signal \nx.n1008\ : std_logic;
signal \nx.n7084_cascade_\ : std_logic;
signal \nx.n838_cascade_\ : std_logic;
signal \nx.n12595_cascade_\ : std_logic;
signal \nx.n9618_cascade_\ : std_logic;
signal \nx.n608\ : std_logic;
signal \nx.n11738_cascade_\ : std_logic;
signal \nx.n708\ : std_logic;
signal \nx.n739_cascade_\ : std_logic;
signal \nx.n11738\ : std_logic;
signal \nx.n807\ : std_logic;
signal \nx.bit_ctr_31\ : std_logic;
signal \nx.n9618\ : std_logic;
signal \nx.bit_ctr_29\ : std_logic;
signal \nx.n11771_cascade_\ : std_logic;
signal \nx.n1470\ : std_logic;
signal \nx.n1403\ : std_logic;
signal \nx.bit_ctr_30\ : std_logic;
signal \nx.n48_adj_704\ : std_logic;
signal \nx.n1407\ : std_logic;
signal \nx.n1474\ : std_logic;
signal \nx.n1506_cascade_\ : std_logic;
signal \nx.n18_adj_632\ : std_logic;
signal \nx.n1475\ : std_logic;
signal \nx.n1408\ : std_logic;
signal \nx.n1401\ : std_logic;
signal \nx.n1468\ : std_logic;
signal \nx.n1472\ : std_logic;
signal \nx.n1405\ : std_logic;
signal \nx.n1473\ : std_logic;
signal \nx.n1406\ : std_logic;
signal neopxl_color_15 : std_logic;
signal \nx.n2700_cascade_\ : std_logic;
signal \nx.n2801_cascade_\ : std_logic;
signal \nx.n29_adj_607\ : std_logic;
signal \nx.n37_adj_608_cascade_\ : std_logic;
signal \nx.n40_adj_609\ : std_logic;
signal \nx.n42_cascade_\ : std_logic;
signal \nx.n2720_cascade_\ : std_logic;
signal \nx.n2797_cascade_\ : std_logic;
signal \bfn_6_21_0_\ : std_logic;
signal \nx.n2809\ : std_logic;
signal \nx.n2876\ : std_logic;
signal \nx.n10813\ : std_logic;
signal \nx.n2808\ : std_logic;
signal \nx.n2875\ : std_logic;
signal \nx.n10814\ : std_logic;
signal \nx.n2807\ : std_logic;
signal \nx.n2874\ : std_logic;
signal \nx.n10815\ : std_logic;
signal \nx.n10816\ : std_logic;
signal \nx.n2805\ : std_logic;
signal \nx.n2872\ : std_logic;
signal \nx.n10817\ : std_logic;
signal \nx.n10818\ : std_logic;
signal \nx.n10819\ : std_logic;
signal \nx.n10820\ : std_logic;
signal \nx.n2802\ : std_logic;
signal \nx.n2869\ : std_logic;
signal \bfn_6_22_0_\ : std_logic;
signal \nx.n10821\ : std_logic;
signal \nx.n2800\ : std_logic;
signal \nx.n2867\ : std_logic;
signal \nx.n10822\ : std_logic;
signal \nx.n2799\ : std_logic;
signal \nx.n2866\ : std_logic;
signal \nx.n10823\ : std_logic;
signal \nx.n2798\ : std_logic;
signal \nx.n2865\ : std_logic;
signal \nx.n10824\ : std_logic;
signal \nx.n2797\ : std_logic;
signal \nx.n2864\ : std_logic;
signal \nx.n10825\ : std_logic;
signal \nx.n10826\ : std_logic;
signal \nx.n2795\ : std_logic;
signal \nx.n2862\ : std_logic;
signal \nx.n10827\ : std_logic;
signal \nx.n10828\ : std_logic;
signal \bfn_6_23_0_\ : std_logic;
signal \nx.n10829\ : std_logic;
signal \nx.n10830\ : std_logic;
signal \nx.n10831\ : std_logic;
signal \nx.n10832\ : std_logic;
signal \nx.n10833\ : std_logic;
signal \nx.n10834\ : std_logic;
signal \nx.n10835\ : std_logic;
signal \nx.n10836\ : std_logic;
signal \bfn_6_24_0_\ : std_logic;
signal \nx.n2885\ : std_logic;
signal \nx.n2858\ : std_logic;
signal \nx.n2791_cascade_\ : std_logic;
signal \nx.n2859\ : std_logic;
signal \nx.n2891\ : std_logic;
signal \nx.n2856\ : std_logic;
signal \nx.n2789_cascade_\ : std_logic;
signal \nx.n2995\ : std_logic;
signal \nx.n3062\ : std_logic;
signal \nx.n3017\ : std_logic;
signal \nx.n3094\ : std_logic;
signal \nx.n28_adj_660_cascade_\ : std_logic;
signal \nx.n16\ : std_logic;
signal \nx.n1928_cascade_\ : std_logic;
signal \nx.n1908_cascade_\ : std_logic;
signal \nx.n24_adj_648\ : std_logic;
signal \nx.n1877\ : std_logic;
signal \nx.n1829_cascade_\ : std_logic;
signal \nx.n1906_cascade_\ : std_logic;
signal \nx.n22_adj_605\ : std_logic;
signal \nx.n1006\ : std_logic;
signal \nx.n1804_cascade_\ : std_logic;
signal \nx.n19_cascade_\ : std_logic;
signal \nx.n26_adj_600\ : std_logic;
signal \nx.bit_ctr_27\ : std_logic;
signal \nx.bit_ctr_28\ : std_logic;
signal \nx.n739\ : std_logic;
signal \nx.bit_ctr_26\ : std_logic;
signal \nx.n977\ : std_logic;
signal \bfn_6_28_0_\ : std_logic;
signal \nx.n7082\ : std_logic;
signal \nx.n976\ : std_logic;
signal \nx.n10474\ : std_logic;
signal \nx.n7342\ : std_logic;
signal \nx.n975\ : std_logic;
signal \nx.n10475\ : std_logic;
signal \nx.n974\ : std_logic;
signal \nx.n10476\ : std_logic;
signal \nx.n906\ : std_logic;
signal \nx.n973\ : std_logic;
signal \nx.n10477\ : std_logic;
signal \nx.n13064\ : std_logic;
signal \nx.n10478\ : std_logic;
signal \nx.n4_adj_596\ : std_logic;
signal \nx.n5260\ : std_logic;
signal \nx.n11559\ : std_logic;
signal \nx.n838\ : std_logic;
signal \nx.n11674\ : std_logic;
signal \nx.n20_adj_634\ : std_logic;
signal \nx.n1532_cascade_\ : std_logic;
signal \nx.n1606_cascade_\ : std_logic;
signal \nx.n22_adj_647_cascade_\ : std_logic;
signal \nx.n1631_cascade_\ : std_logic;
signal \nx.n19_adj_602\ : std_logic;
signal \nx.n1409\ : std_logic;
signal \nx.n1476\ : std_logic;
signal \nx.n1433\ : std_logic;
signal \nx.n1508_cascade_\ : std_logic;
signal \nx.n16_adj_633\ : std_logic;
signal \nx.n1599_cascade_\ : std_logic;
signal \bfn_6_31_0_\ : std_logic;
signal \nx.n10592\ : std_logic;
signal \nx.n1508\ : std_logic;
signal \nx.n1575\ : std_logic;
signal \nx.n10593\ : std_logic;
signal \nx.n1507\ : std_logic;
signal \nx.n1574\ : std_logic;
signal \nx.n10594\ : std_logic;
signal \nx.n10595\ : std_logic;
signal \nx.n1505\ : std_logic;
signal \nx.n1572\ : std_logic;
signal \nx.n10596\ : std_logic;
signal \nx.n1504\ : std_logic;
signal \nx.n1571\ : std_logic;
signal \nx.n10597\ : std_logic;
signal \nx.n10598\ : std_logic;
signal \nx.n10599\ : std_logic;
signal \nx.n1502\ : std_logic;
signal \nx.n1569\ : std_logic;
signal \bfn_6_32_0_\ : std_logic;
signal \nx.n1501\ : std_logic;
signal \nx.n1568\ : std_logic;
signal \nx.n10600\ : std_logic;
signal \nx.n1500\ : std_logic;
signal \nx.n1567\ : std_logic;
signal \nx.n10601\ : std_logic;
signal \nx.n1499\ : std_logic;
signal \nx.n10602\ : std_logic;
signal neopxl_color_13 : std_logic;
signal n11683 : std_logic;
signal timer_0 : std_logic;
signal neo_pixel_transmitter_t0_0 : std_logic;
signal \nx.n33_adj_652\ : std_logic;
signal pin_out_0 : std_logic;
signal pin_out_1 : std_logic;
signal \nx.bit_ctr_8\ : std_logic;
signal \nx.n2777\ : std_logic;
signal \bfn_7_19_0_\ : std_logic;
signal \nx.n2776\ : std_logic;
signal \nx.n10790\ : std_logic;
signal \nx.n2708\ : std_logic;
signal \nx.n2775\ : std_logic;
signal \nx.n10791\ : std_logic;
signal \nx.n2707\ : std_logic;
signal \nx.n2774\ : std_logic;
signal \nx.n10792\ : std_logic;
signal \nx.n2706\ : std_logic;
signal \nx.n2773\ : std_logic;
signal \nx.n10793\ : std_logic;
signal \nx.n10794\ : std_logic;
signal \nx.n2771\ : std_logic;
signal \nx.n10795\ : std_logic;
signal \nx.n2770\ : std_logic;
signal \nx.n10796\ : std_logic;
signal \nx.n10797\ : std_logic;
signal \nx.n2702\ : std_logic;
signal \nx.n2769\ : std_logic;
signal \bfn_7_20_0_\ : std_logic;
signal \nx.n2768\ : std_logic;
signal \nx.n10798\ : std_logic;
signal \nx.n2700\ : std_logic;
signal \nx.n2767\ : std_logic;
signal \nx.n10799\ : std_logic;
signal \nx.n2766\ : std_logic;
signal \nx.n10800\ : std_logic;
signal \nx.n2765\ : std_logic;
signal \nx.n10801\ : std_logic;
signal \nx.n2764\ : std_logic;
signal \nx.n10802\ : std_logic;
signal \nx.n2696\ : std_logic;
signal \nx.n2763\ : std_logic;
signal \nx.n10803\ : std_logic;
signal \nx.n2762\ : std_logic;
signal \nx.n10804\ : std_logic;
signal \nx.n10805\ : std_logic;
signal \bfn_7_21_0_\ : std_logic;
signal \nx.n10806\ : std_logic;
signal \nx.n2759\ : std_logic;
signal \nx.n10807\ : std_logic;
signal \nx.n10808\ : std_logic;
signal \nx.n2757\ : std_logic;
signal \nx.n10809\ : std_logic;
signal \nx.n2756\ : std_logic;
signal \nx.n10810\ : std_logic;
signal \nx.n10811\ : std_logic;
signal \nx.n10812\ : std_logic;
signal neo_pixel_transmitter_t0_22 : std_logic;
signal \nx.n11\ : std_logic;
signal \nx.n2761\ : std_logic;
signal \nx.n2860\ : std_logic;
signal \nx.n2793_cascade_\ : std_logic;
signal \nx.n2892\ : std_logic;
signal \nx.n2758\ : std_logic;
signal \nx.n2760\ : std_logic;
signal \nx.n2873\ : std_logic;
signal \nx.n2806\ : std_logic;
signal \nx.n2905\ : std_logic;
signal \nx.n2793\ : std_logic;
signal \nx.n2791\ : std_logic;
signal \nx.n2792\ : std_logic;
signal \nx.n2786\ : std_logic;
signal \nx.n38_adj_625_cascade_\ : std_logic;
signal \nx.n42_adj_635\ : std_logic;
signal \nx.n41_adj_643\ : std_logic;
signal \nx.n43_cascade_\ : std_logic;
signal \nx.n44\ : std_logic;
signal \nx.n2854\ : std_logic;
signal \nx.n2819_cascade_\ : std_logic;
signal \nx.n2886\ : std_logic;
signal \nx.n2789\ : std_logic;
signal \nx.n26_adj_615\ : std_logic;
signal \nx.n2863\ : std_logic;
signal \nx.n2796\ : std_logic;
signal \nx.n2895\ : std_logic;
signal \nx.n2877\ : std_logic;
signal \nx.bit_ctr_7\ : std_logic;
signal \nx.n2909\ : std_logic;
signal \nx.n2868\ : std_logic;
signal \nx.n2801\ : std_logic;
signal \nx.n2900\ : std_logic;
signal \nx.n2861\ : std_logic;
signal \nx.n2794\ : std_logic;
signal \nx.n2893\ : std_logic;
signal \nx.n2788\ : std_logic;
signal \nx.n2855\ : std_logic;
signal \nx.n2887\ : std_logic;
signal \nx.n2890\ : std_logic;
signal \nx.n2888\ : std_logic;
signal \nx.n2887_cascade_\ : std_logic;
signal \nx.n39_adj_679\ : std_logic;
signal \nx.n2803\ : std_logic;
signal \nx.n2870\ : std_logic;
signal \nx.n2902\ : std_logic;
signal \nx.n2871\ : std_logic;
signal \nx.n2903\ : std_logic;
signal \nx.n2790\ : std_logic;
signal \nx.n2819\ : std_logic;
signal \nx.n2857\ : std_logic;
signal \nx.n2889\ : std_logic;
signal \nx.bit_ctr_16\ : std_logic;
signal \bfn_7_25_0_\ : std_logic;
signal \nx.n1909\ : std_logic;
signal \nx.n13435\ : std_logic;
signal \nx.n10642\ : std_logic;
signal \nx.n1908\ : std_logic;
signal \nx.n10643\ : std_logic;
signal \nx.n1907\ : std_logic;
signal \nx.n10644\ : std_logic;
signal \nx.n1906\ : std_logic;
signal \nx.n10645\ : std_logic;
signal \nx.n10646\ : std_logic;
signal \nx.n1904\ : std_logic;
signal \nx.n10647\ : std_logic;
signal \nx.n1903\ : std_logic;
signal \nx.n10648\ : std_logic;
signal \nx.n10649\ : std_logic;
signal \bfn_7_26_0_\ : std_logic;
signal \nx.n10650\ : std_logic;
signal \nx.n10651\ : std_logic;
signal \nx.n1899\ : std_logic;
signal \nx.n10652\ : std_logic;
signal \nx.n10653\ : std_logic;
signal \nx.n10654\ : std_logic;
signal \nx.n10655\ : std_logic;
signal \nx.n1928\ : std_logic;
signal \nx.n10656\ : std_logic;
signal \nx.n1897\ : std_logic;
signal \nx.n1902\ : std_logic;
signal \nx.n10994\ : std_logic;
signal \nx.n13425\ : std_logic;
signal \nx.n1701_cascade_\ : std_logic;
signal \nx.n1801_cascade_\ : std_logic;
signal \nx.n23\ : std_logic;
signal \nx.n1577\ : std_logic;
signal \nx.bit_ctr_20\ : std_logic;
signal \nx.n1609_cascade_\ : std_logic;
signal \nx.n16_adj_646\ : std_logic;
signal \nx.n1570\ : std_logic;
signal \nx.n1503\ : std_logic;
signal \nx.bit_ctr_19\ : std_logic;
signal \nx.n1677\ : std_logic;
signal \bfn_7_30_0_\ : std_logic;
signal \nx.n1609\ : std_logic;
signal \nx.n1676\ : std_logic;
signal \nx.n10603\ : std_logic;
signal \nx.n10604\ : std_logic;
signal \nx.n1607\ : std_logic;
signal \nx.n1674\ : std_logic;
signal \nx.n10605\ : std_logic;
signal \nx.n10606\ : std_logic;
signal \nx.n1672\ : std_logic;
signal \nx.n10607\ : std_logic;
signal \nx.n10608\ : std_logic;
signal \nx.n1603\ : std_logic;
signal \nx.n1670\ : std_logic;
signal \nx.n10609\ : std_logic;
signal \nx.n10610\ : std_logic;
signal \nx.n1602\ : std_logic;
signal \nx.n1669\ : std_logic;
signal \bfn_7_31_0_\ : std_logic;
signal \nx.n10611\ : std_logic;
signal \nx.n10612\ : std_logic;
signal \nx.n1599\ : std_logic;
signal \nx.n1666\ : std_logic;
signal \nx.n10613\ : std_logic;
signal \nx.n1598\ : std_logic;
signal \nx.n10614\ : std_logic;
signal \nx.n1600\ : std_logic;
signal \nx.n1667\ : std_logic;
signal \n7258_cascade_\ : std_logic;
signal n7236 : std_logic;
signal \n7270_cascade_\ : std_logic;
signal n7254 : std_logic;
signal pin_out_5 : std_logic;
signal \n13152_cascade_\ : std_logic;
signal n13146 : std_logic;
signal \n13462_cascade_\ : std_logic;
signal n13153 : std_logic;
signal pin_out_3 : std_logic;
signal pin_out_2 : std_logic;
signal n13147 : std_logic;
signal n13168 : std_logic;
signal \n13167_cascade_\ : std_logic;
signal n13450 : std_logic;
signal \nx.n2694\ : std_logic;
signal \nx.n2697\ : std_logic;
signal \nx.n2704\ : std_logic;
signal \nx.n2695\ : std_logic;
signal \nx.n2698\ : std_logic;
signal \nx.n2698_cascade_\ : std_logic;
signal \nx.n39_adj_610\ : std_logic;
signal \nx.n2703\ : std_logic;
signal \nx.n2709\ : std_logic;
signal \nx.n2592_cascade_\ : std_logic;
signal \nx.n2689\ : std_logic;
signal \nx.n2690\ : std_logic;
signal \nx.n2689_cascade_\ : std_logic;
signal \nx.n2691\ : std_logic;
signal \nx.n2701\ : std_logic;
signal \nx.n2105_cascade_\ : std_logic;
signal \nx.n2595_cascade_\ : std_logic;
signal \nx.n28_adj_663\ : std_logic;
signal \nx.n26_adj_664_cascade_\ : std_logic;
signal \nx.n25_adj_666\ : std_logic;
signal \nx.n2027_cascade_\ : std_logic;
signal \nx.n2099_cascade_\ : std_logic;
signal \nx.n2904\ : std_logic;
signal \nx.n2971\ : std_logic;
signal \nx.n2918\ : std_logic;
signal \nx.n3003\ : std_logic;
signal \bfn_9_23_0_\ : std_logic;
signal \nx.n10657\ : std_logic;
signal \nx.n10658\ : std_logic;
signal \nx.n10659\ : std_logic;
signal \nx.n2006\ : std_logic;
signal \nx.n2073\ : std_logic;
signal \nx.n10660\ : std_logic;
signal \nx.n2005\ : std_logic;
signal \nx.n2072\ : std_logic;
signal \nx.n10661\ : std_logic;
signal \nx.n2004\ : std_logic;
signal \nx.n2071\ : std_logic;
signal \nx.n10662\ : std_logic;
signal \nx.n10663\ : std_logic;
signal \nx.n10664\ : std_logic;
signal \bfn_9_24_0_\ : std_logic;
signal \nx.n2001\ : std_logic;
signal \nx.n2068\ : std_logic;
signal \nx.n10665\ : std_logic;
signal \nx.n2000\ : std_logic;
signal \nx.n2067\ : std_logic;
signal \nx.n10666\ : std_logic;
signal \nx.n1999\ : std_logic;
signal \nx.n2066\ : std_logic;
signal \nx.n10667\ : std_logic;
signal \nx.n10668\ : std_logic;
signal \nx.n10669\ : std_logic;
signal \nx.n1996\ : std_logic;
signal \nx.n2063\ : std_logic;
signal \nx.n10670\ : std_logic;
signal \nx.n10671\ : std_logic;
signal \nx.n10672\ : std_logic;
signal \nx.n1994\ : std_logic;
signal \bfn_9_25_0_\ : std_logic;
signal \nx.n1901\ : std_logic;
signal \nx.n1905\ : std_logic;
signal \nx.n25_adj_606\ : std_logic;
signal \nx.n22\ : std_logic;
signal \nx.n1900\ : std_logic;
signal \nx.n1799_cascade_\ : std_logic;
signal \nx.n1898\ : std_logic;
signal \nx.n1797_cascade_\ : std_logic;
signal \nx.n1896\ : std_logic;
signal \nx.bit_ctr_17\ : std_logic;
signal \nx.bit_ctr_22\ : std_logic;
signal \nx.n30_adj_703\ : std_logic;
signal \bfn_9_27_0_\ : std_logic;
signal \nx.n1809\ : std_logic;
signal \nx.n1876\ : std_logic;
signal \nx.n10628\ : std_logic;
signal \nx.n1808\ : std_logic;
signal \nx.n1875\ : std_logic;
signal \nx.n10629\ : std_logic;
signal \nx.n1807\ : std_logic;
signal \nx.n1874\ : std_logic;
signal \nx.n10630\ : std_logic;
signal \nx.n1873\ : std_logic;
signal \nx.n10631\ : std_logic;
signal \nx.n1805\ : std_logic;
signal \nx.n1872\ : std_logic;
signal \nx.n10632\ : std_logic;
signal \nx.n1804\ : std_logic;
signal \nx.n1871\ : std_logic;
signal \nx.n10633\ : std_logic;
signal \nx.n1870\ : std_logic;
signal \nx.n10634\ : std_logic;
signal \nx.n10635\ : std_logic;
signal \nx.n1869\ : std_logic;
signal \bfn_9_28_0_\ : std_logic;
signal \nx.n1801\ : std_logic;
signal \nx.n1868\ : std_logic;
signal \nx.n10636\ : std_logic;
signal \nx.n1800\ : std_logic;
signal \nx.n1867\ : std_logic;
signal \nx.n10637\ : std_logic;
signal \nx.n1799\ : std_logic;
signal \nx.n1866\ : std_logic;
signal \nx.n10638\ : std_logic;
signal \nx.n1865\ : std_logic;
signal \nx.n10639\ : std_logic;
signal \nx.n1797\ : std_logic;
signal \nx.n1864\ : std_logic;
signal \nx.n10640\ : std_logic;
signal \nx.n1829\ : std_logic;
signal \nx.n10641\ : std_logic;
signal \nx.n1895\ : std_logic;
signal \nx.n1668\ : std_logic;
signal \nx.n1601\ : std_logic;
signal \nx.n1509\ : std_logic;
signal \nx.n1576\ : std_logic;
signal \nx.n1608_cascade_\ : std_logic;
signal \nx.n18\ : std_logic;
signal \nx.n1506\ : std_logic;
signal \nx.n1573\ : std_logic;
signal \nx.n1532\ : std_logic;
signal \nx.n1605\ : std_logic;
signal \nx.n1604\ : std_logic;
signal \nx.n1671\ : std_logic;
signal \nx.n1606\ : std_logic;
signal \nx.n1673\ : std_logic;
signal \n21_cascade_\ : std_logic;
signal n6150 : std_logic;
signal pin_out_6 : std_logic;
signal n7262 : std_logic;
signal pin_out_7 : std_logic;
signal n8_adj_780 : std_logic;
signal \n8_adj_780_cascade_\ : std_logic;
signal n7274 : std_logic;
signal \nx.n2677\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \nx.n2676\ : std_logic;
signal \nx.n10768\ : std_logic;
signal \nx.n2675\ : std_logic;
signal \nx.n10769\ : std_logic;
signal \nx.n2674\ : std_logic;
signal \nx.n10770\ : std_logic;
signal \nx.n10771\ : std_logic;
signal \nx.n2672\ : std_logic;
signal \nx.n10772\ : std_logic;
signal \nx.n2671\ : std_logic;
signal \nx.n10773\ : std_logic;
signal \nx.n2670\ : std_logic;
signal \nx.n10774\ : std_logic;
signal \nx.n10775\ : std_logic;
signal \nx.n2669\ : std_logic;
signal \bfn_10_18_0_\ : std_logic;
signal \nx.n2668\ : std_logic;
signal \nx.n10776\ : std_logic;
signal \nx.n10777\ : std_logic;
signal \nx.n2666\ : std_logic;
signal \nx.n10778\ : std_logic;
signal \nx.n2665\ : std_logic;
signal \nx.n10779\ : std_logic;
signal \nx.n2664\ : std_logic;
signal \nx.n10780\ : std_logic;
signal \nx.n2663\ : std_logic;
signal \nx.n10781\ : std_logic;
signal \nx.n2595\ : std_logic;
signal \nx.n2662\ : std_logic;
signal \nx.n10782\ : std_logic;
signal \nx.n10783\ : std_logic;
signal \bfn_10_19_0_\ : std_logic;
signal \nx.n10784\ : std_logic;
signal \nx.n2592\ : std_logic;
signal \nx.n2659\ : std_logic;
signal \nx.n10785\ : std_logic;
signal \nx.n2658\ : std_logic;
signal \nx.n10786\ : std_logic;
signal \nx.n2657\ : std_logic;
signal \nx.n10787\ : std_logic;
signal \nx.n10788\ : std_logic;
signal \nx.n10789\ : std_logic;
signal \nx.n2660\ : std_logic;
signal \nx.n2692\ : std_logic;
signal \nx.n34_adj_603_cascade_\ : std_logic;
signal \nx.n39_cascade_\ : std_logic;
signal \nx.n2621_cascade_\ : std_logic;
signal \nx.n2661\ : std_logic;
signal \nx.n2693\ : std_logic;
signal \nx.n2667\ : std_logic;
signal \nx.n2699\ : std_logic;
signal \nx.n2687\ : std_logic;
signal \nx.n2699_cascade_\ : std_logic;
signal \nx.n36\ : std_logic;
signal \nx.n41\ : std_logic;
signal \nx.n2656\ : std_logic;
signal \nx.n31_adj_655_cascade_\ : std_logic;
signal \nx.n24_adj_654\ : std_logic;
signal \nx.n36_adj_656_cascade_\ : std_logic;
signal \nx.n33_adj_659\ : std_logic;
signal \nx.n2423_cascade_\ : std_logic;
signal \nx.n2491_cascade_\ : std_logic;
signal \nx.n2394_cascade_\ : std_logic;
signal \nx.n2077\ : std_logic;
signal \nx.n2070\ : std_logic;
signal \nx.n2069\ : std_logic;
signal \nx.n2076\ : std_logic;
signal \nx.bit_ctr_15\ : std_logic;
signal \nx.n2003\ : std_logic;
signal \nx.n2009\ : std_logic;
signal \nx.n27_adj_665\ : std_logic;
signal \nx.n2074\ : std_logic;
signal \nx.n2064\ : std_logic;
signal \nx.n1997\ : std_logic;
signal \nx.n2062\ : std_logic;
signal \nx.n1995\ : std_logic;
signal \nx.n26_adj_667\ : std_logic;
signal \nx.n30_adj_668_cascade_\ : std_logic;
signal \nx.n28_adj_669\ : std_logic;
signal \nx.n2008\ : std_logic;
signal \nx.n2075\ : std_logic;
signal \nx.n2107_cascade_\ : std_logic;
signal \nx.n29_adj_670\ : std_logic;
signal \nx.n2065\ : std_logic;
signal \nx.n1998\ : std_logic;
signal \nx.n2027\ : std_logic;
signal \nx.n2097_cascade_\ : std_logic;
signal \nx.n27_adj_671\ : std_logic;
signal \nx.n2007\ : std_logic;
signal \nx.n2002\ : std_logic;
signal \nx.n22_adj_662\ : std_logic;
signal \nx.n1803\ : std_logic;
signal \nx.n22_adj_673_cascade_\ : std_logic;
signal \nx.n16_adj_672\ : std_logic;
signal \nx.n1798\ : std_logic;
signal \nx.n1608\ : std_logic;
signal \nx.n1675\ : std_logic;
signal \nx.n1631\ : std_logic;
signal \nx.n1707_cascade_\ : std_logic;
signal \nx.n1806\ : std_logic;
signal \nx.n20_adj_680\ : std_logic;
signal \nx.n24_adj_685\ : std_logic;
signal \nx.n1730_cascade_\ : std_logic;
signal \nx.n1802\ : std_logic;
signal \nx.bit_ctr_18\ : std_logic;
signal \nx.n1777\ : std_logic;
signal \bfn_10_28_0_\ : std_logic;
signal \nx.n1709\ : std_logic;
signal \nx.n1776\ : std_logic;
signal \nx.n10615\ : std_logic;
signal \nx.n1708\ : std_logic;
signal \nx.n1775\ : std_logic;
signal \nx.n10616\ : std_logic;
signal \nx.n1707\ : std_logic;
signal \nx.n1774\ : std_logic;
signal \nx.n10617\ : std_logic;
signal \nx.n1706\ : std_logic;
signal \nx.n1773\ : std_logic;
signal \nx.n10618\ : std_logic;
signal \nx.n1705\ : std_logic;
signal \nx.n1772\ : std_logic;
signal \nx.n10619\ : std_logic;
signal \nx.n1704\ : std_logic;
signal \nx.n1771\ : std_logic;
signal \nx.n10620\ : std_logic;
signal \nx.n1703\ : std_logic;
signal \nx.n1770\ : std_logic;
signal \nx.n10621\ : std_logic;
signal \nx.n10622\ : std_logic;
signal \nx.n1702\ : std_logic;
signal \nx.n1769\ : std_logic;
signal \bfn_10_29_0_\ : std_logic;
signal \nx.n1701\ : std_logic;
signal \nx.n1768\ : std_logic;
signal \nx.n10623\ : std_logic;
signal \nx.n1700\ : std_logic;
signal \nx.n1767\ : std_logic;
signal \nx.n10624\ : std_logic;
signal \nx.n1699\ : std_logic;
signal \nx.n1766\ : std_logic;
signal \nx.n10625\ : std_logic;
signal \nx.n1698\ : std_logic;
signal \nx.n1765\ : std_logic;
signal \nx.n10626\ : std_logic;
signal \nx.n1730\ : std_logic;
signal \nx.n1697\ : std_logic;
signal \nx.n10627\ : std_logic;
signal \nx.n1796\ : std_logic;
signal pin_oe_22 : std_logic;
signal n6158 : std_logic;
signal n8 : std_logic;
signal \n22_adj_740_cascade_\ : std_logic;
signal n5907 : std_logic;
signal n6162 : std_logic;
signal \n6162_cascade_\ : std_logic;
signal n7278 : std_logic;
signal n6156 : std_logic;
signal \n7266_cascade_\ : std_logic;
signal pin_out_4 : std_logic;
signal \nx.n2609\ : std_logic;
signal \nx.bit_ctr_9\ : std_logic;
signal \nx.n2609_cascade_\ : std_logic;
signal \nx.n28_adj_599_cascade_\ : std_logic;
signal \nx.n35\ : std_logic;
signal \nx.n40\ : std_logic;
signal \nx.n2608\ : std_logic;
signal \nx.n2596\ : std_logic;
signal \nx.n2599\ : std_logic;
signal \nx.n2596_cascade_\ : std_logic;
signal \nx.n2604\ : std_logic;
signal \nx.n37\ : std_logic;
signal \nx.n2598\ : std_logic;
signal \nx.n38\ : std_logic;
signal \nx.n2602\ : std_logic;
signal \nx.n2606\ : std_logic;
signal \nx.n2673\ : std_logic;
signal \nx.n2606_cascade_\ : std_logic;
signal \nx.n2621\ : std_logic;
signal \nx.n2705\ : std_logic;
signal \nx.n2772\ : std_logic;
signal \nx.n2705_cascade_\ : std_logic;
signal \nx.n2804\ : std_logic;
signal \nx.n2594\ : std_logic;
signal \nx.n2504_cascade_\ : std_logic;
signal \nx.n2603\ : std_logic;
signal \nx.n2589\ : std_logic;
signal \nx.n2688\ : std_logic;
signal \nx.n2720\ : std_logic;
signal \nx.n2755\ : std_logic;
signal \nx.n2787\ : std_logic;
signal \nx.n2590\ : std_logic;
signal \nx.n2591\ : std_logic;
signal \nx.n2296_cascade_\ : std_logic;
signal \nx.n2395_cascade_\ : std_logic;
signal \nx.n2494_cascade_\ : std_logic;
signal \nx.n2593\ : std_logic;
signal \nx.n2293_cascade_\ : std_logic;
signal \nx.bit_ctr_14\ : std_logic;
signal \bfn_11_23_0_\ : std_logic;
signal \nx.n2109\ : std_logic;
signal \nx.n13436\ : std_logic;
signal \nx.n10673\ : std_logic;
signal \nx.n2108\ : std_logic;
signal \nx.n10674\ : std_logic;
signal \nx.n2107\ : std_logic;
signal \nx.n10675\ : std_logic;
signal \nx.n2106\ : std_logic;
signal \nx.n10676\ : std_logic;
signal \nx.n2105\ : std_logic;
signal \nx.n10677\ : std_logic;
signal \nx.n2104\ : std_logic;
signal \nx.n10678\ : std_logic;
signal \nx.n2103\ : std_logic;
signal \nx.n10679\ : std_logic;
signal \nx.n10680\ : std_logic;
signal \nx.n2102\ : std_logic;
signal \bfn_11_24_0_\ : std_logic;
signal \nx.n2101\ : std_logic;
signal \nx.n10681\ : std_logic;
signal \nx.n2100\ : std_logic;
signal \nx.n10682\ : std_logic;
signal \nx.n2099\ : std_logic;
signal \nx.n10683\ : std_logic;
signal \nx.n2098\ : std_logic;
signal \nx.n10684\ : std_logic;
signal \nx.n2097\ : std_logic;
signal \nx.n10685\ : std_logic;
signal \nx.n2096\ : std_logic;
signal \nx.n10686\ : std_logic;
signal \nx.n2095\ : std_logic;
signal \nx.n10687\ : std_logic;
signal \nx.n10688\ : std_logic;
signal \nx.n2094\ : std_logic;
signal \bfn_11_25_0_\ : std_logic;
signal \nx.n2093\ : std_logic;
signal \nx.n2126\ : std_logic;
signal \nx.n10689\ : std_logic;
signal n12171 : std_logic;
signal n6_adj_761 : std_logic;
signal \n15_cascade_\ : std_logic;
signal n14 : std_logic;
signal n12091 : std_logic;
signal \n24_adj_720_cascade_\ : std_logic;
signal n11898 : std_logic;
signal neopxl_color_7 : std_logic;
signal n22_adj_724 : std_logic;
signal n17_adj_765 : std_logic;
signal \n16_adj_764_cascade_\ : std_logic;
signal n10978 : std_logic;
signal n36 : std_logic;
signal \n7166_cascade_\ : std_logic;
signal n6152 : std_logic;
signal \n8_adj_751_cascade_\ : std_logic;
signal \n7294_cascade_\ : std_logic;
signal pin_out_11 : std_logic;
signal n6154 : std_logic;
signal n8_adj_744 : std_logic;
signal \n13048_cascade_\ : std_logic;
signal n13264 : std_logic;
signal \nx.n2597\ : std_logic;
signal \nx.n2601\ : std_logic;
signal \nx.n2497_cascade_\ : std_logic;
signal \nx.n26_adj_611_cascade_\ : std_logic;
signal \nx.n33\ : std_logic;
signal \nx.n38_adj_612_cascade_\ : std_logic;
signal \nx.n2522_cascade_\ : std_logic;
signal \nx.n2600\ : std_logic;
signal \nx.n2605\ : std_logic;
signal \nx.n35_adj_639\ : std_logic;
signal \nx.bit_ctr_10\ : std_logic;
signal \nx.n2577\ : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal \nx.n2509\ : std_logic;
signal \nx.n2576\ : std_logic;
signal \nx.n10747\ : std_logic;
signal \nx.n10748\ : std_logic;
signal \nx.n2574\ : std_logic;
signal \nx.n10749\ : std_logic;
signal \nx.n2573\ : std_logic;
signal \nx.n10750\ : std_logic;
signal \nx.n2505\ : std_logic;
signal \nx.n2572\ : std_logic;
signal \nx.n10751\ : std_logic;
signal \nx.n2571\ : std_logic;
signal \nx.n10752\ : std_logic;
signal \nx.n2570\ : std_logic;
signal \nx.n10753\ : std_logic;
signal \nx.n10754\ : std_logic;
signal \nx.n2569\ : std_logic;
signal \bfn_12_21_0_\ : std_logic;
signal \nx.n2501\ : std_logic;
signal \nx.n2568\ : std_logic;
signal \nx.n10755\ : std_logic;
signal \nx.n2567\ : std_logic;
signal \nx.n10756\ : std_logic;
signal \nx.n2499\ : std_logic;
signal \nx.n2566\ : std_logic;
signal \nx.n10757\ : std_logic;
signal \nx.n2565\ : std_logic;
signal \nx.n10758\ : std_logic;
signal \nx.n2497\ : std_logic;
signal \nx.n2564\ : std_logic;
signal \nx.n10759\ : std_logic;
signal \nx.n2496\ : std_logic;
signal \nx.n2563\ : std_logic;
signal \nx.n10760\ : std_logic;
signal \nx.n2562\ : std_logic;
signal \nx.n10761\ : std_logic;
signal \nx.n10762\ : std_logic;
signal \nx.n2494\ : std_logic;
signal \nx.n2561\ : std_logic;
signal \bfn_12_22_0_\ : std_logic;
signal \nx.n2493\ : std_logic;
signal \nx.n2560\ : std_logic;
signal \nx.n10763\ : std_logic;
signal \nx.n2492\ : std_logic;
signal \nx.n2559\ : std_logic;
signal \nx.n10764\ : std_logic;
signal \nx.n2491\ : std_logic;
signal \nx.n2558\ : std_logic;
signal \nx.n10765\ : std_logic;
signal \nx.n2557\ : std_logic;
signal \nx.n10766\ : std_logic;
signal \nx.n10767\ : std_logic;
signal \nx.n2588\ : std_logic;
signal \nx.n30_adj_640\ : std_logic;
signal \nx.n34_cascade_\ : std_logic;
signal \nx.n21\ : std_logic;
signal \nx.n2225_cascade_\ : std_logic;
signal \nx.n31\ : std_logic;
signal \nx.n28_adj_601\ : std_logic;
signal neopxl_color_12 : std_logic;
signal neopxl_color_prev_12 : std_logic;
signal \nx.n30\ : std_logic;
signal \nx.n22_adj_604\ : std_logic;
signal delay_counter_0 : std_logic;
signal \bfn_12_26_0_\ : std_logic;
signal delay_counter_1 : std_logic;
signal n10517 : std_logic;
signal delay_counter_2 : std_logic;
signal n10518 : std_logic;
signal delay_counter_3 : std_logic;
signal n10519 : std_logic;
signal delay_counter_4 : std_logic;
signal n10520 : std_logic;
signal delay_counter_5 : std_logic;
signal n10521 : std_logic;
signal delay_counter_6 : std_logic;
signal n10522 : std_logic;
signal delay_counter_7 : std_logic;
signal n10523 : std_logic;
signal n10524 : std_logic;
signal delay_counter_8 : std_logic;
signal \bfn_12_27_0_\ : std_logic;
signal delay_counter_9 : std_logic;
signal n10525 : std_logic;
signal delay_counter_10 : std_logic;
signal n10526 : std_logic;
signal delay_counter_11 : std_logic;
signal n10527 : std_logic;
signal delay_counter_12 : std_logic;
signal n10528 : std_logic;
signal delay_counter_13 : std_logic;
signal n10529 : std_logic;
signal delay_counter_14 : std_logic;
signal n10530 : std_logic;
signal delay_counter_15 : std_logic;
signal n10531 : std_logic;
signal n10532 : std_logic;
signal delay_counter_16 : std_logic;
signal \bfn_12_28_0_\ : std_logic;
signal delay_counter_17 : std_logic;
signal n10533 : std_logic;
signal delay_counter_18 : std_logic;
signal n10534 : std_logic;
signal delay_counter_19 : std_logic;
signal n10535 : std_logic;
signal delay_counter_20 : std_logic;
signal n10536 : std_logic;
signal delay_counter_21 : std_logic;
signal n10537 : std_logic;
signal delay_counter_22 : std_logic;
signal n10538 : std_logic;
signal delay_counter_23 : std_logic;
signal n10539 : std_logic;
signal n10540 : std_logic;
signal delay_counter_24 : std_logic;
signal \bfn_12_29_0_\ : std_logic;
signal delay_counter_25 : std_logic;
signal n10541 : std_logic;
signal delay_counter_26 : std_logic;
signal n10542 : std_logic;
signal delay_counter_27 : std_logic;
signal n10543 : std_logic;
signal delay_counter_28 : std_logic;
signal n10544 : std_logic;
signal delay_counter_29 : std_logic;
signal n10545 : std_logic;
signal delay_counter_30 : std_logic;
signal n10546 : std_logic;
signal n10547 : std_logic;
signal n7442 : std_logic;
signal \n10_adj_779_cascade_\ : std_logic;
signal n10_adj_779 : std_logic;
signal \n7290_cascade_\ : std_logic;
signal pin_out_10 : std_logic;
signal n7135 : std_logic;
signal \n7155_cascade_\ : std_logic;
signal n6190 : std_logic;
signal \n6190_cascade_\ : std_logic;
signal n7334 : std_logic;
signal n6170 : std_logic;
signal n9415 : std_logic;
signal pin_in_8 : std_logic;
signal \n13480_cascade_\ : std_logic;
signal \current_pin_7__N_157_cascade_\ : std_logic;
signal pin_in_0 : std_logic;
signal pin_in_10 : std_logic;
signal \n2289_cascade_\ : std_logic;
signal pin_in_6 : std_logic;
signal n13453 : std_logic;
signal \n13364_cascade_\ : std_logic;
signal n150 : std_logic;
signal n13483 : std_logic;
signal n13360 : std_logic;
signal \nx.n2575\ : std_logic;
signal \nx.n2522\ : std_logic;
signal \nx.n2607\ : std_logic;
signal \nx.n2495\ : std_logic;
signal \nx.n2503\ : std_logic;
signal \nx.n2503_cascade_\ : std_logic;
signal \nx.n36_adj_636\ : std_logic;
signal \nx.n2502\ : std_logic;
signal \nx.n2508\ : std_logic;
signal \nx.n2506\ : std_logic;
signal neopxl_color_5 : std_logic;
signal n22_adj_730 : std_logic;
signal \nx.n2498\ : std_logic;
signal \nx.n2404_cascade_\ : std_logic;
signal \nx.n34_adj_657\ : std_logic;
signal \nx.n2490\ : std_logic;
signal \nx.n2504\ : std_logic;
signal \nx.n22_adj_637_cascade_\ : std_logic;
signal \nx.n2507\ : std_logic;
signal \nx.n37_adj_638\ : std_logic;
signal \nx.n2500\ : std_logic;
signal \nx.n2300_cascade_\ : std_logic;
signal \nx.n33_adj_644\ : std_logic;
signal \nx.n34_adj_641\ : std_logic;
signal \nx.n32_cascade_\ : std_logic;
signal \nx.n2324_cascade_\ : std_logic;
signal \nx.bit_ctr_13\ : std_logic;
signal \nx.n2277\ : std_logic;
signal \bfn_13_23_0_\ : std_logic;
signal \nx.n2209\ : std_logic;
signal \nx.n2276\ : std_logic;
signal \nx.n10690\ : std_logic;
signal \nx.n2208\ : std_logic;
signal \nx.n2275\ : std_logic;
signal \nx.n10691\ : std_logic;
signal \nx.n10692\ : std_logic;
signal \nx.n2206\ : std_logic;
signal \nx.n2273\ : std_logic;
signal \nx.n10693\ : std_logic;
signal \nx.n2205\ : std_logic;
signal \nx.n2272\ : std_logic;
signal \nx.n10694\ : std_logic;
signal \nx.n10695\ : std_logic;
signal \nx.n2203\ : std_logic;
signal \nx.n2270\ : std_logic;
signal \nx.n10696\ : std_logic;
signal \nx.n10697\ : std_logic;
signal \bfn_13_24_0_\ : std_logic;
signal \nx.n2201\ : std_logic;
signal \nx.n2268\ : std_logic;
signal \nx.n10698\ : std_logic;
signal \nx.n10699\ : std_logic;
signal \nx.n10700\ : std_logic;
signal \nx.n10701\ : std_logic;
signal \nx.n2197\ : std_logic;
signal \nx.n2264\ : std_logic;
signal \nx.n10702\ : std_logic;
signal \nx.n2196\ : std_logic;
signal \nx.n2263\ : std_logic;
signal \nx.n10703\ : std_logic;
signal \nx.n2195\ : std_logic;
signal \nx.n2262\ : std_logic;
signal \nx.n10704\ : std_logic;
signal \nx.n10705\ : std_logic;
signal \nx.n2194\ : std_logic;
signal \nx.n2261\ : std_logic;
signal \bfn_13_25_0_\ : std_logic;
signal \nx.n10706\ : std_logic;
signal \nx.n2192\ : std_logic;
signal \nx.n10707\ : std_logic;
signal n7155 : std_logic;
signal n6166 : std_logic;
signal \n6166_cascade_\ : std_logic;
signal n7286 : std_logic;
signal \n7_adj_753_cascade_\ : std_logic;
signal pin_in_2 : std_logic;
signal n22_adj_740 : std_logic;
signal \n21_adj_741_cascade_\ : std_logic;
signal n7128 : std_logic;
signal \n7150_cascade_\ : std_logic;
signal pin_in_11 : std_logic;
signal n2355 : std_logic;
signal n21_adj_714 : std_logic;
signal \n7_adj_719_cascade_\ : std_logic;
signal n7150 : std_logic;
signal pin_in_9 : std_logic;
signal n2337 : std_logic;
signal \n2343_cascade_\ : std_logic;
signal n2325 : std_logic;
signal pin_in_3 : std_logic;
signal pin_in_1 : std_logic;
signal n2361 : std_logic;
signal \n13474_cascade_\ : std_logic;
signal pin_in_12 : std_logic;
signal n13477 : std_logic;
signal pin_in_13 : std_logic;
signal pin_in_15 : std_logic;
signal n2367 : std_logic;
signal n33 : std_logic;
signal \n2379_cascade_\ : std_logic;
signal n45_adj_772 : std_logic;
signal neopxl_color_4 : std_logic;
signal n22_adj_732 : std_logic;
signal n7232 : std_logic;
signal n43 : std_logic;
signal n52_adj_770 : std_logic;
signal neopxl_color_6 : std_logic;
signal n22_adj_728 : std_logic;
signal \nx.bit_ctr_11\ : std_logic;
signal \nx.n2477\ : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal \nx.n2409\ : std_logic;
signal \nx.n2476\ : std_logic;
signal \nx.n10727\ : std_logic;
signal \nx.n2408\ : std_logic;
signal \nx.n2475\ : std_logic;
signal \nx.n10728\ : std_logic;
signal \nx.n2407\ : std_logic;
signal \nx.n2474\ : std_logic;
signal \nx.n10729\ : std_logic;
signal \nx.n2473\ : std_logic;
signal \nx.n10730\ : std_logic;
signal \nx.n2405\ : std_logic;
signal \nx.n2472\ : std_logic;
signal \nx.n10731\ : std_logic;
signal \nx.n2404\ : std_logic;
signal \nx.n2471\ : std_logic;
signal \nx.n10732\ : std_logic;
signal \nx.n2470\ : std_logic;
signal \nx.n10733\ : std_logic;
signal \nx.n10734\ : std_logic;
signal \nx.n2469\ : std_logic;
signal \bfn_14_22_0_\ : std_logic;
signal \nx.n2401\ : std_logic;
signal \nx.n2468\ : std_logic;
signal \nx.n10735\ : std_logic;
signal \nx.n2467\ : std_logic;
signal \nx.n10736\ : std_logic;
signal \nx.n2399\ : std_logic;
signal \nx.n2466\ : std_logic;
signal \nx.n10737\ : std_logic;
signal \nx.n2465\ : std_logic;
signal \nx.n10738\ : std_logic;
signal \nx.n2464\ : std_logic;
signal \nx.n10739\ : std_logic;
signal \nx.n2463\ : std_logic;
signal \nx.n10740\ : std_logic;
signal \nx.n2395\ : std_logic;
signal \nx.n2462\ : std_logic;
signal \nx.n10741\ : std_logic;
signal \nx.n10742\ : std_logic;
signal \nx.n2394\ : std_logic;
signal \nx.n2461\ : std_logic;
signal \bfn_14_23_0_\ : std_logic;
signal \nx.n2393\ : std_logic;
signal \nx.n2460\ : std_logic;
signal \nx.n10743\ : std_logic;
signal \nx.n2392\ : std_logic;
signal \nx.n2459\ : std_logic;
signal \nx.n10744\ : std_logic;
signal \nx.n2458\ : std_logic;
signal \nx.n10745\ : std_logic;
signal \nx.n2423\ : std_logic;
signal \nx.n10746\ : std_logic;
signal \nx.n2489\ : std_logic;
signal \nx.n2207\ : std_logic;
signal \nx.n2274\ : std_logic;
signal \nx.n2391\ : std_logic;
signal \nx.n2271\ : std_logic;
signal \nx.n2204\ : std_logic;
signal \nx.n2265\ : std_logic;
signal \nx.n2198\ : std_logic;
signal \nx.n2297_cascade_\ : std_logic;
signal \nx.n9650\ : std_logic;
signal \nx.n31_adj_645\ : std_logic;
signal \nx.n2269\ : std_logic;
signal \nx.n2202\ : std_logic;
signal \nx.n2267\ : std_logic;
signal \nx.n2200\ : std_logic;
signal \nx.n2266\ : std_logic;
signal \nx.n2199\ : std_logic;
signal \nx.n2260\ : std_logic;
signal \nx.n2193\ : std_logic;
signal \nx.n2225\ : std_logic;
signal \nx.n2396\ : std_logic;
signal \n13177_cascade_\ : std_logic;
signal \LED_c\ : std_logic;
signal n13176 : std_logic;
signal n21_adj_741 : std_logic;
signal n6172 : std_logic;
signal n7298 : std_logic;
signal \n6172_cascade_\ : std_logic;
signal n6174 : std_logic;
signal n7302 : std_logic;
signal n7_adj_753 : std_logic;
signal n6176 : std_logic;
signal \n7306_cascade_\ : std_logic;
signal pin_out_9 : std_logic;
signal n13162 : std_logic;
signal \n13161_cascade_\ : std_logic;
signal n8_adj_751 : std_logic;
signal n6164 : std_logic;
signal \n7282_cascade_\ : std_logic;
signal pin_out_8 : std_logic;
signal n6184 : std_logic;
signal \n7322_cascade_\ : std_logic;
signal n13471 : std_logic;
signal n13465 : std_logic;
signal n10_adj_736 : std_logic;
signal pin_in_14 : std_logic;
signal n7145 : std_logic;
signal n7314 : std_logic;
signal n6 : std_logic;
signal n6182 : std_logic;
signal \n7318_cascade_\ : std_logic;
signal n9_adj_733 : std_logic;
signal n6188 : std_logic;
signal n7330 : std_logic;
signal pin_out_18 : std_logic;
signal pin_out_16 : std_logic;
signal \n13438_cascade_\ : std_logic;
signal pin_out_17 : std_logic;
signal \n13441_cascade_\ : std_logic;
signal \n13142_cascade_\ : std_logic;
signal n13362 : std_logic;
signal \n149_cascade_\ : std_logic;
signal pin_out_19 : std_logic;
signal n8_adj_746 : std_logic;
signal n6186 : std_logic;
signal n7326 : std_logic;
signal n11_adj_734 : std_logic;
signal \n11_adj_734_cascade_\ : std_logic;
signal n36_adj_773 : std_logic;
signal pin_out_21 : std_logic;
signal pin_out_20 : std_logic;
signal \n19_adj_735_cascade_\ : std_logic;
signal n13141 : std_logic;
signal n1 : std_logic;
signal n8_adj_747 : std_logic;
signal n9426 : std_logic;
signal n6178 : std_logic;
signal \n7310_cascade_\ : std_logic;
signal \nx.n2398\ : std_logic;
signal \nx.n2397\ : std_logic;
signal neopxl_color_14 : std_logic;
signal neopxl_color_prev_14 : std_logic;
signal \nx.n2400\ : std_logic;
signal \nx.n2400_cascade_\ : std_logic;
signal \nx.n2403\ : std_logic;
signal \nx.n35_adj_658\ : std_logic;
signal \nx.n2402\ : std_logic;
signal \nx.n2406\ : std_logic;
signal \nx.bit_ctr_12\ : std_logic;
signal \nx.n2377\ : std_logic;
signal \bfn_15_23_0_\ : std_logic;
signal \nx.n2309\ : std_logic;
signal \nx.n2376\ : std_logic;
signal \nx.n10708\ : std_logic;
signal \nx.n2308\ : std_logic;
signal \nx.n2375\ : std_logic;
signal \nx.n10709\ : std_logic;
signal \nx.n2307\ : std_logic;
signal \nx.n2374\ : std_logic;
signal \nx.n10710\ : std_logic;
signal \nx.n2306\ : std_logic;
signal \nx.n2373\ : std_logic;
signal \nx.n10711\ : std_logic;
signal \nx.n2305\ : std_logic;
signal \nx.n2372\ : std_logic;
signal \nx.n10712\ : std_logic;
signal \nx.n2304\ : std_logic;
signal \nx.n2371\ : std_logic;
signal \nx.n10713\ : std_logic;
signal \nx.n2303\ : std_logic;
signal \nx.n2370\ : std_logic;
signal \nx.n10714\ : std_logic;
signal \nx.n10715\ : std_logic;
signal \nx.n2302\ : std_logic;
signal \nx.n2369\ : std_logic;
signal \bfn_15_24_0_\ : std_logic;
signal \nx.n2301\ : std_logic;
signal \nx.n2368\ : std_logic;
signal \nx.n10716\ : std_logic;
signal \nx.n2300\ : std_logic;
signal \nx.n2367\ : std_logic;
signal \nx.n10717\ : std_logic;
signal \nx.n2299\ : std_logic;
signal \nx.n2366\ : std_logic;
signal \nx.n10718\ : std_logic;
signal \nx.n2298\ : std_logic;
signal \nx.n2365\ : std_logic;
signal \nx.n10719\ : std_logic;
signal \nx.n2297\ : std_logic;
signal \nx.n2364\ : std_logic;
signal \nx.n10720\ : std_logic;
signal \nx.n2296\ : std_logic;
signal \nx.n2363\ : std_logic;
signal \nx.n10721\ : std_logic;
signal \nx.n2295\ : std_logic;
signal \nx.n2362\ : std_logic;
signal \nx.n10722\ : std_logic;
signal \nx.n10723\ : std_logic;
signal \nx.n2294\ : std_logic;
signal \nx.n2361\ : std_logic;
signal \bfn_15_25_0_\ : std_logic;
signal \nx.n2293\ : std_logic;
signal \nx.n2360\ : std_logic;
signal \nx.n10724\ : std_logic;
signal \nx.n2292\ : std_logic;
signal \nx.n2359\ : std_logic;
signal \nx.n10725\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \nx.n2291\ : std_logic;
signal \nx.n2324\ : std_logic;
signal \nx.n10726\ : std_logic;
signal \nx.n2390\ : std_logic;
signal n26 : std_logic;
signal \bfn_15_26_0_\ : std_logic;
signal n25 : std_logic;
signal n10548 : std_logic;
signal n24 : std_logic;
signal n10549 : std_logic;
signal n23 : std_logic;
signal n10550 : std_logic;
signal n22 : std_logic;
signal n10551 : std_logic;
signal n21_adj_737 : std_logic;
signal n10552 : std_logic;
signal n20 : std_logic;
signal n10553 : std_logic;
signal n19_adj_718 : std_logic;
signal n10554 : std_logic;
signal n10555 : std_logic;
signal n18 : std_logic;
signal \bfn_15_27_0_\ : std_logic;
signal n17 : std_logic;
signal n10556 : std_logic;
signal n16 : std_logic;
signal n10557 : std_logic;
signal n15_adj_759 : std_logic;
signal n10558 : std_logic;
signal n14_adj_745 : std_logic;
signal n10559 : std_logic;
signal n13 : std_logic;
signal n10560 : std_logic;
signal n12 : std_logic;
signal n10561 : std_logic;
signal n11_adj_758 : std_logic;
signal n10562 : std_logic;
signal n10563 : std_logic;
signal n10_adj_757 : std_logic;
signal \bfn_15_28_0_\ : std_logic;
signal n9 : std_logic;
signal n10564 : std_logic;
signal n8_adj_755 : std_logic;
signal n10565 : std_logic;
signal n7 : std_logic;
signal n10566 : std_logic;
signal n6_adj_756 : std_logic;
signal n10567 : std_logic;
signal blink_counter_21 : std_logic;
signal n10568 : std_logic;
signal blink_counter_22 : std_logic;
signal n10569 : std_logic;
signal blink_counter_23 : std_logic;
signal n10570 : std_logic;
signal n10571 : std_logic;
signal blink_counter_24 : std_logic;
signal \bfn_15_29_0_\ : std_logic;
signal n10572 : std_logic;
signal blink_counter_25 : std_logic;
signal n45 : std_logic;
signal \bfn_16_15_0_\ : std_logic;
signal n10510 : std_logic;
signal n10511 : std_logic;
signal n10512 : std_logic;
signal n10513 : std_logic;
signal n10514 : std_logic;
signal n10515 : std_logic;
signal n10516 : std_logic;
signal \n8_adj_763_cascade_\ : std_logic;
signal \current_pin_7__N_155\ : std_logic;
signal n7_adj_719 : std_logic;
signal n21 : std_logic;
signal \current_pin_7__N_155_cascade_\ : std_logic;
signal n7166 : std_logic;
signal n6180 : std_logic;
signal n6971 : std_logic;
signal n12135 : std_logic;
signal n149 : std_logic;
signal n7231 : std_logic;
signal n12208 : std_logic;
signal \n7500_cascade_\ : std_logic;
signal pin_out_22 : std_logic;
signal n8_adj_723 : std_logic;
signal n4_adj_778 : std_logic;
signal n7142 : std_logic;
signal \n7142_cascade_\ : std_logic;
signal counter_7 : std_logic;
signal counter_6 : std_logic;
signal n73 : std_logic;
signal pin_in_7 : std_logic;
signal n2385 : std_logic;
signal \n12123_cascade_\ : std_logic;
signal n48_adj_771 : std_logic;
signal pin_in_4 : std_logic;
signal n2313 : std_logic;
signal \n13144_cascade_\ : std_logic;
signal n13279 : std_logic;
signal n14_adj_717 : std_logic;
signal n11 : std_logic;
signal n30 : std_logic;
signal delay_counter_31 : std_logic;
signal n11612 : std_logic;
signal n11481 : std_logic;
signal n13273 : std_logic;
signal \state_7_N_167_0\ : std_logic;
signal counter_3 : std_logic;
signal counter_4 : std_logic;
signal counter_0 : std_logic;
signal counter_2 : std_logic;
signal counter_1 : std_logic;
signal \n10_adj_762_cascade_\ : std_logic;
signal counter_5 : std_logic;
signal n18_adj_742 : std_logic;
signal n4 : std_logic;
signal pin_out_13 : std_logic;
signal pin_out_12 : std_logic;
signal \n13164_cascade_\ : std_logic;
signal n13468 : std_logic;
signal n6_adj_748 : std_logic;
signal pin_in_22 : std_logic;
signal \n6_adj_748_cascade_\ : std_logic;
signal pin_out_15 : std_logic;
signal pin_out_14 : std_logic;
signal n13165 : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal n10384 : std_logic;
signal n10385 : std_logic;
signal n10386 : std_logic;
signal current_pin_4 : std_logic;
signal n10387 : std_logic;
signal current_pin_5 : std_logic;
signal n10388 : std_logic;
signal current_pin_6 : std_logic;
signal n10389 : std_logic;
signal n10390 : std_logic;
signal current_pin_7 : std_logic;
signal \CLK_c\ : std_logic;
signal n7223 : std_logic;
signal n7401 : std_logic;
signal n7409 : std_logic;
signal n11_adj_743 : std_logic;
signal n2421 : std_logic;
signal n2373 : std_logic;
signal n11_adj_739 : std_logic;
signal n39 : std_logic;
signal n42 : std_logic;
signal \n40_cascade_\ : std_logic;
signal n41 : std_logic;
signal pin_in_19 : std_logic;
signal pin_in_18 : std_logic;
signal pin_in_16 : std_logic;
signal \n13444_cascade_\ : std_logic;
signal pin_in_17 : std_logic;
signal n13447 : std_logic;
signal n14_adj_752 : std_logic;
signal pin_in_5 : std_logic;
signal \n15_adj_749_cascade_\ : std_logic;
signal n15_adj_750 : std_logic;
signal n37 : std_logic;
signal current_pin_0 : std_logic;
signal pin_in_21 : std_logic;
signal pin_in_20 : std_logic;
signal n19_adj_715 : std_logic;
signal n6_adj_766 : std_logic;
signal n54_adj_768 : std_logic;
signal n53_adj_769 : std_logic;
signal \n13037_cascade_\ : std_logic;
signal n55_adj_767 : std_logic;
signal n7249 : std_logic;
signal \n7249_cascade_\ : std_logic;
signal n7395 : std_logic;
signal current_pin_3 : std_logic;
signal n10 : std_logic;
signal current_pin_2 : std_logic;
signal current_pin_1 : std_logic;
signal n9456 : std_logic;
signal state_0 : std_logic;
signal state_1 : std_logic;
signal state_2 : std_logic;
signal n15_adj_721 : std_logic;
signal \_gnd_net_\ : std_logic;

signal \LED_wire\ : std_logic;
signal \NEOPXL_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    LED <= \LED_wire\;
    NEOPXL <= \NEOPXL_wire\;
    \CLK_wire\ <= CLK;

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51103\,
            DIN => \N__51102\,
            DOUT => \N__51101\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51103\,
            PADOUT => \N__51102\,
            PADIN => \N__51101\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__42351\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \NEOPXL_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__51094\,
            DIN => \N__51093\,
            DOUT => \N__51092\,
            PACKAGEPIN => \NEOPXL_wire\
        );

    \NEOPXL_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51094\,
            PADOUT => \N__51093\,
            PADIN => \N__51092\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__18414\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \pin0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__51085\,
            DIN => \N__51084\,
            DOUT => \N__51083\,
            PACKAGEPIN => USBPU
        );

    \pin0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51085\,
            PADOUT => \N__51084\,
            PADIN => \N__51083\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_0,
            DIN1 => OPEN,
            DOUT0 => \N__28623\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35735\
        );

    \pin1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__51076\,
            DIN => \N__51075\,
            DOUT => \N__51074\,
            PACKAGEPIN => ENCODER0_A
        );

    \pin1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51076\,
            PADOUT => \N__51075\,
            PADIN => \N__51074\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_1,
            DIN1 => OPEN,
            DOUT0 => \N__28587\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35801\
        );

    \pin10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__51067\,
            DIN => \N__51066\,
            DOUT => \N__51065\,
            PACKAGEPIN => TX
        );

    \pin10_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51067\,
            PADOUT => \N__51066\,
            PADIN => \N__51065\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_10,
            DIN1 => OPEN,
            DOUT0 => \N__38943\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35670\
        );

    \pin11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__51058\,
            DIN => \N__51057\,
            DOUT => \N__51056\,
            PACKAGEPIN => RX
        );

    \pin11_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51058\,
            PADOUT => \N__51057\,
            PADIN => \N__51056\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_11,
            DIN1 => OPEN,
            DOUT0 => \N__37560\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35734\
        );

    \pin12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__51049\,
            DIN => \N__51048\,
            DOUT => \N__51047\,
            PACKAGEPIN => CS_CLK
        );

    \pin12_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51049\,
            PADOUT => \N__51048\,
            PADIN => \N__51047\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_12,
            DIN1 => OPEN,
            DOUT0 => \N__48045\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35723\
        );

    \pin13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__51040\,
            DIN => \N__51039\,
            DOUT => \N__51038\,
            PACKAGEPIN => CS
        );

    \pin13_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51040\,
            PADOUT => \N__51039\,
            PADIN => \N__51038\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_13,
            DIN1 => OPEN,
            DOUT0 => \N__48084\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35737\
        );

    \pin14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__51031\,
            DIN => \N__51030\,
            DOUT => \N__51029\,
            PACKAGEPIN => CS_MISO
        );

    \pin14_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51031\,
            PADOUT => \N__51030\,
            PADIN => \N__51029\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_14,
            DIN1 => OPEN,
            DOUT0 => \N__47850\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35668\
        );

    \pin15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__51022\,
            DIN => \N__51021\,
            DOUT => \N__51020\,
            PACKAGEPIN => SCL
        );

    \pin15_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51022\,
            PADOUT => \N__51021\,
            PADIN => \N__51020\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_15,
            DIN1 => OPEN,
            DOUT0 => \N__47882\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35768\
        );

    \pin16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__51013\,
            DIN => \N__51012\,
            DOUT => \N__51011\,
            PACKAGEPIN => SDA
        );

    \pin16_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51013\,
            PADOUT => \N__51012\,
            PADIN => \N__51011\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_16,
            DIN1 => OPEN,
            DOUT0 => \N__43101\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35793\
        );

    \pin17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__51004\,
            DIN => \N__51003\,
            DOUT => \N__51002\,
            PACKAGEPIN => INLC
        );

    \pin17_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__51004\,
            PADOUT => \N__51003\,
            PADIN => \N__51002\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_17,
            DIN1 => OPEN,
            DOUT0 => \N__43065\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35796\
        );

    \pin18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50995\,
            DIN => \N__50994\,
            DOUT => \N__50993\,
            PACKAGEPIN => INHC
        );

    \pin18_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50995\,
            PADOUT => \N__50994\,
            PADIN => \N__50993\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_18,
            DIN1 => OPEN,
            DOUT0 => \N__42555\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35795\
        );

    \pin19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50986\,
            DIN => \N__50985\,
            DOUT => \N__50984\,
            PACKAGEPIN => INLB
        );

    \pin19_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50986\,
            PADOUT => \N__50985\,
            PADIN => \N__50984\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_19,
            DIN1 => OPEN,
            DOUT0 => \N__43011\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35772\
        );

    \pin2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50977\,
            DIN => \N__50976\,
            DOUT => \N__50975\,
            PACKAGEPIN => ENCODER0_B
        );

    \pin2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50977\,
            PADOUT => \N__50976\,
            PADIN => \N__50975\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_2,
            DIN1 => OPEN,
            DOUT0 => \N__31374\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35725\
        );

    \pin20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50968\,
            DIN => \N__50967\,
            DOUT => \N__50966\,
            PACKAGEPIN => INHB
        );

    \pin20_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50968\,
            PADOUT => \N__50967\,
            PADIN => \N__50966\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_20,
            DIN1 => OPEN,
            DOUT0 => \N__42867\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35794\
        );

    \pin21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50959\,
            DIN => \N__50958\,
            DOUT => \N__50957\,
            PACKAGEPIN => INLA
        );

    \pin21_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50959\,
            PADOUT => \N__50958\,
            PADIN => \N__50957\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_21,
            DIN1 => OPEN,
            DOUT0 => \N__42909\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35736\
        );

    \pin22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50950\,
            DIN => \N__50949\,
            DOUT => \N__50948\,
            PACKAGEPIN => INHA
        );

    \pin22_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50950\,
            PADOUT => \N__50949\,
            PADIN => \N__50948\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_22,
            DIN1 => OPEN,
            DOUT0 => \N__47337\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35679\
        );

    \pin3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50941\,
            DIN => \N__50940\,
            DOUT => \N__50939\,
            PACKAGEPIN => ENCODER1_A
        );

    \pin3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50941\,
            PADOUT => \N__50940\,
            PADIN => \N__50939\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_3,
            DIN1 => OPEN,
            DOUT0 => \N__31401\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35724\
        );

    \pin4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50932\,
            DIN => \N__50931\,
            DOUT => \N__50930\,
            PACKAGEPIN => ENCODER1_B
        );

    \pin4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50932\,
            PADOUT => \N__50931\,
            PADIN => \N__50930\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_4,
            DIN1 => OPEN,
            DOUT0 => \N__35964\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35733\
        );

    \pin5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50923\,
            DIN => \N__50922\,
            DOUT => \N__50921\,
            PACKAGEPIN => HALL1
        );

    \pin5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50923\,
            PADOUT => \N__50922\,
            PADIN => \N__50921\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_5,
            DIN1 => OPEN,
            DOUT0 => \N__31230\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35800\
        );

    \pin6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50914\,
            DIN => \N__50913\,
            DOUT => \N__50912\,
            PACKAGEPIN => HALL2
        );

    \pin6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50914\,
            PADOUT => \N__50913\,
            PADIN => \N__50912\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_6,
            DIN1 => OPEN,
            DOUT0 => \N__33561\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35782\
        );

    \pin7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50905\,
            DIN => \N__50904\,
            DOUT => \N__50903\,
            PACKAGEPIN => HALL3
        );

    \pin7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50905\,
            PADOUT => \N__50904\,
            PADIN => \N__50903\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_7,
            DIN1 => OPEN,
            DOUT0 => \N__33516\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35783\
        );

    \pin8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50896\,
            DIN => \N__50895\,
            DOUT => \N__50894\,
            PACKAGEPIN => FAULT_N
        );

    \pin8_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50896\,
            PADOUT => \N__50895\,
            PADIN => \N__50894\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_8,
            DIN1 => OPEN,
            DOUT0 => \N__42411\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35802\
        );

    \pin9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__50887\,
            DIN => \N__50886\,
            DOUT => \N__50885\,
            PACKAGEPIN => DE
        );

    \pin9_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50887\,
            PADOUT => \N__50886\,
            PADIN => \N__50885\,
            CLOCKENABLE => 'H',
            DIN0 => pin_in_9,
            DIN1 => OPEN,
            DOUT0 => \N__42507\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__35669\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50878\,
            DIN => \N__50877\,
            DOUT => \N__50876\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__50878\,
            PADOUT => \N__50877\,
            PADIN => \N__50876\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__12374\ : InMux
    port map (
            O => \N__50859\,
            I => \N__50856\
        );

    \I__12373\ : LocalMux
    port map (
            O => \N__50856\,
            I => n6_adj_766
        );

    \I__12372\ : InMux
    port map (
            O => \N__50853\,
            I => \N__50850\
        );

    \I__12371\ : LocalMux
    port map (
            O => \N__50850\,
            I => \N__50847\
        );

    \I__12370\ : Odrv4
    port map (
            O => \N__50847\,
            I => n54_adj_768
        );

    \I__12369\ : InMux
    port map (
            O => \N__50844\,
            I => \N__50841\
        );

    \I__12368\ : LocalMux
    port map (
            O => \N__50841\,
            I => \N__50838\
        );

    \I__12367\ : Span4Mux_h
    port map (
            O => \N__50838\,
            I => \N__50835\
        );

    \I__12366\ : Odrv4
    port map (
            O => \N__50835\,
            I => n53_adj_769
        );

    \I__12365\ : CascadeMux
    port map (
            O => \N__50832\,
            I => \n13037_cascade_\
        );

    \I__12364\ : InMux
    port map (
            O => \N__50829\,
            I => \N__50826\
        );

    \I__12363\ : LocalMux
    port map (
            O => \N__50826\,
            I => \N__50823\
        );

    \I__12362\ : Odrv4
    port map (
            O => \N__50823\,
            I => n55_adj_767
        );

    \I__12361\ : CEMux
    port map (
            O => \N__50820\,
            I => \N__50817\
        );

    \I__12360\ : LocalMux
    port map (
            O => \N__50817\,
            I => \N__50812\
        );

    \I__12359\ : CEMux
    port map (
            O => \N__50816\,
            I => \N__50809\
        );

    \I__12358\ : InMux
    port map (
            O => \N__50815\,
            I => \N__50806\
        );

    \I__12357\ : Span4Mux_h
    port map (
            O => \N__50812\,
            I => \N__50803\
        );

    \I__12356\ : LocalMux
    port map (
            O => \N__50809\,
            I => \N__50800\
        );

    \I__12355\ : LocalMux
    port map (
            O => \N__50806\,
            I => \N__50797\
        );

    \I__12354\ : Odrv4
    port map (
            O => \N__50803\,
            I => n7249
        );

    \I__12353\ : Odrv12
    port map (
            O => \N__50800\,
            I => n7249
        );

    \I__12352\ : Odrv4
    port map (
            O => \N__50797\,
            I => n7249
        );

    \I__12351\ : CascadeMux
    port map (
            O => \N__50790\,
            I => \n7249_cascade_\
        );

    \I__12350\ : SRMux
    port map (
            O => \N__50787\,
            I => \N__50784\
        );

    \I__12349\ : LocalMux
    port map (
            O => \N__50784\,
            I => \N__50781\
        );

    \I__12348\ : Odrv12
    port map (
            O => \N__50781\,
            I => n7395
        );

    \I__12347\ : CascadeMux
    port map (
            O => \N__50778\,
            I => \N__50774\
        );

    \I__12346\ : InMux
    port map (
            O => \N__50777\,
            I => \N__50767\
        );

    \I__12345\ : InMux
    port map (
            O => \N__50774\,
            I => \N__50762\
        );

    \I__12344\ : InMux
    port map (
            O => \N__50773\,
            I => \N__50762\
        );

    \I__12343\ : InMux
    port map (
            O => \N__50772\,
            I => \N__50749\
        );

    \I__12342\ : InMux
    port map (
            O => \N__50771\,
            I => \N__50744\
        );

    \I__12341\ : InMux
    port map (
            O => \N__50770\,
            I => \N__50744\
        );

    \I__12340\ : LocalMux
    port map (
            O => \N__50767\,
            I => \N__50739\
        );

    \I__12339\ : LocalMux
    port map (
            O => \N__50762\,
            I => \N__50739\
        );

    \I__12338\ : InMux
    port map (
            O => \N__50761\,
            I => \N__50734\
        );

    \I__12337\ : InMux
    port map (
            O => \N__50760\,
            I => \N__50734\
        );

    \I__12336\ : InMux
    port map (
            O => \N__50759\,
            I => \N__50731\
        );

    \I__12335\ : InMux
    port map (
            O => \N__50758\,
            I => \N__50727\
        );

    \I__12334\ : CascadeMux
    port map (
            O => \N__50757\,
            I => \N__50723\
        );

    \I__12333\ : InMux
    port map (
            O => \N__50756\,
            I => \N__50718\
        );

    \I__12332\ : InMux
    port map (
            O => \N__50755\,
            I => \N__50715\
        );

    \I__12331\ : CascadeMux
    port map (
            O => \N__50754\,
            I => \N__50709\
        );

    \I__12330\ : InMux
    port map (
            O => \N__50753\,
            I => \N__50706\
        );

    \I__12329\ : InMux
    port map (
            O => \N__50752\,
            I => \N__50703\
        );

    \I__12328\ : LocalMux
    port map (
            O => \N__50749\,
            I => \N__50696\
        );

    \I__12327\ : LocalMux
    port map (
            O => \N__50744\,
            I => \N__50696\
        );

    \I__12326\ : Span4Mux_v
    port map (
            O => \N__50739\,
            I => \N__50696\
        );

    \I__12325\ : LocalMux
    port map (
            O => \N__50734\,
            I => \N__50691\
        );

    \I__12324\ : LocalMux
    port map (
            O => \N__50731\,
            I => \N__50691\
        );

    \I__12323\ : InMux
    port map (
            O => \N__50730\,
            I => \N__50688\
        );

    \I__12322\ : LocalMux
    port map (
            O => \N__50727\,
            I => \N__50684\
        );

    \I__12321\ : InMux
    port map (
            O => \N__50726\,
            I => \N__50675\
        );

    \I__12320\ : InMux
    port map (
            O => \N__50723\,
            I => \N__50675\
        );

    \I__12319\ : InMux
    port map (
            O => \N__50722\,
            I => \N__50675\
        );

    \I__12318\ : InMux
    port map (
            O => \N__50721\,
            I => \N__50675\
        );

    \I__12317\ : LocalMux
    port map (
            O => \N__50718\,
            I => \N__50670\
        );

    \I__12316\ : LocalMux
    port map (
            O => \N__50715\,
            I => \N__50670\
        );

    \I__12315\ : InMux
    port map (
            O => \N__50714\,
            I => \N__50665\
        );

    \I__12314\ : InMux
    port map (
            O => \N__50713\,
            I => \N__50665\
        );

    \I__12313\ : InMux
    port map (
            O => \N__50712\,
            I => \N__50662\
        );

    \I__12312\ : InMux
    port map (
            O => \N__50709\,
            I => \N__50659\
        );

    \I__12311\ : LocalMux
    port map (
            O => \N__50706\,
            I => \N__50656\
        );

    \I__12310\ : LocalMux
    port map (
            O => \N__50703\,
            I => \N__50653\
        );

    \I__12309\ : Span4Mux_h
    port map (
            O => \N__50696\,
            I => \N__50648\
        );

    \I__12308\ : Span4Mux_v
    port map (
            O => \N__50691\,
            I => \N__50648\
        );

    \I__12307\ : LocalMux
    port map (
            O => \N__50688\,
            I => \N__50645\
        );

    \I__12306\ : InMux
    port map (
            O => \N__50687\,
            I => \N__50642\
        );

    \I__12305\ : Span4Mux_v
    port map (
            O => \N__50684\,
            I => \N__50633\
        );

    \I__12304\ : LocalMux
    port map (
            O => \N__50675\,
            I => \N__50633\
        );

    \I__12303\ : Span4Mux_v
    port map (
            O => \N__50670\,
            I => \N__50633\
        );

    \I__12302\ : LocalMux
    port map (
            O => \N__50665\,
            I => \N__50633\
        );

    \I__12301\ : LocalMux
    port map (
            O => \N__50662\,
            I => current_pin_3
        );

    \I__12300\ : LocalMux
    port map (
            O => \N__50659\,
            I => current_pin_3
        );

    \I__12299\ : Odrv4
    port map (
            O => \N__50656\,
            I => current_pin_3
        );

    \I__12298\ : Odrv4
    port map (
            O => \N__50653\,
            I => current_pin_3
        );

    \I__12297\ : Odrv4
    port map (
            O => \N__50648\,
            I => current_pin_3
        );

    \I__12296\ : Odrv12
    port map (
            O => \N__50645\,
            I => current_pin_3
        );

    \I__12295\ : LocalMux
    port map (
            O => \N__50642\,
            I => current_pin_3
        );

    \I__12294\ : Odrv4
    port map (
            O => \N__50633\,
            I => current_pin_3
        );

    \I__12293\ : InMux
    port map (
            O => \N__50616\,
            I => \N__50612\
        );

    \I__12292\ : CascadeMux
    port map (
            O => \N__50615\,
            I => \N__50608\
        );

    \I__12291\ : LocalMux
    port map (
            O => \N__50612\,
            I => \N__50604\
        );

    \I__12290\ : InMux
    port map (
            O => \N__50611\,
            I => \N__50599\
        );

    \I__12289\ : InMux
    port map (
            O => \N__50608\,
            I => \N__50599\
        );

    \I__12288\ : CascadeMux
    port map (
            O => \N__50607\,
            I => \N__50596\
        );

    \I__12287\ : Span4Mux_v
    port map (
            O => \N__50604\,
            I => \N__50590\
        );

    \I__12286\ : LocalMux
    port map (
            O => \N__50599\,
            I => \N__50590\
        );

    \I__12285\ : InMux
    port map (
            O => \N__50596\,
            I => \N__50587\
        );

    \I__12284\ : InMux
    port map (
            O => \N__50595\,
            I => \N__50584\
        );

    \I__12283\ : Span4Mux_h
    port map (
            O => \N__50590\,
            I => \N__50579\
        );

    \I__12282\ : LocalMux
    port map (
            O => \N__50587\,
            I => \N__50579\
        );

    \I__12281\ : LocalMux
    port map (
            O => \N__50584\,
            I => n10
        );

    \I__12280\ : Odrv4
    port map (
            O => \N__50579\,
            I => n10
        );

    \I__12279\ : CascadeMux
    port map (
            O => \N__50574\,
            I => \N__50570\
        );

    \I__12278\ : InMux
    port map (
            O => \N__50573\,
            I => \N__50559\
        );

    \I__12277\ : InMux
    port map (
            O => \N__50570\,
            I => \N__50551\
        );

    \I__12276\ : InMux
    port map (
            O => \N__50569\,
            I => \N__50548\
        );

    \I__12275\ : InMux
    port map (
            O => \N__50568\,
            I => \N__50545\
        );

    \I__12274\ : CascadeMux
    port map (
            O => \N__50567\,
            I => \N__50541\
        );

    \I__12273\ : CascadeMux
    port map (
            O => \N__50566\,
            I => \N__50538\
        );

    \I__12272\ : InMux
    port map (
            O => \N__50565\,
            I => \N__50528\
        );

    \I__12271\ : InMux
    port map (
            O => \N__50564\,
            I => \N__50525\
        );

    \I__12270\ : InMux
    port map (
            O => \N__50563\,
            I => \N__50520\
        );

    \I__12269\ : InMux
    port map (
            O => \N__50562\,
            I => \N__50520\
        );

    \I__12268\ : LocalMux
    port map (
            O => \N__50559\,
            I => \N__50517\
        );

    \I__12267\ : InMux
    port map (
            O => \N__50558\,
            I => \N__50512\
        );

    \I__12266\ : InMux
    port map (
            O => \N__50557\,
            I => \N__50512\
        );

    \I__12265\ : InMux
    port map (
            O => \N__50556\,
            I => \N__50509\
        );

    \I__12264\ : InMux
    port map (
            O => \N__50555\,
            I => \N__50506\
        );

    \I__12263\ : InMux
    port map (
            O => \N__50554\,
            I => \N__50503\
        );

    \I__12262\ : LocalMux
    port map (
            O => \N__50551\,
            I => \N__50500\
        );

    \I__12261\ : LocalMux
    port map (
            O => \N__50548\,
            I => \N__50496\
        );

    \I__12260\ : LocalMux
    port map (
            O => \N__50545\,
            I => \N__50493\
        );

    \I__12259\ : InMux
    port map (
            O => \N__50544\,
            I => \N__50487\
        );

    \I__12258\ : InMux
    port map (
            O => \N__50541\,
            I => \N__50482\
        );

    \I__12257\ : InMux
    port map (
            O => \N__50538\,
            I => \N__50482\
        );

    \I__12256\ : InMux
    port map (
            O => \N__50537\,
            I => \N__50479\
        );

    \I__12255\ : InMux
    port map (
            O => \N__50536\,
            I => \N__50476\
        );

    \I__12254\ : InMux
    port map (
            O => \N__50535\,
            I => \N__50473\
        );

    \I__12253\ : InMux
    port map (
            O => \N__50534\,
            I => \N__50470\
        );

    \I__12252\ : InMux
    port map (
            O => \N__50533\,
            I => \N__50467\
        );

    \I__12251\ : InMux
    port map (
            O => \N__50532\,
            I => \N__50462\
        );

    \I__12250\ : InMux
    port map (
            O => \N__50531\,
            I => \N__50462\
        );

    \I__12249\ : LocalMux
    port map (
            O => \N__50528\,
            I => \N__50459\
        );

    \I__12248\ : LocalMux
    port map (
            O => \N__50525\,
            I => \N__50454\
        );

    \I__12247\ : LocalMux
    port map (
            O => \N__50520\,
            I => \N__50454\
        );

    \I__12246\ : Span4Mux_h
    port map (
            O => \N__50517\,
            I => \N__50449\
        );

    \I__12245\ : LocalMux
    port map (
            O => \N__50512\,
            I => \N__50449\
        );

    \I__12244\ : LocalMux
    port map (
            O => \N__50509\,
            I => \N__50446\
        );

    \I__12243\ : LocalMux
    port map (
            O => \N__50506\,
            I => \N__50437\
        );

    \I__12242\ : LocalMux
    port map (
            O => \N__50503\,
            I => \N__50437\
        );

    \I__12241\ : Span12Mux_v
    port map (
            O => \N__50500\,
            I => \N__50437\
        );

    \I__12240\ : InMux
    port map (
            O => \N__50499\,
            I => \N__50434\
        );

    \I__12239\ : Span4Mux_v
    port map (
            O => \N__50496\,
            I => \N__50429\
        );

    \I__12238\ : Span4Mux_h
    port map (
            O => \N__50493\,
            I => \N__50429\
        );

    \I__12237\ : InMux
    port map (
            O => \N__50492\,
            I => \N__50424\
        );

    \I__12236\ : InMux
    port map (
            O => \N__50491\,
            I => \N__50424\
        );

    \I__12235\ : InMux
    port map (
            O => \N__50490\,
            I => \N__50421\
        );

    \I__12234\ : LocalMux
    port map (
            O => \N__50487\,
            I => \N__50418\
        );

    \I__12233\ : LocalMux
    port map (
            O => \N__50482\,
            I => \N__50411\
        );

    \I__12232\ : LocalMux
    port map (
            O => \N__50479\,
            I => \N__50411\
        );

    \I__12231\ : LocalMux
    port map (
            O => \N__50476\,
            I => \N__50411\
        );

    \I__12230\ : LocalMux
    port map (
            O => \N__50473\,
            I => \N__50398\
        );

    \I__12229\ : LocalMux
    port map (
            O => \N__50470\,
            I => \N__50398\
        );

    \I__12228\ : LocalMux
    port map (
            O => \N__50467\,
            I => \N__50398\
        );

    \I__12227\ : LocalMux
    port map (
            O => \N__50462\,
            I => \N__50398\
        );

    \I__12226\ : Span4Mux_v
    port map (
            O => \N__50459\,
            I => \N__50398\
        );

    \I__12225\ : Span4Mux_h
    port map (
            O => \N__50454\,
            I => \N__50398\
        );

    \I__12224\ : Span4Mux_h
    port map (
            O => \N__50449\,
            I => \N__50393\
        );

    \I__12223\ : Span4Mux_h
    port map (
            O => \N__50446\,
            I => \N__50393\
        );

    \I__12222\ : InMux
    port map (
            O => \N__50445\,
            I => \N__50388\
        );

    \I__12221\ : InMux
    port map (
            O => \N__50444\,
            I => \N__50388\
        );

    \I__12220\ : Span12Mux_h
    port map (
            O => \N__50437\,
            I => \N__50385\
        );

    \I__12219\ : LocalMux
    port map (
            O => \N__50434\,
            I => \N__50378\
        );

    \I__12218\ : Span4Mux_h
    port map (
            O => \N__50429\,
            I => \N__50378\
        );

    \I__12217\ : LocalMux
    port map (
            O => \N__50424\,
            I => \N__50378\
        );

    \I__12216\ : LocalMux
    port map (
            O => \N__50421\,
            I => \N__50369\
        );

    \I__12215\ : Span4Mux_h
    port map (
            O => \N__50418\,
            I => \N__50369\
        );

    \I__12214\ : Span4Mux_v
    port map (
            O => \N__50411\,
            I => \N__50369\
        );

    \I__12213\ : Span4Mux_h
    port map (
            O => \N__50398\,
            I => \N__50369\
        );

    \I__12212\ : Odrv4
    port map (
            O => \N__50393\,
            I => current_pin_2
        );

    \I__12211\ : LocalMux
    port map (
            O => \N__50388\,
            I => current_pin_2
        );

    \I__12210\ : Odrv12
    port map (
            O => \N__50385\,
            I => current_pin_2
        );

    \I__12209\ : Odrv4
    port map (
            O => \N__50378\,
            I => current_pin_2
        );

    \I__12208\ : Odrv4
    port map (
            O => \N__50369\,
            I => current_pin_2
        );

    \I__12207\ : CascadeMux
    port map (
            O => \N__50358\,
            I => \N__50349\
        );

    \I__12206\ : InMux
    port map (
            O => \N__50357\,
            I => \N__50339\
        );

    \I__12205\ : InMux
    port map (
            O => \N__50356\,
            I => \N__50329\
        );

    \I__12204\ : InMux
    port map (
            O => \N__50355\,
            I => \N__50322\
        );

    \I__12203\ : InMux
    port map (
            O => \N__50354\,
            I => \N__50322\
        );

    \I__12202\ : InMux
    port map (
            O => \N__50353\,
            I => \N__50317\
        );

    \I__12201\ : InMux
    port map (
            O => \N__50352\,
            I => \N__50317\
        );

    \I__12200\ : InMux
    port map (
            O => \N__50349\,
            I => \N__50310\
        );

    \I__12199\ : InMux
    port map (
            O => \N__50348\,
            I => \N__50310\
        );

    \I__12198\ : InMux
    port map (
            O => \N__50347\,
            I => \N__50305\
        );

    \I__12197\ : InMux
    port map (
            O => \N__50346\,
            I => \N__50305\
        );

    \I__12196\ : InMux
    port map (
            O => \N__50345\,
            I => \N__50298\
        );

    \I__12195\ : InMux
    port map (
            O => \N__50344\,
            I => \N__50298\
        );

    \I__12194\ : InMux
    port map (
            O => \N__50343\,
            I => \N__50298\
        );

    \I__12193\ : InMux
    port map (
            O => \N__50342\,
            I => \N__50295\
        );

    \I__12192\ : LocalMux
    port map (
            O => \N__50339\,
            I => \N__50292\
        );

    \I__12191\ : CascadeMux
    port map (
            O => \N__50338\,
            I => \N__50289\
        );

    \I__12190\ : InMux
    port map (
            O => \N__50337\,
            I => \N__50281\
        );

    \I__12189\ : InMux
    port map (
            O => \N__50336\,
            I => \N__50272\
        );

    \I__12188\ : InMux
    port map (
            O => \N__50335\,
            I => \N__50272\
        );

    \I__12187\ : InMux
    port map (
            O => \N__50334\,
            I => \N__50272\
        );

    \I__12186\ : InMux
    port map (
            O => \N__50333\,
            I => \N__50272\
        );

    \I__12185\ : CascadeMux
    port map (
            O => \N__50332\,
            I => \N__50269\
        );

    \I__12184\ : LocalMux
    port map (
            O => \N__50329\,
            I => \N__50266\
        );

    \I__12183\ : InMux
    port map (
            O => \N__50328\,
            I => \N__50257\
        );

    \I__12182\ : InMux
    port map (
            O => \N__50327\,
            I => \N__50257\
        );

    \I__12181\ : LocalMux
    port map (
            O => \N__50322\,
            I => \N__50253\
        );

    \I__12180\ : LocalMux
    port map (
            O => \N__50317\,
            I => \N__50250\
        );

    \I__12179\ : InMux
    port map (
            O => \N__50316\,
            I => \N__50247\
        );

    \I__12178\ : InMux
    port map (
            O => \N__50315\,
            I => \N__50244\
        );

    \I__12177\ : LocalMux
    port map (
            O => \N__50310\,
            I => \N__50241\
        );

    \I__12176\ : LocalMux
    port map (
            O => \N__50305\,
            I => \N__50236\
        );

    \I__12175\ : LocalMux
    port map (
            O => \N__50298\,
            I => \N__50236\
        );

    \I__12174\ : LocalMux
    port map (
            O => \N__50295\,
            I => \N__50231\
        );

    \I__12173\ : Span4Mux_h
    port map (
            O => \N__50292\,
            I => \N__50231\
        );

    \I__12172\ : InMux
    port map (
            O => \N__50289\,
            I => \N__50224\
        );

    \I__12171\ : InMux
    port map (
            O => \N__50288\,
            I => \N__50224\
        );

    \I__12170\ : InMux
    port map (
            O => \N__50287\,
            I => \N__50224\
        );

    \I__12169\ : InMux
    port map (
            O => \N__50286\,
            I => \N__50217\
        );

    \I__12168\ : InMux
    port map (
            O => \N__50285\,
            I => \N__50217\
        );

    \I__12167\ : InMux
    port map (
            O => \N__50284\,
            I => \N__50217\
        );

    \I__12166\ : LocalMux
    port map (
            O => \N__50281\,
            I => \N__50212\
        );

    \I__12165\ : LocalMux
    port map (
            O => \N__50272\,
            I => \N__50212\
        );

    \I__12164\ : InMux
    port map (
            O => \N__50269\,
            I => \N__50209\
        );

    \I__12163\ : Span12Mux_v
    port map (
            O => \N__50266\,
            I => \N__50206\
        );

    \I__12162\ : InMux
    port map (
            O => \N__50265\,
            I => \N__50197\
        );

    \I__12161\ : InMux
    port map (
            O => \N__50264\,
            I => \N__50197\
        );

    \I__12160\ : InMux
    port map (
            O => \N__50263\,
            I => \N__50197\
        );

    \I__12159\ : InMux
    port map (
            O => \N__50262\,
            I => \N__50194\
        );

    \I__12158\ : LocalMux
    port map (
            O => \N__50257\,
            I => \N__50191\
        );

    \I__12157\ : InMux
    port map (
            O => \N__50256\,
            I => \N__50188\
        );

    \I__12156\ : Span4Mux_v
    port map (
            O => \N__50253\,
            I => \N__50185\
        );

    \I__12155\ : Span4Mux_h
    port map (
            O => \N__50250\,
            I => \N__50182\
        );

    \I__12154\ : LocalMux
    port map (
            O => \N__50247\,
            I => \N__50173\
        );

    \I__12153\ : LocalMux
    port map (
            O => \N__50244\,
            I => \N__50173\
        );

    \I__12152\ : Span4Mux_h
    port map (
            O => \N__50241\,
            I => \N__50173\
        );

    \I__12151\ : Span4Mux_v
    port map (
            O => \N__50236\,
            I => \N__50173\
        );

    \I__12150\ : Span4Mux_h
    port map (
            O => \N__50231\,
            I => \N__50164\
        );

    \I__12149\ : LocalMux
    port map (
            O => \N__50224\,
            I => \N__50164\
        );

    \I__12148\ : LocalMux
    port map (
            O => \N__50217\,
            I => \N__50164\
        );

    \I__12147\ : Span4Mux_h
    port map (
            O => \N__50212\,
            I => \N__50164\
        );

    \I__12146\ : LocalMux
    port map (
            O => \N__50209\,
            I => \N__50159\
        );

    \I__12145\ : Span12Mux_h
    port map (
            O => \N__50206\,
            I => \N__50159\
        );

    \I__12144\ : InMux
    port map (
            O => \N__50205\,
            I => \N__50154\
        );

    \I__12143\ : InMux
    port map (
            O => \N__50204\,
            I => \N__50154\
        );

    \I__12142\ : LocalMux
    port map (
            O => \N__50197\,
            I => \N__50147\
        );

    \I__12141\ : LocalMux
    port map (
            O => \N__50194\,
            I => \N__50147\
        );

    \I__12140\ : Span12Mux_s11_h
    port map (
            O => \N__50191\,
            I => \N__50147\
        );

    \I__12139\ : LocalMux
    port map (
            O => \N__50188\,
            I => current_pin_1
        );

    \I__12138\ : Odrv4
    port map (
            O => \N__50185\,
            I => current_pin_1
        );

    \I__12137\ : Odrv4
    port map (
            O => \N__50182\,
            I => current_pin_1
        );

    \I__12136\ : Odrv4
    port map (
            O => \N__50173\,
            I => current_pin_1
        );

    \I__12135\ : Odrv4
    port map (
            O => \N__50164\,
            I => current_pin_1
        );

    \I__12134\ : Odrv12
    port map (
            O => \N__50159\,
            I => current_pin_1
        );

    \I__12133\ : LocalMux
    port map (
            O => \N__50154\,
            I => current_pin_1
        );

    \I__12132\ : Odrv12
    port map (
            O => \N__50147\,
            I => current_pin_1
        );

    \I__12131\ : InMux
    port map (
            O => \N__50130\,
            I => \N__50122\
        );

    \I__12130\ : InMux
    port map (
            O => \N__50129\,
            I => \N__50119\
        );

    \I__12129\ : InMux
    port map (
            O => \N__50128\,
            I => \N__50116\
        );

    \I__12128\ : InMux
    port map (
            O => \N__50127\,
            I => \N__50113\
        );

    \I__12127\ : InMux
    port map (
            O => \N__50126\,
            I => \N__50110\
        );

    \I__12126\ : InMux
    port map (
            O => \N__50125\,
            I => \N__50107\
        );

    \I__12125\ : LocalMux
    port map (
            O => \N__50122\,
            I => \N__50104\
        );

    \I__12124\ : LocalMux
    port map (
            O => \N__50119\,
            I => \N__50099\
        );

    \I__12123\ : LocalMux
    port map (
            O => \N__50116\,
            I => \N__50099\
        );

    \I__12122\ : LocalMux
    port map (
            O => \N__50113\,
            I => \N__50094\
        );

    \I__12121\ : LocalMux
    port map (
            O => \N__50110\,
            I => \N__50094\
        );

    \I__12120\ : LocalMux
    port map (
            O => \N__50107\,
            I => \N__50089\
        );

    \I__12119\ : Span4Mux_v
    port map (
            O => \N__50104\,
            I => \N__50089\
        );

    \I__12118\ : Span4Mux_h
    port map (
            O => \N__50099\,
            I => \N__50086\
        );

    \I__12117\ : Odrv12
    port map (
            O => \N__50094\,
            I => n9456
        );

    \I__12116\ : Odrv4
    port map (
            O => \N__50089\,
            I => n9456
        );

    \I__12115\ : Odrv4
    port map (
            O => \N__50086\,
            I => n9456
        );

    \I__12114\ : InMux
    port map (
            O => \N__50079\,
            I => \N__50072\
        );

    \I__12113\ : InMux
    port map (
            O => \N__50078\,
            I => \N__50069\
        );

    \I__12112\ : CascadeMux
    port map (
            O => \N__50077\,
            I => \N__50063\
        );

    \I__12111\ : InMux
    port map (
            O => \N__50076\,
            I => \N__50060\
        );

    \I__12110\ : InMux
    port map (
            O => \N__50075\,
            I => \N__50057\
        );

    \I__12109\ : LocalMux
    port map (
            O => \N__50072\,
            I => \N__50054\
        );

    \I__12108\ : LocalMux
    port map (
            O => \N__50069\,
            I => \N__50051\
        );

    \I__12107\ : InMux
    port map (
            O => \N__50068\,
            I => \N__50048\
        );

    \I__12106\ : InMux
    port map (
            O => \N__50067\,
            I => \N__50045\
        );

    \I__12105\ : CascadeMux
    port map (
            O => \N__50066\,
            I => \N__50041\
        );

    \I__12104\ : InMux
    port map (
            O => \N__50063\,
            I => \N__50038\
        );

    \I__12103\ : LocalMux
    port map (
            O => \N__50060\,
            I => \N__50035\
        );

    \I__12102\ : LocalMux
    port map (
            O => \N__50057\,
            I => \N__50031\
        );

    \I__12101\ : Span4Mux_v
    port map (
            O => \N__50054\,
            I => \N__50028\
        );

    \I__12100\ : Span4Mux_v
    port map (
            O => \N__50051\,
            I => \N__50023\
        );

    \I__12099\ : LocalMux
    port map (
            O => \N__50048\,
            I => \N__50023\
        );

    \I__12098\ : LocalMux
    port map (
            O => \N__50045\,
            I => \N__50020\
        );

    \I__12097\ : InMux
    port map (
            O => \N__50044\,
            I => \N__50017\
        );

    \I__12096\ : InMux
    port map (
            O => \N__50041\,
            I => \N__50011\
        );

    \I__12095\ : LocalMux
    port map (
            O => \N__50038\,
            I => \N__50008\
        );

    \I__12094\ : Span4Mux_v
    port map (
            O => \N__50035\,
            I => \N__50002\
        );

    \I__12093\ : InMux
    port map (
            O => \N__50034\,
            I => \N__49996\
        );

    \I__12092\ : Span4Mux_h
    port map (
            O => \N__50031\,
            I => \N__49993\
        );

    \I__12091\ : Span4Mux_h
    port map (
            O => \N__50028\,
            I => \N__49990\
        );

    \I__12090\ : Span4Mux_h
    port map (
            O => \N__50023\,
            I => \N__49987\
        );

    \I__12089\ : Span4Mux_h
    port map (
            O => \N__50020\,
            I => \N__49979\
        );

    \I__12088\ : LocalMux
    port map (
            O => \N__50017\,
            I => \N__49979\
        );

    \I__12087\ : InMux
    port map (
            O => \N__50016\,
            I => \N__49974\
        );

    \I__12086\ : InMux
    port map (
            O => \N__50015\,
            I => \N__49974\
        );

    \I__12085\ : InMux
    port map (
            O => \N__50014\,
            I => \N__49971\
        );

    \I__12084\ : LocalMux
    port map (
            O => \N__50011\,
            I => \N__49968\
        );

    \I__12083\ : Span4Mux_v
    port map (
            O => \N__50008\,
            I => \N__49965\
        );

    \I__12082\ : InMux
    port map (
            O => \N__50007\,
            I => \N__49962\
        );

    \I__12081\ : InMux
    port map (
            O => \N__50006\,
            I => \N__49957\
        );

    \I__12080\ : InMux
    port map (
            O => \N__50005\,
            I => \N__49957\
        );

    \I__12079\ : Sp12to4
    port map (
            O => \N__50002\,
            I => \N__49951\
        );

    \I__12078\ : InMux
    port map (
            O => \N__50001\,
            I => \N__49948\
        );

    \I__12077\ : InMux
    port map (
            O => \N__50000\,
            I => \N__49943\
        );

    \I__12076\ : InMux
    port map (
            O => \N__49999\,
            I => \N__49943\
        );

    \I__12075\ : LocalMux
    port map (
            O => \N__49996\,
            I => \N__49934\
        );

    \I__12074\ : Span4Mux_v
    port map (
            O => \N__49993\,
            I => \N__49934\
        );

    \I__12073\ : Span4Mux_h
    port map (
            O => \N__49990\,
            I => \N__49934\
        );

    \I__12072\ : Span4Mux_v
    port map (
            O => \N__49987\,
            I => \N__49931\
        );

    \I__12071\ : InMux
    port map (
            O => \N__49986\,
            I => \N__49924\
        );

    \I__12070\ : InMux
    port map (
            O => \N__49985\,
            I => \N__49924\
        );

    \I__12069\ : InMux
    port map (
            O => \N__49984\,
            I => \N__49924\
        );

    \I__12068\ : Span4Mux_h
    port map (
            O => \N__49979\,
            I => \N__49920\
        );

    \I__12067\ : LocalMux
    port map (
            O => \N__49974\,
            I => \N__49915\
        );

    \I__12066\ : LocalMux
    port map (
            O => \N__49971\,
            I => \N__49915\
        );

    \I__12065\ : Span4Mux_v
    port map (
            O => \N__49968\,
            I => \N__49906\
        );

    \I__12064\ : Span4Mux_h
    port map (
            O => \N__49965\,
            I => \N__49906\
        );

    \I__12063\ : LocalMux
    port map (
            O => \N__49962\,
            I => \N__49906\
        );

    \I__12062\ : LocalMux
    port map (
            O => \N__49957\,
            I => \N__49906\
        );

    \I__12061\ : InMux
    port map (
            O => \N__49956\,
            I => \N__49903\
        );

    \I__12060\ : InMux
    port map (
            O => \N__49955\,
            I => \N__49898\
        );

    \I__12059\ : InMux
    port map (
            O => \N__49954\,
            I => \N__49898\
        );

    \I__12058\ : Span12Mux_v
    port map (
            O => \N__49951\,
            I => \N__49893\
        );

    \I__12057\ : LocalMux
    port map (
            O => \N__49948\,
            I => \N__49893\
        );

    \I__12056\ : LocalMux
    port map (
            O => \N__49943\,
            I => \N__49890\
        );

    \I__12055\ : InMux
    port map (
            O => \N__49942\,
            I => \N__49885\
        );

    \I__12054\ : InMux
    port map (
            O => \N__49941\,
            I => \N__49885\
        );

    \I__12053\ : Span4Mux_h
    port map (
            O => \N__49934\,
            I => \N__49878\
        );

    \I__12052\ : Span4Mux_v
    port map (
            O => \N__49931\,
            I => \N__49878\
        );

    \I__12051\ : LocalMux
    port map (
            O => \N__49924\,
            I => \N__49878\
        );

    \I__12050\ : InMux
    port map (
            O => \N__49923\,
            I => \N__49875\
        );

    \I__12049\ : Span4Mux_v
    port map (
            O => \N__49920\,
            I => \N__49868\
        );

    \I__12048\ : Span4Mux_h
    port map (
            O => \N__49915\,
            I => \N__49868\
        );

    \I__12047\ : Span4Mux_h
    port map (
            O => \N__49906\,
            I => \N__49868\
        );

    \I__12046\ : LocalMux
    port map (
            O => \N__49903\,
            I => state_0
        );

    \I__12045\ : LocalMux
    port map (
            O => \N__49898\,
            I => state_0
        );

    \I__12044\ : Odrv12
    port map (
            O => \N__49893\,
            I => state_0
        );

    \I__12043\ : Odrv12
    port map (
            O => \N__49890\,
            I => state_0
        );

    \I__12042\ : LocalMux
    port map (
            O => \N__49885\,
            I => state_0
        );

    \I__12041\ : Odrv4
    port map (
            O => \N__49878\,
            I => state_0
        );

    \I__12040\ : LocalMux
    port map (
            O => \N__49875\,
            I => state_0
        );

    \I__12039\ : Odrv4
    port map (
            O => \N__49868\,
            I => state_0
        );

    \I__12038\ : CascadeMux
    port map (
            O => \N__49851\,
            I => \N__49847\
        );

    \I__12037\ : InMux
    port map (
            O => \N__49850\,
            I => \N__49844\
        );

    \I__12036\ : InMux
    port map (
            O => \N__49847\,
            I => \N__49839\
        );

    \I__12035\ : LocalMux
    port map (
            O => \N__49844\,
            I => \N__49835\
        );

    \I__12034\ : InMux
    port map (
            O => \N__49843\,
            I => \N__49831\
        );

    \I__12033\ : InMux
    port map (
            O => \N__49842\,
            I => \N__49825\
        );

    \I__12032\ : LocalMux
    port map (
            O => \N__49839\,
            I => \N__49822\
        );

    \I__12031\ : InMux
    port map (
            O => \N__49838\,
            I => \N__49819\
        );

    \I__12030\ : Span4Mux_v
    port map (
            O => \N__49835\,
            I => \N__49815\
        );

    \I__12029\ : InMux
    port map (
            O => \N__49834\,
            I => \N__49812\
        );

    \I__12028\ : LocalMux
    port map (
            O => \N__49831\,
            I => \N__49808\
        );

    \I__12027\ : InMux
    port map (
            O => \N__49830\,
            I => \N__49804\
        );

    \I__12026\ : InMux
    port map (
            O => \N__49829\,
            I => \N__49800\
        );

    \I__12025\ : CascadeMux
    port map (
            O => \N__49828\,
            I => \N__49797\
        );

    \I__12024\ : LocalMux
    port map (
            O => \N__49825\,
            I => \N__49793\
        );

    \I__12023\ : Span4Mux_v
    port map (
            O => \N__49822\,
            I => \N__49790\
        );

    \I__12022\ : LocalMux
    port map (
            O => \N__49819\,
            I => \N__49787\
        );

    \I__12021\ : InMux
    port map (
            O => \N__49818\,
            I => \N__49784\
        );

    \I__12020\ : Span4Mux_h
    port map (
            O => \N__49815\,
            I => \N__49779\
        );

    \I__12019\ : LocalMux
    port map (
            O => \N__49812\,
            I => \N__49779\
        );

    \I__12018\ : CascadeMux
    port map (
            O => \N__49811\,
            I => \N__49776\
        );

    \I__12017\ : Span4Mux_h
    port map (
            O => \N__49808\,
            I => \N__49768\
        );

    \I__12016\ : InMux
    port map (
            O => \N__49807\,
            I => \N__49765\
        );

    \I__12015\ : LocalMux
    port map (
            O => \N__49804\,
            I => \N__49762\
        );

    \I__12014\ : InMux
    port map (
            O => \N__49803\,
            I => \N__49759\
        );

    \I__12013\ : LocalMux
    port map (
            O => \N__49800\,
            I => \N__49754\
        );

    \I__12012\ : InMux
    port map (
            O => \N__49797\,
            I => \N__49746\
        );

    \I__12011\ : CascadeMux
    port map (
            O => \N__49796\,
            I => \N__49743\
        );

    \I__12010\ : Span4Mux_v
    port map (
            O => \N__49793\,
            I => \N__49738\
        );

    \I__12009\ : Span4Mux_h
    port map (
            O => \N__49790\,
            I => \N__49738\
        );

    \I__12008\ : Span4Mux_v
    port map (
            O => \N__49787\,
            I => \N__49735\
        );

    \I__12007\ : LocalMux
    port map (
            O => \N__49784\,
            I => \N__49730\
        );

    \I__12006\ : Span4Mux_v
    port map (
            O => \N__49779\,
            I => \N__49730\
        );

    \I__12005\ : InMux
    port map (
            O => \N__49776\,
            I => \N__49723\
        );

    \I__12004\ : InMux
    port map (
            O => \N__49775\,
            I => \N__49723\
        );

    \I__12003\ : InMux
    port map (
            O => \N__49774\,
            I => \N__49723\
        );

    \I__12002\ : InMux
    port map (
            O => \N__49773\,
            I => \N__49719\
        );

    \I__12001\ : CascadeMux
    port map (
            O => \N__49772\,
            I => \N__49716\
        );

    \I__12000\ : InMux
    port map (
            O => \N__49771\,
            I => \N__49713\
        );

    \I__11999\ : Span4Mux_h
    port map (
            O => \N__49768\,
            I => \N__49704\
        );

    \I__11998\ : LocalMux
    port map (
            O => \N__49765\,
            I => \N__49704\
        );

    \I__11997\ : Span4Mux_v
    port map (
            O => \N__49762\,
            I => \N__49704\
        );

    \I__11996\ : LocalMux
    port map (
            O => \N__49759\,
            I => \N__49704\
        );

    \I__11995\ : InMux
    port map (
            O => \N__49758\,
            I => \N__49701\
        );

    \I__11994\ : CascadeMux
    port map (
            O => \N__49757\,
            I => \N__49698\
        );

    \I__11993\ : Sp12to4
    port map (
            O => \N__49754\,
            I => \N__49694\
        );

    \I__11992\ : InMux
    port map (
            O => \N__49753\,
            I => \N__49691\
        );

    \I__11991\ : InMux
    port map (
            O => \N__49752\,
            I => \N__49688\
        );

    \I__11990\ : InMux
    port map (
            O => \N__49751\,
            I => \N__49685\
        );

    \I__11989\ : InMux
    port map (
            O => \N__49750\,
            I => \N__49680\
        );

    \I__11988\ : InMux
    port map (
            O => \N__49749\,
            I => \N__49680\
        );

    \I__11987\ : LocalMux
    port map (
            O => \N__49746\,
            I => \N__49677\
        );

    \I__11986\ : InMux
    port map (
            O => \N__49743\,
            I => \N__49674\
        );

    \I__11985\ : Span4Mux_h
    port map (
            O => \N__49738\,
            I => \N__49665\
        );

    \I__11984\ : Span4Mux_v
    port map (
            O => \N__49735\,
            I => \N__49665\
        );

    \I__11983\ : Span4Mux_v
    port map (
            O => \N__49730\,
            I => \N__49665\
        );

    \I__11982\ : LocalMux
    port map (
            O => \N__49723\,
            I => \N__49665\
        );

    \I__11981\ : InMux
    port map (
            O => \N__49722\,
            I => \N__49662\
        );

    \I__11980\ : LocalMux
    port map (
            O => \N__49719\,
            I => \N__49659\
        );

    \I__11979\ : InMux
    port map (
            O => \N__49716\,
            I => \N__49656\
        );

    \I__11978\ : LocalMux
    port map (
            O => \N__49713\,
            I => \N__49649\
        );

    \I__11977\ : Span4Mux_h
    port map (
            O => \N__49704\,
            I => \N__49649\
        );

    \I__11976\ : LocalMux
    port map (
            O => \N__49701\,
            I => \N__49649\
        );

    \I__11975\ : InMux
    port map (
            O => \N__49698\,
            I => \N__49646\
        );

    \I__11974\ : InMux
    port map (
            O => \N__49697\,
            I => \N__49643\
        );

    \I__11973\ : Span12Mux_v
    port map (
            O => \N__49694\,
            I => \N__49638\
        );

    \I__11972\ : LocalMux
    port map (
            O => \N__49691\,
            I => \N__49638\
        );

    \I__11971\ : LocalMux
    port map (
            O => \N__49688\,
            I => \N__49633\
        );

    \I__11970\ : LocalMux
    port map (
            O => \N__49685\,
            I => \N__49633\
        );

    \I__11969\ : LocalMux
    port map (
            O => \N__49680\,
            I => \N__49620\
        );

    \I__11968\ : Span4Mux_h
    port map (
            O => \N__49677\,
            I => \N__49620\
        );

    \I__11967\ : LocalMux
    port map (
            O => \N__49674\,
            I => \N__49620\
        );

    \I__11966\ : Span4Mux_h
    port map (
            O => \N__49665\,
            I => \N__49620\
        );

    \I__11965\ : LocalMux
    port map (
            O => \N__49662\,
            I => \N__49620\
        );

    \I__11964\ : Span4Mux_v
    port map (
            O => \N__49659\,
            I => \N__49620\
        );

    \I__11963\ : LocalMux
    port map (
            O => \N__49656\,
            I => \N__49615\
        );

    \I__11962\ : Span4Mux_v
    port map (
            O => \N__49649\,
            I => \N__49615\
        );

    \I__11961\ : LocalMux
    port map (
            O => \N__49646\,
            I => state_1
        );

    \I__11960\ : LocalMux
    port map (
            O => \N__49643\,
            I => state_1
        );

    \I__11959\ : Odrv12
    port map (
            O => \N__49638\,
            I => state_1
        );

    \I__11958\ : Odrv4
    port map (
            O => \N__49633\,
            I => state_1
        );

    \I__11957\ : Odrv4
    port map (
            O => \N__49620\,
            I => state_1
        );

    \I__11956\ : Odrv4
    port map (
            O => \N__49615\,
            I => state_1
        );

    \I__11955\ : CascadeMux
    port map (
            O => \N__49602\,
            I => \N__49597\
        );

    \I__11954\ : CascadeMux
    port map (
            O => \N__49601\,
            I => \N__49594\
        );

    \I__11953\ : CascadeMux
    port map (
            O => \N__49600\,
            I => \N__49590\
        );

    \I__11952\ : InMux
    port map (
            O => \N__49597\,
            I => \N__49585\
        );

    \I__11951\ : InMux
    port map (
            O => \N__49594\,
            I => \N__49582\
        );

    \I__11950\ : InMux
    port map (
            O => \N__49593\,
            I => \N__49577\
        );

    \I__11949\ : InMux
    port map (
            O => \N__49590\,
            I => \N__49574\
        );

    \I__11948\ : InMux
    port map (
            O => \N__49589\,
            I => \N__49571\
        );

    \I__11947\ : CascadeMux
    port map (
            O => \N__49588\,
            I => \N__49567\
        );

    \I__11946\ : LocalMux
    port map (
            O => \N__49585\,
            I => \N__49564\
        );

    \I__11945\ : LocalMux
    port map (
            O => \N__49582\,
            I => \N__49561\
        );

    \I__11944\ : InMux
    port map (
            O => \N__49581\,
            I => \N__49558\
        );

    \I__11943\ : InMux
    port map (
            O => \N__49580\,
            I => \N__49555\
        );

    \I__11942\ : LocalMux
    port map (
            O => \N__49577\,
            I => \N__49548\
        );

    \I__11941\ : LocalMux
    port map (
            O => \N__49574\,
            I => \N__49548\
        );

    \I__11940\ : LocalMux
    port map (
            O => \N__49571\,
            I => \N__49545\
        );

    \I__11939\ : InMux
    port map (
            O => \N__49570\,
            I => \N__49542\
        );

    \I__11938\ : InMux
    port map (
            O => \N__49567\,
            I => \N__49539\
        );

    \I__11937\ : Span4Mux_v
    port map (
            O => \N__49564\,
            I => \N__49536\
        );

    \I__11936\ : Span4Mux_v
    port map (
            O => \N__49561\,
            I => \N__49533\
        );

    \I__11935\ : LocalMux
    port map (
            O => \N__49558\,
            I => \N__49528\
        );

    \I__11934\ : LocalMux
    port map (
            O => \N__49555\,
            I => \N__49528\
        );

    \I__11933\ : InMux
    port map (
            O => \N__49554\,
            I => \N__49521\
        );

    \I__11932\ : InMux
    port map (
            O => \N__49553\,
            I => \N__49518\
        );

    \I__11931\ : Span4Mux_v
    port map (
            O => \N__49548\,
            I => \N__49511\
        );

    \I__11930\ : Span4Mux_v
    port map (
            O => \N__49545\,
            I => \N__49511\
        );

    \I__11929\ : LocalMux
    port map (
            O => \N__49542\,
            I => \N__49503\
        );

    \I__11928\ : LocalMux
    port map (
            O => \N__49539\,
            I => \N__49503\
        );

    \I__11927\ : Sp12to4
    port map (
            O => \N__49536\,
            I => \N__49498\
        );

    \I__11926\ : Sp12to4
    port map (
            O => \N__49533\,
            I => \N__49498\
        );

    \I__11925\ : Span4Mux_v
    port map (
            O => \N__49528\,
            I => \N__49495\
        );

    \I__11924\ : InMux
    port map (
            O => \N__49527\,
            I => \N__49490\
        );

    \I__11923\ : InMux
    port map (
            O => \N__49526\,
            I => \N__49490\
        );

    \I__11922\ : InMux
    port map (
            O => \N__49525\,
            I => \N__49484\
        );

    \I__11921\ : InMux
    port map (
            O => \N__49524\,
            I => \N__49484\
        );

    \I__11920\ : LocalMux
    port map (
            O => \N__49521\,
            I => \N__49481\
        );

    \I__11919\ : LocalMux
    port map (
            O => \N__49518\,
            I => \N__49478\
        );

    \I__11918\ : InMux
    port map (
            O => \N__49517\,
            I => \N__49475\
        );

    \I__11917\ : InMux
    port map (
            O => \N__49516\,
            I => \N__49472\
        );

    \I__11916\ : Sp12to4
    port map (
            O => \N__49511\,
            I => \N__49469\
        );

    \I__11915\ : InMux
    port map (
            O => \N__49510\,
            I => \N__49466\
        );

    \I__11914\ : InMux
    port map (
            O => \N__49509\,
            I => \N__49463\
        );

    \I__11913\ : InMux
    port map (
            O => \N__49508\,
            I => \N__49460\
        );

    \I__11912\ : Span12Mux_h
    port map (
            O => \N__49503\,
            I => \N__49455\
        );

    \I__11911\ : Span12Mux_h
    port map (
            O => \N__49498\,
            I => \N__49455\
        );

    \I__11910\ : Span4Mux_h
    port map (
            O => \N__49495\,
            I => \N__49450\
        );

    \I__11909\ : LocalMux
    port map (
            O => \N__49490\,
            I => \N__49450\
        );

    \I__11908\ : InMux
    port map (
            O => \N__49489\,
            I => \N__49447\
        );

    \I__11907\ : LocalMux
    port map (
            O => \N__49484\,
            I => \N__49444\
        );

    \I__11906\ : Span4Mux_v
    port map (
            O => \N__49481\,
            I => \N__49435\
        );

    \I__11905\ : Span4Mux_h
    port map (
            O => \N__49478\,
            I => \N__49435\
        );

    \I__11904\ : LocalMux
    port map (
            O => \N__49475\,
            I => \N__49435\
        );

    \I__11903\ : LocalMux
    port map (
            O => \N__49472\,
            I => \N__49435\
        );

    \I__11902\ : Span12Mux_s11_h
    port map (
            O => \N__49469\,
            I => \N__49426\
        );

    \I__11901\ : LocalMux
    port map (
            O => \N__49466\,
            I => \N__49426\
        );

    \I__11900\ : LocalMux
    port map (
            O => \N__49463\,
            I => \N__49426\
        );

    \I__11899\ : LocalMux
    port map (
            O => \N__49460\,
            I => \N__49426\
        );

    \I__11898\ : Odrv12
    port map (
            O => \N__49455\,
            I => state_2
        );

    \I__11897\ : Odrv4
    port map (
            O => \N__49450\,
            I => state_2
        );

    \I__11896\ : LocalMux
    port map (
            O => \N__49447\,
            I => state_2
        );

    \I__11895\ : Odrv4
    port map (
            O => \N__49444\,
            I => state_2
        );

    \I__11894\ : Odrv4
    port map (
            O => \N__49435\,
            I => state_2
        );

    \I__11893\ : Odrv12
    port map (
            O => \N__49426\,
            I => state_2
        );

    \I__11892\ : CascadeMux
    port map (
            O => \N__49413\,
            I => \N__49407\
        );

    \I__11891\ : InMux
    port map (
            O => \N__49412\,
            I => \N__49403\
        );

    \I__11890\ : InMux
    port map (
            O => \N__49411\,
            I => \N__49396\
        );

    \I__11889\ : InMux
    port map (
            O => \N__49410\,
            I => \N__49396\
        );

    \I__11888\ : InMux
    port map (
            O => \N__49407\,
            I => \N__49396\
        );

    \I__11887\ : InMux
    port map (
            O => \N__49406\,
            I => \N__49393\
        );

    \I__11886\ : LocalMux
    port map (
            O => \N__49403\,
            I => \N__49390\
        );

    \I__11885\ : LocalMux
    port map (
            O => \N__49396\,
            I => \N__49387\
        );

    \I__11884\ : LocalMux
    port map (
            O => \N__49393\,
            I => \N__49384\
        );

    \I__11883\ : Span4Mux_h
    port map (
            O => \N__49390\,
            I => \N__49381\
        );

    \I__11882\ : Span4Mux_h
    port map (
            O => \N__49387\,
            I => \N__49378\
        );

    \I__11881\ : Span4Mux_h
    port map (
            O => \N__49384\,
            I => \N__49375\
        );

    \I__11880\ : Odrv4
    port map (
            O => \N__49381\,
            I => n15_adj_721
        );

    \I__11879\ : Odrv4
    port map (
            O => \N__49378\,
            I => n15_adj_721
        );

    \I__11878\ : Odrv4
    port map (
            O => \N__49375\,
            I => n15_adj_721
        );

    \I__11877\ : InMux
    port map (
            O => \N__49368\,
            I => \N__49365\
        );

    \I__11876\ : LocalMux
    port map (
            O => \N__49365\,
            I => \N__49362\
        );

    \I__11875\ : Odrv4
    port map (
            O => \N__49362\,
            I => n2421
        );

    \I__11874\ : InMux
    port map (
            O => \N__49359\,
            I => \N__49356\
        );

    \I__11873\ : LocalMux
    port map (
            O => \N__49356\,
            I => \N__49353\
        );

    \I__11872\ : Odrv12
    port map (
            O => \N__49353\,
            I => n2373
        );

    \I__11871\ : CascadeMux
    port map (
            O => \N__49350\,
            I => \N__49346\
        );

    \I__11870\ : CascadeMux
    port map (
            O => \N__49349\,
            I => \N__49343\
        );

    \I__11869\ : InMux
    port map (
            O => \N__49346\,
            I => \N__49340\
        );

    \I__11868\ : InMux
    port map (
            O => \N__49343\,
            I => \N__49337\
        );

    \I__11867\ : LocalMux
    port map (
            O => \N__49340\,
            I => \N__49334\
        );

    \I__11866\ : LocalMux
    port map (
            O => \N__49337\,
            I => \N__49331\
        );

    \I__11865\ : Span4Mux_v
    port map (
            O => \N__49334\,
            I => \N__49326\
        );

    \I__11864\ : Span4Mux_h
    port map (
            O => \N__49331\,
            I => \N__49326\
        );

    \I__11863\ : Odrv4
    port map (
            O => \N__49326\,
            I => n11_adj_739
        );

    \I__11862\ : InMux
    port map (
            O => \N__49323\,
            I => \N__49320\
        );

    \I__11861\ : LocalMux
    port map (
            O => \N__49320\,
            I => \N__49317\
        );

    \I__11860\ : Span4Mux_h
    port map (
            O => \N__49317\,
            I => \N__49314\
        );

    \I__11859\ : Odrv4
    port map (
            O => \N__49314\,
            I => n39
        );

    \I__11858\ : InMux
    port map (
            O => \N__49311\,
            I => \N__49308\
        );

    \I__11857\ : LocalMux
    port map (
            O => \N__49308\,
            I => n42
        );

    \I__11856\ : CascadeMux
    port map (
            O => \N__49305\,
            I => \n40_cascade_\
        );

    \I__11855\ : InMux
    port map (
            O => \N__49302\,
            I => \N__49299\
        );

    \I__11854\ : LocalMux
    port map (
            O => \N__49299\,
            I => \N__49296\
        );

    \I__11853\ : Span4Mux_v
    port map (
            O => \N__49296\,
            I => \N__49293\
        );

    \I__11852\ : Odrv4
    port map (
            O => \N__49293\,
            I => n41
        );

    \I__11851\ : InMux
    port map (
            O => \N__49290\,
            I => \N__49287\
        );

    \I__11850\ : LocalMux
    port map (
            O => \N__49287\,
            I => \N__49284\
        );

    \I__11849\ : Span4Mux_v
    port map (
            O => \N__49284\,
            I => \N__49280\
        );

    \I__11848\ : InMux
    port map (
            O => \N__49283\,
            I => \N__49277\
        );

    \I__11847\ : Sp12to4
    port map (
            O => \N__49280\,
            I => \N__49272\
        );

    \I__11846\ : LocalMux
    port map (
            O => \N__49277\,
            I => \N__49272\
        );

    \I__11845\ : Span12Mux_h
    port map (
            O => \N__49272\,
            I => \N__49269\
        );

    \I__11844\ : Span12Mux_v
    port map (
            O => \N__49269\,
            I => \N__49266\
        );

    \I__11843\ : Odrv12
    port map (
            O => \N__49266\,
            I => pin_in_19
        );

    \I__11842\ : InMux
    port map (
            O => \N__49263\,
            I => \N__49260\
        );

    \I__11841\ : LocalMux
    port map (
            O => \N__49260\,
            I => \N__49256\
        );

    \I__11840\ : CascadeMux
    port map (
            O => \N__49259\,
            I => \N__49253\
        );

    \I__11839\ : Span4Mux_v
    port map (
            O => \N__49256\,
            I => \N__49250\
        );

    \I__11838\ : InMux
    port map (
            O => \N__49253\,
            I => \N__49247\
        );

    \I__11837\ : Sp12to4
    port map (
            O => \N__49250\,
            I => \N__49242\
        );

    \I__11836\ : LocalMux
    port map (
            O => \N__49247\,
            I => \N__49242\
        );

    \I__11835\ : Span12Mux_h
    port map (
            O => \N__49242\,
            I => \N__49239\
        );

    \I__11834\ : Span12Mux_v
    port map (
            O => \N__49239\,
            I => \N__49236\
        );

    \I__11833\ : Odrv12
    port map (
            O => \N__49236\,
            I => pin_in_18
        );

    \I__11832\ : CascadeMux
    port map (
            O => \N__49233\,
            I => \N__49230\
        );

    \I__11831\ : InMux
    port map (
            O => \N__49230\,
            I => \N__49227\
        );

    \I__11830\ : LocalMux
    port map (
            O => \N__49227\,
            I => \N__49223\
        );

    \I__11829\ : InMux
    port map (
            O => \N__49226\,
            I => \N__49220\
        );

    \I__11828\ : Span4Mux_h
    port map (
            O => \N__49223\,
            I => \N__49217\
        );

    \I__11827\ : LocalMux
    port map (
            O => \N__49220\,
            I => \N__49214\
        );

    \I__11826\ : Sp12to4
    port map (
            O => \N__49217\,
            I => \N__49211\
        );

    \I__11825\ : Span4Mux_v
    port map (
            O => \N__49214\,
            I => \N__49208\
        );

    \I__11824\ : Span12Mux_v
    port map (
            O => \N__49211\,
            I => \N__49203\
        );

    \I__11823\ : Sp12to4
    port map (
            O => \N__49208\,
            I => \N__49203\
        );

    \I__11822\ : Span12Mux_v
    port map (
            O => \N__49203\,
            I => \N__49200\
        );

    \I__11821\ : Span12Mux_h
    port map (
            O => \N__49200\,
            I => \N__49197\
        );

    \I__11820\ : Odrv12
    port map (
            O => \N__49197\,
            I => pin_in_16
        );

    \I__11819\ : CascadeMux
    port map (
            O => \N__49194\,
            I => \n13444_cascade_\
        );

    \I__11818\ : InMux
    port map (
            O => \N__49191\,
            I => \N__49188\
        );

    \I__11817\ : LocalMux
    port map (
            O => \N__49188\,
            I => \N__49184\
        );

    \I__11816\ : InMux
    port map (
            O => \N__49187\,
            I => \N__49181\
        );

    \I__11815\ : Span4Mux_v
    port map (
            O => \N__49184\,
            I => \N__49178\
        );

    \I__11814\ : LocalMux
    port map (
            O => \N__49181\,
            I => \N__49175\
        );

    \I__11813\ : Span4Mux_h
    port map (
            O => \N__49178\,
            I => \N__49172\
        );

    \I__11812\ : Sp12to4
    port map (
            O => \N__49175\,
            I => \N__49169\
        );

    \I__11811\ : Sp12to4
    port map (
            O => \N__49172\,
            I => \N__49166\
        );

    \I__11810\ : Span12Mux_v
    port map (
            O => \N__49169\,
            I => \N__49163\
        );

    \I__11809\ : Span12Mux_h
    port map (
            O => \N__49166\,
            I => \N__49160\
        );

    \I__11808\ : Span12Mux_h
    port map (
            O => \N__49163\,
            I => \N__49157\
        );

    \I__11807\ : Odrv12
    port map (
            O => \N__49160\,
            I => pin_in_17
        );

    \I__11806\ : Odrv12
    port map (
            O => \N__49157\,
            I => pin_in_17
        );

    \I__11805\ : InMux
    port map (
            O => \N__49152\,
            I => \N__49149\
        );

    \I__11804\ : LocalMux
    port map (
            O => \N__49149\,
            I => n13447
        );

    \I__11803\ : InMux
    port map (
            O => \N__49146\,
            I => \N__49138\
        );

    \I__11802\ : InMux
    port map (
            O => \N__49145\,
            I => \N__49133\
        );

    \I__11801\ : InMux
    port map (
            O => \N__49144\,
            I => \N__49133\
        );

    \I__11800\ : InMux
    port map (
            O => \N__49143\,
            I => \N__49130\
        );

    \I__11799\ : InMux
    port map (
            O => \N__49142\,
            I => \N__49127\
        );

    \I__11798\ : InMux
    port map (
            O => \N__49141\,
            I => \N__49124\
        );

    \I__11797\ : LocalMux
    port map (
            O => \N__49138\,
            I => \N__49120\
        );

    \I__11796\ : LocalMux
    port map (
            O => \N__49133\,
            I => \N__49113\
        );

    \I__11795\ : LocalMux
    port map (
            O => \N__49130\,
            I => \N__49113\
        );

    \I__11794\ : LocalMux
    port map (
            O => \N__49127\,
            I => \N__49113\
        );

    \I__11793\ : LocalMux
    port map (
            O => \N__49124\,
            I => \N__49110\
        );

    \I__11792\ : InMux
    port map (
            O => \N__49123\,
            I => \N__49107\
        );

    \I__11791\ : Span4Mux_v
    port map (
            O => \N__49120\,
            I => \N__49102\
        );

    \I__11790\ : Span4Mux_v
    port map (
            O => \N__49113\,
            I => \N__49102\
        );

    \I__11789\ : Odrv4
    port map (
            O => \N__49110\,
            I => n14_adj_752
        );

    \I__11788\ : LocalMux
    port map (
            O => \N__49107\,
            I => n14_adj_752
        );

    \I__11787\ : Odrv4
    port map (
            O => \N__49102\,
            I => n14_adj_752
        );

    \I__11786\ : InMux
    port map (
            O => \N__49095\,
            I => \N__49092\
        );

    \I__11785\ : LocalMux
    port map (
            O => \N__49092\,
            I => \N__49088\
        );

    \I__11784\ : InMux
    port map (
            O => \N__49091\,
            I => \N__49085\
        );

    \I__11783\ : Sp12to4
    port map (
            O => \N__49088\,
            I => \N__49082\
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__49085\,
            I => \N__49079\
        );

    \I__11781\ : Span12Mux_v
    port map (
            O => \N__49082\,
            I => \N__49076\
        );

    \I__11780\ : Sp12to4
    port map (
            O => \N__49079\,
            I => \N__49073\
        );

    \I__11779\ : Span12Mux_h
    port map (
            O => \N__49076\,
            I => \N__49068\
        );

    \I__11778\ : Span12Mux_v
    port map (
            O => \N__49073\,
            I => \N__49068\
        );

    \I__11777\ : Odrv12
    port map (
            O => \N__49068\,
            I => pin_in_5
        );

    \I__11776\ : CascadeMux
    port map (
            O => \N__49065\,
            I => \n15_adj_749_cascade_\
        );

    \I__11775\ : InMux
    port map (
            O => \N__49062\,
            I => \N__49059\
        );

    \I__11774\ : LocalMux
    port map (
            O => \N__49059\,
            I => n15_adj_750
        );

    \I__11773\ : InMux
    port map (
            O => \N__49056\,
            I => \N__49053\
        );

    \I__11772\ : LocalMux
    port map (
            O => \N__49053\,
            I => n37
        );

    \I__11771\ : CascadeMux
    port map (
            O => \N__49050\,
            I => \N__49045\
        );

    \I__11770\ : CascadeMux
    port map (
            O => \N__49049\,
            I => \N__49037\
        );

    \I__11769\ : CascadeMux
    port map (
            O => \N__49048\,
            I => \N__49034\
        );

    \I__11768\ : InMux
    port map (
            O => \N__49045\,
            I => \N__49021\
        );

    \I__11767\ : InMux
    port map (
            O => \N__49044\,
            I => \N__49021\
        );

    \I__11766\ : InMux
    port map (
            O => \N__49043\,
            I => \N__49021\
        );

    \I__11765\ : InMux
    port map (
            O => \N__49042\,
            I => \N__49021\
        );

    \I__11764\ : InMux
    port map (
            O => \N__49041\,
            I => \N__49018\
        );

    \I__11763\ : CascadeMux
    port map (
            O => \N__49040\,
            I => \N__49011\
        );

    \I__11762\ : InMux
    port map (
            O => \N__49037\,
            I => \N__49008\
        );

    \I__11761\ : InMux
    port map (
            O => \N__49034\,
            I => \N__49005\
        );

    \I__11760\ : InMux
    port map (
            O => \N__49033\,
            I => \N__48989\
        );

    \I__11759\ : InMux
    port map (
            O => \N__49032\,
            I => \N__48986\
        );

    \I__11758\ : InMux
    port map (
            O => \N__49031\,
            I => \N__48979\
        );

    \I__11757\ : InMux
    port map (
            O => \N__49030\,
            I => \N__48979\
        );

    \I__11756\ : LocalMux
    port map (
            O => \N__49021\,
            I => \N__48976\
        );

    \I__11755\ : LocalMux
    port map (
            O => \N__49018\,
            I => \N__48973\
        );

    \I__11754\ : InMux
    port map (
            O => \N__49017\,
            I => \N__48970\
        );

    \I__11753\ : InMux
    port map (
            O => \N__49016\,
            I => \N__48964\
        );

    \I__11752\ : InMux
    port map (
            O => \N__49015\,
            I => \N__48961\
        );

    \I__11751\ : InMux
    port map (
            O => \N__49014\,
            I => \N__48956\
        );

    \I__11750\ : InMux
    port map (
            O => \N__49011\,
            I => \N__48956\
        );

    \I__11749\ : LocalMux
    port map (
            O => \N__49008\,
            I => \N__48950\
        );

    \I__11748\ : LocalMux
    port map (
            O => \N__49005\,
            I => \N__48950\
        );

    \I__11747\ : InMux
    port map (
            O => \N__49004\,
            I => \N__48947\
        );

    \I__11746\ : InMux
    port map (
            O => \N__49003\,
            I => \N__48940\
        );

    \I__11745\ : InMux
    port map (
            O => \N__49002\,
            I => \N__48940\
        );

    \I__11744\ : InMux
    port map (
            O => \N__49001\,
            I => \N__48940\
        );

    \I__11743\ : InMux
    port map (
            O => \N__49000\,
            I => \N__48937\
        );

    \I__11742\ : InMux
    port map (
            O => \N__48999\,
            I => \N__48928\
        );

    \I__11741\ : InMux
    port map (
            O => \N__48998\,
            I => \N__48928\
        );

    \I__11740\ : InMux
    port map (
            O => \N__48997\,
            I => \N__48928\
        );

    \I__11739\ : InMux
    port map (
            O => \N__48996\,
            I => \N__48928\
        );

    \I__11738\ : InMux
    port map (
            O => \N__48995\,
            I => \N__48925\
        );

    \I__11737\ : CascadeMux
    port map (
            O => \N__48994\,
            I => \N__48922\
        );

    \I__11736\ : InMux
    port map (
            O => \N__48993\,
            I => \N__48914\
        );

    \I__11735\ : InMux
    port map (
            O => \N__48992\,
            I => \N__48914\
        );

    \I__11734\ : LocalMux
    port map (
            O => \N__48989\,
            I => \N__48910\
        );

    \I__11733\ : LocalMux
    port map (
            O => \N__48986\,
            I => \N__48907\
        );

    \I__11732\ : InMux
    port map (
            O => \N__48985\,
            I => \N__48902\
        );

    \I__11731\ : InMux
    port map (
            O => \N__48984\,
            I => \N__48902\
        );

    \I__11730\ : LocalMux
    port map (
            O => \N__48979\,
            I => \N__48895\
        );

    \I__11729\ : Span4Mux_v
    port map (
            O => \N__48976\,
            I => \N__48895\
        );

    \I__11728\ : Span4Mux_h
    port map (
            O => \N__48973\,
            I => \N__48895\
        );

    \I__11727\ : LocalMux
    port map (
            O => \N__48970\,
            I => \N__48891\
        );

    \I__11726\ : InMux
    port map (
            O => \N__48969\,
            I => \N__48884\
        );

    \I__11725\ : InMux
    port map (
            O => \N__48968\,
            I => \N__48884\
        );

    \I__11724\ : InMux
    port map (
            O => \N__48967\,
            I => \N__48884\
        );

    \I__11723\ : LocalMux
    port map (
            O => \N__48964\,
            I => \N__48877\
        );

    \I__11722\ : LocalMux
    port map (
            O => \N__48961\,
            I => \N__48877\
        );

    \I__11721\ : LocalMux
    port map (
            O => \N__48956\,
            I => \N__48877\
        );

    \I__11720\ : InMux
    port map (
            O => \N__48955\,
            I => \N__48874\
        );

    \I__11719\ : Span4Mux_v
    port map (
            O => \N__48950\,
            I => \N__48869\
        );

    \I__11718\ : LocalMux
    port map (
            O => \N__48947\,
            I => \N__48869\
        );

    \I__11717\ : LocalMux
    port map (
            O => \N__48940\,
            I => \N__48862\
        );

    \I__11716\ : LocalMux
    port map (
            O => \N__48937\,
            I => \N__48862\
        );

    \I__11715\ : LocalMux
    port map (
            O => \N__48928\,
            I => \N__48862\
        );

    \I__11714\ : LocalMux
    port map (
            O => \N__48925\,
            I => \N__48859\
        );

    \I__11713\ : InMux
    port map (
            O => \N__48922\,
            I => \N__48854\
        );

    \I__11712\ : InMux
    port map (
            O => \N__48921\,
            I => \N__48854\
        );

    \I__11711\ : InMux
    port map (
            O => \N__48920\,
            I => \N__48849\
        );

    \I__11710\ : InMux
    port map (
            O => \N__48919\,
            I => \N__48849\
        );

    \I__11709\ : LocalMux
    port map (
            O => \N__48914\,
            I => \N__48846\
        );

    \I__11708\ : InMux
    port map (
            O => \N__48913\,
            I => \N__48839\
        );

    \I__11707\ : Span4Mux_h
    port map (
            O => \N__48910\,
            I => \N__48836\
        );

    \I__11706\ : Span4Mux_v
    port map (
            O => \N__48907\,
            I => \N__48829\
        );

    \I__11705\ : LocalMux
    port map (
            O => \N__48902\,
            I => \N__48829\
        );

    \I__11704\ : Span4Mux_h
    port map (
            O => \N__48895\,
            I => \N__48829\
        );

    \I__11703\ : InMux
    port map (
            O => \N__48894\,
            I => \N__48826\
        );

    \I__11702\ : Span4Mux_h
    port map (
            O => \N__48891\,
            I => \N__48819\
        );

    \I__11701\ : LocalMux
    port map (
            O => \N__48884\,
            I => \N__48819\
        );

    \I__11700\ : Span4Mux_h
    port map (
            O => \N__48877\,
            I => \N__48819\
        );

    \I__11699\ : LocalMux
    port map (
            O => \N__48874\,
            I => \N__48810\
        );

    \I__11698\ : Span4Mux_h
    port map (
            O => \N__48869\,
            I => \N__48810\
        );

    \I__11697\ : Span4Mux_v
    port map (
            O => \N__48862\,
            I => \N__48810\
        );

    \I__11696\ : Span4Mux_v
    port map (
            O => \N__48859\,
            I => \N__48810\
        );

    \I__11695\ : LocalMux
    port map (
            O => \N__48854\,
            I => \N__48803\
        );

    \I__11694\ : LocalMux
    port map (
            O => \N__48849\,
            I => \N__48803\
        );

    \I__11693\ : Span12Mux_h
    port map (
            O => \N__48846\,
            I => \N__48803\
        );

    \I__11692\ : InMux
    port map (
            O => \N__48845\,
            I => \N__48794\
        );

    \I__11691\ : InMux
    port map (
            O => \N__48844\,
            I => \N__48794\
        );

    \I__11690\ : InMux
    port map (
            O => \N__48843\,
            I => \N__48794\
        );

    \I__11689\ : InMux
    port map (
            O => \N__48842\,
            I => \N__48794\
        );

    \I__11688\ : LocalMux
    port map (
            O => \N__48839\,
            I => \N__48787\
        );

    \I__11687\ : Span4Mux_h
    port map (
            O => \N__48836\,
            I => \N__48787\
        );

    \I__11686\ : Span4Mux_h
    port map (
            O => \N__48829\,
            I => \N__48787\
        );

    \I__11685\ : LocalMux
    port map (
            O => \N__48826\,
            I => current_pin_0
        );

    \I__11684\ : Odrv4
    port map (
            O => \N__48819\,
            I => current_pin_0
        );

    \I__11683\ : Odrv4
    port map (
            O => \N__48810\,
            I => current_pin_0
        );

    \I__11682\ : Odrv12
    port map (
            O => \N__48803\,
            I => current_pin_0
        );

    \I__11681\ : LocalMux
    port map (
            O => \N__48794\,
            I => current_pin_0
        );

    \I__11680\ : Odrv4
    port map (
            O => \N__48787\,
            I => current_pin_0
        );

    \I__11679\ : InMux
    port map (
            O => \N__48774\,
            I => \N__48770\
        );

    \I__11678\ : InMux
    port map (
            O => \N__48773\,
            I => \N__48767\
        );

    \I__11677\ : LocalMux
    port map (
            O => \N__48770\,
            I => \N__48764\
        );

    \I__11676\ : LocalMux
    port map (
            O => \N__48767\,
            I => \N__48761\
        );

    \I__11675\ : Span4Mux_h
    port map (
            O => \N__48764\,
            I => \N__48756\
        );

    \I__11674\ : Span4Mux_h
    port map (
            O => \N__48761\,
            I => \N__48756\
        );

    \I__11673\ : Span4Mux_h
    port map (
            O => \N__48756\,
            I => \N__48753\
        );

    \I__11672\ : Sp12to4
    port map (
            O => \N__48753\,
            I => \N__48750\
        );

    \I__11671\ : Odrv12
    port map (
            O => \N__48750\,
            I => pin_in_21
        );

    \I__11670\ : InMux
    port map (
            O => \N__48747\,
            I => \N__48743\
        );

    \I__11669\ : InMux
    port map (
            O => \N__48746\,
            I => \N__48740\
        );

    \I__11668\ : LocalMux
    port map (
            O => \N__48743\,
            I => \N__48737\
        );

    \I__11667\ : LocalMux
    port map (
            O => \N__48740\,
            I => \N__48734\
        );

    \I__11666\ : Span4Mux_v
    port map (
            O => \N__48737\,
            I => \N__48731\
        );

    \I__11665\ : Span4Mux_v
    port map (
            O => \N__48734\,
            I => \N__48728\
        );

    \I__11664\ : Sp12to4
    port map (
            O => \N__48731\,
            I => \N__48723\
        );

    \I__11663\ : Sp12to4
    port map (
            O => \N__48728\,
            I => \N__48723\
        );

    \I__11662\ : Span12Mux_h
    port map (
            O => \N__48723\,
            I => \N__48720\
        );

    \I__11661\ : Odrv12
    port map (
            O => \N__48720\,
            I => pin_in_20
        );

    \I__11660\ : InMux
    port map (
            O => \N__48717\,
            I => \N__48714\
        );

    \I__11659\ : LocalMux
    port map (
            O => \N__48714\,
            I => n19_adj_715
        );

    \I__11658\ : InMux
    port map (
            O => \N__48711\,
            I => n10384
        );

    \I__11657\ : InMux
    port map (
            O => \N__48708\,
            I => n10385
        );

    \I__11656\ : InMux
    port map (
            O => \N__48705\,
            I => n10386
        );

    \I__11655\ : CascadeMux
    port map (
            O => \N__48702\,
            I => \N__48692\
        );

    \I__11654\ : InMux
    port map (
            O => \N__48701\,
            I => \N__48686\
        );

    \I__11653\ : InMux
    port map (
            O => \N__48700\,
            I => \N__48686\
        );

    \I__11652\ : InMux
    port map (
            O => \N__48699\,
            I => \N__48683\
        );

    \I__11651\ : InMux
    port map (
            O => \N__48698\,
            I => \N__48677\
        );

    \I__11650\ : InMux
    port map (
            O => \N__48697\,
            I => \N__48672\
        );

    \I__11649\ : InMux
    port map (
            O => \N__48696\,
            I => \N__48672\
        );

    \I__11648\ : CascadeMux
    port map (
            O => \N__48695\,
            I => \N__48667\
        );

    \I__11647\ : InMux
    port map (
            O => \N__48692\,
            I => \N__48663\
        );

    \I__11646\ : InMux
    port map (
            O => \N__48691\,
            I => \N__48660\
        );

    \I__11645\ : LocalMux
    port map (
            O => \N__48686\,
            I => \N__48657\
        );

    \I__11644\ : LocalMux
    port map (
            O => \N__48683\,
            I => \N__48654\
        );

    \I__11643\ : InMux
    port map (
            O => \N__48682\,
            I => \N__48651\
        );

    \I__11642\ : InMux
    port map (
            O => \N__48681\,
            I => \N__48648\
        );

    \I__11641\ : InMux
    port map (
            O => \N__48680\,
            I => \N__48642\
        );

    \I__11640\ : LocalMux
    port map (
            O => \N__48677\,
            I => \N__48637\
        );

    \I__11639\ : LocalMux
    port map (
            O => \N__48672\,
            I => \N__48637\
        );

    \I__11638\ : InMux
    port map (
            O => \N__48671\,
            I => \N__48628\
        );

    \I__11637\ : InMux
    port map (
            O => \N__48670\,
            I => \N__48628\
        );

    \I__11636\ : InMux
    port map (
            O => \N__48667\,
            I => \N__48628\
        );

    \I__11635\ : InMux
    port map (
            O => \N__48666\,
            I => \N__48628\
        );

    \I__11634\ : LocalMux
    port map (
            O => \N__48663\,
            I => \N__48625\
        );

    \I__11633\ : LocalMux
    port map (
            O => \N__48660\,
            I => \N__48620\
        );

    \I__11632\ : Span4Mux_h
    port map (
            O => \N__48657\,
            I => \N__48620\
        );

    \I__11631\ : Span4Mux_v
    port map (
            O => \N__48654\,
            I => \N__48613\
        );

    \I__11630\ : LocalMux
    port map (
            O => \N__48651\,
            I => \N__48613\
        );

    \I__11629\ : LocalMux
    port map (
            O => \N__48648\,
            I => \N__48613\
        );

    \I__11628\ : InMux
    port map (
            O => \N__48647\,
            I => \N__48610\
        );

    \I__11627\ : InMux
    port map (
            O => \N__48646\,
            I => \N__48607\
        );

    \I__11626\ : InMux
    port map (
            O => \N__48645\,
            I => \N__48604\
        );

    \I__11625\ : LocalMux
    port map (
            O => \N__48642\,
            I => \N__48597\
        );

    \I__11624\ : Span4Mux_h
    port map (
            O => \N__48637\,
            I => \N__48597\
        );

    \I__11623\ : LocalMux
    port map (
            O => \N__48628\,
            I => \N__48597\
        );

    \I__11622\ : Span4Mux_h
    port map (
            O => \N__48625\,
            I => \N__48594\
        );

    \I__11621\ : Span4Mux_h
    port map (
            O => \N__48620\,
            I => \N__48589\
        );

    \I__11620\ : Span4Mux_h
    port map (
            O => \N__48613\,
            I => \N__48589\
        );

    \I__11619\ : LocalMux
    port map (
            O => \N__48610\,
            I => current_pin_4
        );

    \I__11618\ : LocalMux
    port map (
            O => \N__48607\,
            I => current_pin_4
        );

    \I__11617\ : LocalMux
    port map (
            O => \N__48604\,
            I => current_pin_4
        );

    \I__11616\ : Odrv4
    port map (
            O => \N__48597\,
            I => current_pin_4
        );

    \I__11615\ : Odrv4
    port map (
            O => \N__48594\,
            I => current_pin_4
        );

    \I__11614\ : Odrv4
    port map (
            O => \N__48589\,
            I => current_pin_4
        );

    \I__11613\ : InMux
    port map (
            O => \N__48576\,
            I => n10387
        );

    \I__11612\ : InMux
    port map (
            O => \N__48573\,
            I => \N__48569\
        );

    \I__11611\ : InMux
    port map (
            O => \N__48572\,
            I => \N__48566\
        );

    \I__11610\ : LocalMux
    port map (
            O => \N__48569\,
            I => \N__48563\
        );

    \I__11609\ : LocalMux
    port map (
            O => \N__48566\,
            I => \N__48560\
        );

    \I__11608\ : Span4Mux_v
    port map (
            O => \N__48563\,
            I => \N__48554\
        );

    \I__11607\ : Span4Mux_h
    port map (
            O => \N__48560\,
            I => \N__48554\
        );

    \I__11606\ : InMux
    port map (
            O => \N__48559\,
            I => \N__48550\
        );

    \I__11605\ : Span4Mux_h
    port map (
            O => \N__48554\,
            I => \N__48547\
        );

    \I__11604\ : InMux
    port map (
            O => \N__48553\,
            I => \N__48544\
        );

    \I__11603\ : LocalMux
    port map (
            O => \N__48550\,
            I => current_pin_5
        );

    \I__11602\ : Odrv4
    port map (
            O => \N__48547\,
            I => current_pin_5
        );

    \I__11601\ : LocalMux
    port map (
            O => \N__48544\,
            I => current_pin_5
        );

    \I__11600\ : InMux
    port map (
            O => \N__48537\,
            I => n10388
        );

    \I__11599\ : InMux
    port map (
            O => \N__48534\,
            I => \N__48531\
        );

    \I__11598\ : LocalMux
    port map (
            O => \N__48531\,
            I => \N__48528\
        );

    \I__11597\ : Span4Mux_h
    port map (
            O => \N__48528\,
            I => \N__48523\
        );

    \I__11596\ : InMux
    port map (
            O => \N__48527\,
            I => \N__48520\
        );

    \I__11595\ : InMux
    port map (
            O => \N__48526\,
            I => \N__48516\
        );

    \I__11594\ : Span4Mux_h
    port map (
            O => \N__48523\,
            I => \N__48513\
        );

    \I__11593\ : LocalMux
    port map (
            O => \N__48520\,
            I => \N__48510\
        );

    \I__11592\ : InMux
    port map (
            O => \N__48519\,
            I => \N__48507\
        );

    \I__11591\ : LocalMux
    port map (
            O => \N__48516\,
            I => current_pin_6
        );

    \I__11590\ : Odrv4
    port map (
            O => \N__48513\,
            I => current_pin_6
        );

    \I__11589\ : Odrv12
    port map (
            O => \N__48510\,
            I => current_pin_6
        );

    \I__11588\ : LocalMux
    port map (
            O => \N__48507\,
            I => current_pin_6
        );

    \I__11587\ : InMux
    port map (
            O => \N__48498\,
            I => n10389
        );

    \I__11586\ : InMux
    port map (
            O => \N__48495\,
            I => n10390
        );

    \I__11585\ : CascadeMux
    port map (
            O => \N__48492\,
            I => \N__48489\
        );

    \I__11584\ : InMux
    port map (
            O => \N__48489\,
            I => \N__48486\
        );

    \I__11583\ : LocalMux
    port map (
            O => \N__48486\,
            I => \N__48483\
        );

    \I__11582\ : Span4Mux_h
    port map (
            O => \N__48483\,
            I => \N__48478\
        );

    \I__11581\ : InMux
    port map (
            O => \N__48482\,
            I => \N__48475\
        );

    \I__11580\ : InMux
    port map (
            O => \N__48481\,
            I => \N__48471\
        );

    \I__11579\ : Span4Mux_h
    port map (
            O => \N__48478\,
            I => \N__48468\
        );

    \I__11578\ : LocalMux
    port map (
            O => \N__48475\,
            I => \N__48465\
        );

    \I__11577\ : InMux
    port map (
            O => \N__48474\,
            I => \N__48462\
        );

    \I__11576\ : LocalMux
    port map (
            O => \N__48471\,
            I => current_pin_7
        );

    \I__11575\ : Odrv4
    port map (
            O => \N__48468\,
            I => current_pin_7
        );

    \I__11574\ : Odrv12
    port map (
            O => \N__48465\,
            I => current_pin_7
        );

    \I__11573\ : LocalMux
    port map (
            O => \N__48462\,
            I => current_pin_7
        );

    \I__11572\ : ClkMux
    port map (
            O => \N__48453\,
            I => \N__48240\
        );

    \I__11571\ : ClkMux
    port map (
            O => \N__48452\,
            I => \N__48240\
        );

    \I__11570\ : ClkMux
    port map (
            O => \N__48451\,
            I => \N__48240\
        );

    \I__11569\ : ClkMux
    port map (
            O => \N__48450\,
            I => \N__48240\
        );

    \I__11568\ : ClkMux
    port map (
            O => \N__48449\,
            I => \N__48240\
        );

    \I__11567\ : ClkMux
    port map (
            O => \N__48448\,
            I => \N__48240\
        );

    \I__11566\ : ClkMux
    port map (
            O => \N__48447\,
            I => \N__48240\
        );

    \I__11565\ : ClkMux
    port map (
            O => \N__48446\,
            I => \N__48240\
        );

    \I__11564\ : ClkMux
    port map (
            O => \N__48445\,
            I => \N__48240\
        );

    \I__11563\ : ClkMux
    port map (
            O => \N__48444\,
            I => \N__48240\
        );

    \I__11562\ : ClkMux
    port map (
            O => \N__48443\,
            I => \N__48240\
        );

    \I__11561\ : ClkMux
    port map (
            O => \N__48442\,
            I => \N__48240\
        );

    \I__11560\ : ClkMux
    port map (
            O => \N__48441\,
            I => \N__48240\
        );

    \I__11559\ : ClkMux
    port map (
            O => \N__48440\,
            I => \N__48240\
        );

    \I__11558\ : ClkMux
    port map (
            O => \N__48439\,
            I => \N__48240\
        );

    \I__11557\ : ClkMux
    port map (
            O => \N__48438\,
            I => \N__48240\
        );

    \I__11556\ : ClkMux
    port map (
            O => \N__48437\,
            I => \N__48240\
        );

    \I__11555\ : ClkMux
    port map (
            O => \N__48436\,
            I => \N__48240\
        );

    \I__11554\ : ClkMux
    port map (
            O => \N__48435\,
            I => \N__48240\
        );

    \I__11553\ : ClkMux
    port map (
            O => \N__48434\,
            I => \N__48240\
        );

    \I__11552\ : ClkMux
    port map (
            O => \N__48433\,
            I => \N__48240\
        );

    \I__11551\ : ClkMux
    port map (
            O => \N__48432\,
            I => \N__48240\
        );

    \I__11550\ : ClkMux
    port map (
            O => \N__48431\,
            I => \N__48240\
        );

    \I__11549\ : ClkMux
    port map (
            O => \N__48430\,
            I => \N__48240\
        );

    \I__11548\ : ClkMux
    port map (
            O => \N__48429\,
            I => \N__48240\
        );

    \I__11547\ : ClkMux
    port map (
            O => \N__48428\,
            I => \N__48240\
        );

    \I__11546\ : ClkMux
    port map (
            O => \N__48427\,
            I => \N__48240\
        );

    \I__11545\ : ClkMux
    port map (
            O => \N__48426\,
            I => \N__48240\
        );

    \I__11544\ : ClkMux
    port map (
            O => \N__48425\,
            I => \N__48240\
        );

    \I__11543\ : ClkMux
    port map (
            O => \N__48424\,
            I => \N__48240\
        );

    \I__11542\ : ClkMux
    port map (
            O => \N__48423\,
            I => \N__48240\
        );

    \I__11541\ : ClkMux
    port map (
            O => \N__48422\,
            I => \N__48240\
        );

    \I__11540\ : ClkMux
    port map (
            O => \N__48421\,
            I => \N__48240\
        );

    \I__11539\ : ClkMux
    port map (
            O => \N__48420\,
            I => \N__48240\
        );

    \I__11538\ : ClkMux
    port map (
            O => \N__48419\,
            I => \N__48240\
        );

    \I__11537\ : ClkMux
    port map (
            O => \N__48418\,
            I => \N__48240\
        );

    \I__11536\ : ClkMux
    port map (
            O => \N__48417\,
            I => \N__48240\
        );

    \I__11535\ : ClkMux
    port map (
            O => \N__48416\,
            I => \N__48240\
        );

    \I__11534\ : ClkMux
    port map (
            O => \N__48415\,
            I => \N__48240\
        );

    \I__11533\ : ClkMux
    port map (
            O => \N__48414\,
            I => \N__48240\
        );

    \I__11532\ : ClkMux
    port map (
            O => \N__48413\,
            I => \N__48240\
        );

    \I__11531\ : ClkMux
    port map (
            O => \N__48412\,
            I => \N__48240\
        );

    \I__11530\ : ClkMux
    port map (
            O => \N__48411\,
            I => \N__48240\
        );

    \I__11529\ : ClkMux
    port map (
            O => \N__48410\,
            I => \N__48240\
        );

    \I__11528\ : ClkMux
    port map (
            O => \N__48409\,
            I => \N__48240\
        );

    \I__11527\ : ClkMux
    port map (
            O => \N__48408\,
            I => \N__48240\
        );

    \I__11526\ : ClkMux
    port map (
            O => \N__48407\,
            I => \N__48240\
        );

    \I__11525\ : ClkMux
    port map (
            O => \N__48406\,
            I => \N__48240\
        );

    \I__11524\ : ClkMux
    port map (
            O => \N__48405\,
            I => \N__48240\
        );

    \I__11523\ : ClkMux
    port map (
            O => \N__48404\,
            I => \N__48240\
        );

    \I__11522\ : ClkMux
    port map (
            O => \N__48403\,
            I => \N__48240\
        );

    \I__11521\ : ClkMux
    port map (
            O => \N__48402\,
            I => \N__48240\
        );

    \I__11520\ : ClkMux
    port map (
            O => \N__48401\,
            I => \N__48240\
        );

    \I__11519\ : ClkMux
    port map (
            O => \N__48400\,
            I => \N__48240\
        );

    \I__11518\ : ClkMux
    port map (
            O => \N__48399\,
            I => \N__48240\
        );

    \I__11517\ : ClkMux
    port map (
            O => \N__48398\,
            I => \N__48240\
        );

    \I__11516\ : ClkMux
    port map (
            O => \N__48397\,
            I => \N__48240\
        );

    \I__11515\ : ClkMux
    port map (
            O => \N__48396\,
            I => \N__48240\
        );

    \I__11514\ : ClkMux
    port map (
            O => \N__48395\,
            I => \N__48240\
        );

    \I__11513\ : ClkMux
    port map (
            O => \N__48394\,
            I => \N__48240\
        );

    \I__11512\ : ClkMux
    port map (
            O => \N__48393\,
            I => \N__48240\
        );

    \I__11511\ : ClkMux
    port map (
            O => \N__48392\,
            I => \N__48240\
        );

    \I__11510\ : ClkMux
    port map (
            O => \N__48391\,
            I => \N__48240\
        );

    \I__11509\ : ClkMux
    port map (
            O => \N__48390\,
            I => \N__48240\
        );

    \I__11508\ : ClkMux
    port map (
            O => \N__48389\,
            I => \N__48240\
        );

    \I__11507\ : ClkMux
    port map (
            O => \N__48388\,
            I => \N__48240\
        );

    \I__11506\ : ClkMux
    port map (
            O => \N__48387\,
            I => \N__48240\
        );

    \I__11505\ : ClkMux
    port map (
            O => \N__48386\,
            I => \N__48240\
        );

    \I__11504\ : ClkMux
    port map (
            O => \N__48385\,
            I => \N__48240\
        );

    \I__11503\ : ClkMux
    port map (
            O => \N__48384\,
            I => \N__48240\
        );

    \I__11502\ : ClkMux
    port map (
            O => \N__48383\,
            I => \N__48240\
        );

    \I__11501\ : GlobalMux
    port map (
            O => \N__48240\,
            I => \N__48237\
        );

    \I__11500\ : gio2CtrlBuf
    port map (
            O => \N__48237\,
            I => \CLK_c\
        );

    \I__11499\ : CEMux
    port map (
            O => \N__48234\,
            I => \N__48230\
        );

    \I__11498\ : InMux
    port map (
            O => \N__48233\,
            I => \N__48227\
        );

    \I__11497\ : LocalMux
    port map (
            O => \N__48230\,
            I => n7223
        );

    \I__11496\ : LocalMux
    port map (
            O => \N__48227\,
            I => n7223
        );

    \I__11495\ : SRMux
    port map (
            O => \N__48222\,
            I => \N__48219\
        );

    \I__11494\ : LocalMux
    port map (
            O => \N__48219\,
            I => \N__48216\
        );

    \I__11493\ : Odrv4
    port map (
            O => \N__48216\,
            I => n7401
        );

    \I__11492\ : SRMux
    port map (
            O => \N__48213\,
            I => \N__48210\
        );

    \I__11491\ : LocalMux
    port map (
            O => \N__48210\,
            I => \N__48207\
        );

    \I__11490\ : Sp12to4
    port map (
            O => \N__48207\,
            I => \N__48204\
        );

    \I__11489\ : Odrv12
    port map (
            O => \N__48204\,
            I => n7409
        );

    \I__11488\ : CascadeMux
    port map (
            O => \N__48201\,
            I => \N__48198\
        );

    \I__11487\ : InMux
    port map (
            O => \N__48198\,
            I => \N__48194\
        );

    \I__11486\ : CascadeMux
    port map (
            O => \N__48197\,
            I => \N__48191\
        );

    \I__11485\ : LocalMux
    port map (
            O => \N__48194\,
            I => \N__48188\
        );

    \I__11484\ : InMux
    port map (
            O => \N__48191\,
            I => \N__48185\
        );

    \I__11483\ : Span4Mux_h
    port map (
            O => \N__48188\,
            I => \N__48182\
        );

    \I__11482\ : LocalMux
    port map (
            O => \N__48185\,
            I => n11_adj_743
        );

    \I__11481\ : Odrv4
    port map (
            O => \N__48182\,
            I => n11_adj_743
        );

    \I__11480\ : InMux
    port map (
            O => \N__48177\,
            I => \N__48173\
        );

    \I__11479\ : InMux
    port map (
            O => \N__48176\,
            I => \N__48170\
        );

    \I__11478\ : LocalMux
    port map (
            O => \N__48173\,
            I => counter_1
        );

    \I__11477\ : LocalMux
    port map (
            O => \N__48170\,
            I => counter_1
        );

    \I__11476\ : CascadeMux
    port map (
            O => \N__48165\,
            I => \n10_adj_762_cascade_\
        );

    \I__11475\ : InMux
    port map (
            O => \N__48162\,
            I => \N__48158\
        );

    \I__11474\ : InMux
    port map (
            O => \N__48161\,
            I => \N__48155\
        );

    \I__11473\ : LocalMux
    port map (
            O => \N__48158\,
            I => counter_5
        );

    \I__11472\ : LocalMux
    port map (
            O => \N__48155\,
            I => counter_5
        );

    \I__11471\ : InMux
    port map (
            O => \N__48150\,
            I => \N__48144\
        );

    \I__11470\ : InMux
    port map (
            O => \N__48149\,
            I => \N__48141\
        );

    \I__11469\ : InMux
    port map (
            O => \N__48148\,
            I => \N__48138\
        );

    \I__11468\ : CascadeMux
    port map (
            O => \N__48147\,
            I => \N__48134\
        );

    \I__11467\ : LocalMux
    port map (
            O => \N__48144\,
            I => \N__48129\
        );

    \I__11466\ : LocalMux
    port map (
            O => \N__48141\,
            I => \N__48124\
        );

    \I__11465\ : LocalMux
    port map (
            O => \N__48138\,
            I => \N__48124\
        );

    \I__11464\ : InMux
    port map (
            O => \N__48137\,
            I => \N__48121\
        );

    \I__11463\ : InMux
    port map (
            O => \N__48134\,
            I => \N__48116\
        );

    \I__11462\ : InMux
    port map (
            O => \N__48133\,
            I => \N__48116\
        );

    \I__11461\ : InMux
    port map (
            O => \N__48132\,
            I => \N__48113\
        );

    \I__11460\ : Span4Mux_v
    port map (
            O => \N__48129\,
            I => \N__48108\
        );

    \I__11459\ : Span4Mux_h
    port map (
            O => \N__48124\,
            I => \N__48108\
        );

    \I__11458\ : LocalMux
    port map (
            O => \N__48121\,
            I => \N__48103\
        );

    \I__11457\ : LocalMux
    port map (
            O => \N__48116\,
            I => \N__48103\
        );

    \I__11456\ : LocalMux
    port map (
            O => \N__48113\,
            I => n18_adj_742
        );

    \I__11455\ : Odrv4
    port map (
            O => \N__48108\,
            I => n18_adj_742
        );

    \I__11454\ : Odrv12
    port map (
            O => \N__48103\,
            I => n18_adj_742
        );

    \I__11453\ : InMux
    port map (
            O => \N__48096\,
            I => \N__48093\
        );

    \I__11452\ : LocalMux
    port map (
            O => \N__48093\,
            I => \N__48090\
        );

    \I__11451\ : Span4Mux_v
    port map (
            O => \N__48090\,
            I => \N__48087\
        );

    \I__11450\ : Odrv4
    port map (
            O => \N__48087\,
            I => n4
        );

    \I__11449\ : IoInMux
    port map (
            O => \N__48084\,
            I => \N__48081\
        );

    \I__11448\ : LocalMux
    port map (
            O => \N__48081\,
            I => \N__48078\
        );

    \I__11447\ : IoSpan4Mux
    port map (
            O => \N__48078\,
            I => \N__48074\
        );

    \I__11446\ : InMux
    port map (
            O => \N__48077\,
            I => \N__48070\
        );

    \I__11445\ : Sp12to4
    port map (
            O => \N__48074\,
            I => \N__48067\
        );

    \I__11444\ : CascadeMux
    port map (
            O => \N__48073\,
            I => \N__48064\
        );

    \I__11443\ : LocalMux
    port map (
            O => \N__48070\,
            I => \N__48061\
        );

    \I__11442\ : Span12Mux_s9_h
    port map (
            O => \N__48067\,
            I => \N__48058\
        );

    \I__11441\ : InMux
    port map (
            O => \N__48064\,
            I => \N__48055\
        );

    \I__11440\ : Span4Mux_h
    port map (
            O => \N__48061\,
            I => \N__48052\
        );

    \I__11439\ : Odrv12
    port map (
            O => \N__48058\,
            I => pin_out_13
        );

    \I__11438\ : LocalMux
    port map (
            O => \N__48055\,
            I => pin_out_13
        );

    \I__11437\ : Odrv4
    port map (
            O => \N__48052\,
            I => pin_out_13
        );

    \I__11436\ : IoInMux
    port map (
            O => \N__48045\,
            I => \N__48042\
        );

    \I__11435\ : LocalMux
    port map (
            O => \N__48042\,
            I => \N__48039\
        );

    \I__11434\ : Span12Mux_s5_h
    port map (
            O => \N__48039\,
            I => \N__48035\
        );

    \I__11433\ : InMux
    port map (
            O => \N__48038\,
            I => \N__48032\
        );

    \I__11432\ : Span12Mux_h
    port map (
            O => \N__48035\,
            I => \N__48029\
        );

    \I__11431\ : LocalMux
    port map (
            O => \N__48032\,
            I => \N__48025\
        );

    \I__11430\ : Span12Mux_v
    port map (
            O => \N__48029\,
            I => \N__48022\
        );

    \I__11429\ : InMux
    port map (
            O => \N__48028\,
            I => \N__48019\
        );

    \I__11428\ : Span4Mux_h
    port map (
            O => \N__48025\,
            I => \N__48016\
        );

    \I__11427\ : Odrv12
    port map (
            O => \N__48022\,
            I => pin_out_12
        );

    \I__11426\ : LocalMux
    port map (
            O => \N__48019\,
            I => pin_out_12
        );

    \I__11425\ : Odrv4
    port map (
            O => \N__48016\,
            I => pin_out_12
        );

    \I__11424\ : CascadeMux
    port map (
            O => \N__48009\,
            I => \n13164_cascade_\
        );

    \I__11423\ : InMux
    port map (
            O => \N__48006\,
            I => \N__48003\
        );

    \I__11422\ : LocalMux
    port map (
            O => \N__48003\,
            I => \N__48000\
        );

    \I__11421\ : Odrv4
    port map (
            O => \N__48000\,
            I => n13468
        );

    \I__11420\ : CascadeMux
    port map (
            O => \N__47997\,
            I => \N__47988\
        );

    \I__11419\ : InMux
    port map (
            O => \N__47996\,
            I => \N__47985\
        );

    \I__11418\ : InMux
    port map (
            O => \N__47995\,
            I => \N__47982\
        );

    \I__11417\ : InMux
    port map (
            O => \N__47994\,
            I => \N__47978\
        );

    \I__11416\ : InMux
    port map (
            O => \N__47993\,
            I => \N__47975\
        );

    \I__11415\ : InMux
    port map (
            O => \N__47992\,
            I => \N__47970\
        );

    \I__11414\ : InMux
    port map (
            O => \N__47991\,
            I => \N__47970\
        );

    \I__11413\ : InMux
    port map (
            O => \N__47988\,
            I => \N__47967\
        );

    \I__11412\ : LocalMux
    port map (
            O => \N__47985\,
            I => \N__47964\
        );

    \I__11411\ : LocalMux
    port map (
            O => \N__47982\,
            I => \N__47961\
        );

    \I__11410\ : InMux
    port map (
            O => \N__47981\,
            I => \N__47958\
        );

    \I__11409\ : LocalMux
    port map (
            O => \N__47978\,
            I => \N__47955\
        );

    \I__11408\ : LocalMux
    port map (
            O => \N__47975\,
            I => \N__47950\
        );

    \I__11407\ : LocalMux
    port map (
            O => \N__47970\,
            I => \N__47950\
        );

    \I__11406\ : LocalMux
    port map (
            O => \N__47967\,
            I => \N__47945\
        );

    \I__11405\ : Span4Mux_v
    port map (
            O => \N__47964\,
            I => \N__47945\
        );

    \I__11404\ : Span12Mux_v
    port map (
            O => \N__47961\,
            I => \N__47940\
        );

    \I__11403\ : LocalMux
    port map (
            O => \N__47958\,
            I => \N__47940\
        );

    \I__11402\ : Span4Mux_h
    port map (
            O => \N__47955\,
            I => \N__47935\
        );

    \I__11401\ : Span4Mux_h
    port map (
            O => \N__47950\,
            I => \N__47935\
        );

    \I__11400\ : Odrv4
    port map (
            O => \N__47945\,
            I => n6_adj_748
        );

    \I__11399\ : Odrv12
    port map (
            O => \N__47940\,
            I => n6_adj_748
        );

    \I__11398\ : Odrv4
    port map (
            O => \N__47935\,
            I => n6_adj_748
        );

    \I__11397\ : InMux
    port map (
            O => \N__47928\,
            I => \N__47924\
        );

    \I__11396\ : CascadeMux
    port map (
            O => \N__47927\,
            I => \N__47921\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__47924\,
            I => \N__47918\
        );

    \I__11394\ : InMux
    port map (
            O => \N__47921\,
            I => \N__47915\
        );

    \I__11393\ : Span4Mux_v
    port map (
            O => \N__47918\,
            I => \N__47912\
        );

    \I__11392\ : LocalMux
    port map (
            O => \N__47915\,
            I => \N__47909\
        );

    \I__11391\ : Sp12to4
    port map (
            O => \N__47912\,
            I => \N__47906\
        );

    \I__11390\ : Span4Mux_h
    port map (
            O => \N__47909\,
            I => \N__47903\
        );

    \I__11389\ : Span12Mux_h
    port map (
            O => \N__47906\,
            I => \N__47900\
        );

    \I__11388\ : Span4Mux_h
    port map (
            O => \N__47903\,
            I => \N__47897\
        );

    \I__11387\ : Span12Mux_v
    port map (
            O => \N__47900\,
            I => \N__47894\
        );

    \I__11386\ : Sp12to4
    port map (
            O => \N__47897\,
            I => \N__47891\
        );

    \I__11385\ : Odrv12
    port map (
            O => \N__47894\,
            I => pin_in_22
        );

    \I__11384\ : Odrv12
    port map (
            O => \N__47891\,
            I => pin_in_22
        );

    \I__11383\ : CascadeMux
    port map (
            O => \N__47886\,
            I => \n6_adj_748_cascade_\
        );

    \I__11382\ : InMux
    port map (
            O => \N__47883\,
            I => \N__47879\
        );

    \I__11381\ : IoInMux
    port map (
            O => \N__47882\,
            I => \N__47876\
        );

    \I__11380\ : LocalMux
    port map (
            O => \N__47879\,
            I => \N__47873\
        );

    \I__11379\ : LocalMux
    port map (
            O => \N__47876\,
            I => \N__47870\
        );

    \I__11378\ : Span4Mux_h
    port map (
            O => \N__47873\,
            I => \N__47866\
        );

    \I__11377\ : Span12Mux_s6_h
    port map (
            O => \N__47870\,
            I => \N__47863\
        );

    \I__11376\ : InMux
    port map (
            O => \N__47869\,
            I => \N__47860\
        );

    \I__11375\ : Span4Mux_v
    port map (
            O => \N__47866\,
            I => \N__47857\
        );

    \I__11374\ : Odrv12
    port map (
            O => \N__47863\,
            I => pin_out_15
        );

    \I__11373\ : LocalMux
    port map (
            O => \N__47860\,
            I => pin_out_15
        );

    \I__11372\ : Odrv4
    port map (
            O => \N__47857\,
            I => pin_out_15
        );

    \I__11371\ : IoInMux
    port map (
            O => \N__47850\,
            I => \N__47847\
        );

    \I__11370\ : LocalMux
    port map (
            O => \N__47847\,
            I => \N__47844\
        );

    \I__11369\ : Span12Mux_s5_h
    port map (
            O => \N__47844\,
            I => \N__47840\
        );

    \I__11368\ : InMux
    port map (
            O => \N__47843\,
            I => \N__47836\
        );

    \I__11367\ : Span12Mux_h
    port map (
            O => \N__47840\,
            I => \N__47833\
        );

    \I__11366\ : InMux
    port map (
            O => \N__47839\,
            I => \N__47830\
        );

    \I__11365\ : LocalMux
    port map (
            O => \N__47836\,
            I => \N__47827\
        );

    \I__11364\ : Odrv12
    port map (
            O => \N__47833\,
            I => pin_out_14
        );

    \I__11363\ : LocalMux
    port map (
            O => \N__47830\,
            I => pin_out_14
        );

    \I__11362\ : Odrv4
    port map (
            O => \N__47827\,
            I => pin_out_14
        );

    \I__11361\ : InMux
    port map (
            O => \N__47820\,
            I => \N__47817\
        );

    \I__11360\ : LocalMux
    port map (
            O => \N__47817\,
            I => n13165
        );

    \I__11359\ : InMux
    port map (
            O => \N__47814\,
            I => \bfn_17_17_0_\
        );

    \I__11358\ : CascadeMux
    port map (
            O => \N__47811\,
            I => \n13144_cascade_\
        );

    \I__11357\ : InMux
    port map (
            O => \N__47808\,
            I => \N__47805\
        );

    \I__11356\ : LocalMux
    port map (
            O => \N__47805\,
            I => \N__47802\
        );

    \I__11355\ : Odrv4
    port map (
            O => \N__47802\,
            I => n13279
        );

    \I__11354\ : InMux
    port map (
            O => \N__47799\,
            I => \N__47792\
        );

    \I__11353\ : InMux
    port map (
            O => \N__47798\,
            I => \N__47789\
        );

    \I__11352\ : InMux
    port map (
            O => \N__47797\,
            I => \N__47784\
        );

    \I__11351\ : InMux
    port map (
            O => \N__47796\,
            I => \N__47784\
        );

    \I__11350\ : InMux
    port map (
            O => \N__47795\,
            I => \N__47781\
        );

    \I__11349\ : LocalMux
    port map (
            O => \N__47792\,
            I => \N__47775\
        );

    \I__11348\ : LocalMux
    port map (
            O => \N__47789\,
            I => \N__47770\
        );

    \I__11347\ : LocalMux
    port map (
            O => \N__47784\,
            I => \N__47770\
        );

    \I__11346\ : LocalMux
    port map (
            O => \N__47781\,
            I => \N__47767\
        );

    \I__11345\ : InMux
    port map (
            O => \N__47780\,
            I => \N__47760\
        );

    \I__11344\ : InMux
    port map (
            O => \N__47779\,
            I => \N__47760\
        );

    \I__11343\ : InMux
    port map (
            O => \N__47778\,
            I => \N__47760\
        );

    \I__11342\ : Span4Mux_h
    port map (
            O => \N__47775\,
            I => \N__47757\
        );

    \I__11341\ : Span4Mux_h
    port map (
            O => \N__47770\,
            I => \N__47754\
        );

    \I__11340\ : Span4Mux_h
    port map (
            O => \N__47767\,
            I => \N__47749\
        );

    \I__11339\ : LocalMux
    port map (
            O => \N__47760\,
            I => \N__47749\
        );

    \I__11338\ : Odrv4
    port map (
            O => \N__47757\,
            I => n14_adj_717
        );

    \I__11337\ : Odrv4
    port map (
            O => \N__47754\,
            I => n14_adj_717
        );

    \I__11336\ : Odrv4
    port map (
            O => \N__47749\,
            I => n14_adj_717
        );

    \I__11335\ : InMux
    port map (
            O => \N__47742\,
            I => \N__47738\
        );

    \I__11334\ : InMux
    port map (
            O => \N__47741\,
            I => \N__47735\
        );

    \I__11333\ : LocalMux
    port map (
            O => \N__47738\,
            I => \N__47732\
        );

    \I__11332\ : LocalMux
    port map (
            O => \N__47735\,
            I => n11
        );

    \I__11331\ : Odrv4
    port map (
            O => \N__47732\,
            I => n11
        );

    \I__11330\ : InMux
    port map (
            O => \N__47727\,
            I => \N__47724\
        );

    \I__11329\ : LocalMux
    port map (
            O => \N__47724\,
            I => \N__47721\
        );

    \I__11328\ : Odrv12
    port map (
            O => \N__47721\,
            I => n30
        );

    \I__11327\ : InMux
    port map (
            O => \N__47718\,
            I => \N__47715\
        );

    \I__11326\ : LocalMux
    port map (
            O => \N__47715\,
            I => \N__47712\
        );

    \I__11325\ : Span4Mux_v
    port map (
            O => \N__47712\,
            I => \N__47708\
        );

    \I__11324\ : InMux
    port map (
            O => \N__47711\,
            I => \N__47704\
        );

    \I__11323\ : Span4Mux_v
    port map (
            O => \N__47708\,
            I => \N__47701\
        );

    \I__11322\ : InMux
    port map (
            O => \N__47707\,
            I => \N__47698\
        );

    \I__11321\ : LocalMux
    port map (
            O => \N__47704\,
            I => \N__47695\
        );

    \I__11320\ : Span4Mux_h
    port map (
            O => \N__47701\,
            I => \N__47692\
        );

    \I__11319\ : LocalMux
    port map (
            O => \N__47698\,
            I => delay_counter_31
        );

    \I__11318\ : Odrv12
    port map (
            O => \N__47695\,
            I => delay_counter_31
        );

    \I__11317\ : Odrv4
    port map (
            O => \N__47692\,
            I => delay_counter_31
        );

    \I__11316\ : InMux
    port map (
            O => \N__47685\,
            I => \N__47682\
        );

    \I__11315\ : LocalMux
    port map (
            O => \N__47682\,
            I => \N__47679\
        );

    \I__11314\ : Span4Mux_v
    port map (
            O => \N__47679\,
            I => \N__47675\
        );

    \I__11313\ : InMux
    port map (
            O => \N__47678\,
            I => \N__47672\
        );

    \I__11312\ : Span4Mux_h
    port map (
            O => \N__47675\,
            I => \N__47669\
        );

    \I__11311\ : LocalMux
    port map (
            O => \N__47672\,
            I => n11612
        );

    \I__11310\ : Odrv4
    port map (
            O => \N__47669\,
            I => n11612
        );

    \I__11309\ : CascadeMux
    port map (
            O => \N__47664\,
            I => \N__47661\
        );

    \I__11308\ : InMux
    port map (
            O => \N__47661\,
            I => \N__47658\
        );

    \I__11307\ : LocalMux
    port map (
            O => \N__47658\,
            I => \N__47655\
        );

    \I__11306\ : Span12Mux_h
    port map (
            O => \N__47655\,
            I => \N__47651\
        );

    \I__11305\ : InMux
    port map (
            O => \N__47654\,
            I => \N__47648\
        );

    \I__11304\ : Odrv12
    port map (
            O => \N__47651\,
            I => n11481
        );

    \I__11303\ : LocalMux
    port map (
            O => \N__47648\,
            I => n11481
        );

    \I__11302\ : InMux
    port map (
            O => \N__47643\,
            I => \N__47640\
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__47640\,
            I => \N__47637\
        );

    \I__11300\ : Span4Mux_v
    port map (
            O => \N__47637\,
            I => \N__47634\
        );

    \I__11299\ : Odrv4
    port map (
            O => \N__47634\,
            I => n13273
        );

    \I__11298\ : InMux
    port map (
            O => \N__47631\,
            I => \N__47627\
        );

    \I__11297\ : CascadeMux
    port map (
            O => \N__47630\,
            I => \N__47624\
        );

    \I__11296\ : LocalMux
    port map (
            O => \N__47627\,
            I => \N__47621\
        );

    \I__11295\ : InMux
    port map (
            O => \N__47624\,
            I => \N__47618\
        );

    \I__11294\ : Span4Mux_v
    port map (
            O => \N__47621\,
            I => \N__47612\
        );

    \I__11293\ : LocalMux
    port map (
            O => \N__47618\,
            I => \N__47612\
        );

    \I__11292\ : InMux
    port map (
            O => \N__47617\,
            I => \N__47609\
        );

    \I__11291\ : Span4Mux_v
    port map (
            O => \N__47612\,
            I => \N__47604\
        );

    \I__11290\ : LocalMux
    port map (
            O => \N__47609\,
            I => \N__47604\
        );

    \I__11289\ : Span4Mux_h
    port map (
            O => \N__47604\,
            I => \N__47601\
        );

    \I__11288\ : Odrv4
    port map (
            O => \N__47601\,
            I => \state_7_N_167_0\
        );

    \I__11287\ : InMux
    port map (
            O => \N__47598\,
            I => \N__47594\
        );

    \I__11286\ : InMux
    port map (
            O => \N__47597\,
            I => \N__47591\
        );

    \I__11285\ : LocalMux
    port map (
            O => \N__47594\,
            I => counter_3
        );

    \I__11284\ : LocalMux
    port map (
            O => \N__47591\,
            I => counter_3
        );

    \I__11283\ : CascadeMux
    port map (
            O => \N__47586\,
            I => \N__47583\
        );

    \I__11282\ : InMux
    port map (
            O => \N__47583\,
            I => \N__47579\
        );

    \I__11281\ : InMux
    port map (
            O => \N__47582\,
            I => \N__47576\
        );

    \I__11280\ : LocalMux
    port map (
            O => \N__47579\,
            I => counter_4
        );

    \I__11279\ : LocalMux
    port map (
            O => \N__47576\,
            I => counter_4
        );

    \I__11278\ : CascadeMux
    port map (
            O => \N__47571\,
            I => \N__47567\
        );

    \I__11277\ : InMux
    port map (
            O => \N__47570\,
            I => \N__47564\
        );

    \I__11276\ : InMux
    port map (
            O => \N__47567\,
            I => \N__47561\
        );

    \I__11275\ : LocalMux
    port map (
            O => \N__47564\,
            I => counter_0
        );

    \I__11274\ : LocalMux
    port map (
            O => \N__47561\,
            I => counter_0
        );

    \I__11273\ : CascadeMux
    port map (
            O => \N__47556\,
            I => \N__47553\
        );

    \I__11272\ : InMux
    port map (
            O => \N__47553\,
            I => \N__47550\
        );

    \I__11271\ : LocalMux
    port map (
            O => \N__47550\,
            I => \N__47546\
        );

    \I__11270\ : InMux
    port map (
            O => \N__47549\,
            I => \N__47543\
        );

    \I__11269\ : Odrv4
    port map (
            O => \N__47546\,
            I => counter_2
        );

    \I__11268\ : LocalMux
    port map (
            O => \N__47543\,
            I => counter_2
        );

    \I__11267\ : CEMux
    port map (
            O => \N__47538\,
            I => \N__47535\
        );

    \I__11266\ : LocalMux
    port map (
            O => \N__47535\,
            I => \N__47531\
        );

    \I__11265\ : CascadeMux
    port map (
            O => \N__47534\,
            I => \N__47520\
        );

    \I__11264\ : Span4Mux_v
    port map (
            O => \N__47531\,
            I => \N__47515\
        );

    \I__11263\ : CEMux
    port map (
            O => \N__47530\,
            I => \N__47512\
        );

    \I__11262\ : InMux
    port map (
            O => \N__47529\,
            I => \N__47507\
        );

    \I__11261\ : InMux
    port map (
            O => \N__47528\,
            I => \N__47507\
        );

    \I__11260\ : CascadeMux
    port map (
            O => \N__47527\,
            I => \N__47498\
        );

    \I__11259\ : InMux
    port map (
            O => \N__47526\,
            I => \N__47490\
        );

    \I__11258\ : InMux
    port map (
            O => \N__47525\,
            I => \N__47487\
        );

    \I__11257\ : InMux
    port map (
            O => \N__47524\,
            I => \N__47484\
        );

    \I__11256\ : InMux
    port map (
            O => \N__47523\,
            I => \N__47477\
        );

    \I__11255\ : InMux
    port map (
            O => \N__47520\,
            I => \N__47477\
        );

    \I__11254\ : InMux
    port map (
            O => \N__47519\,
            I => \N__47477\
        );

    \I__11253\ : InMux
    port map (
            O => \N__47518\,
            I => \N__47473\
        );

    \I__11252\ : Span4Mux_v
    port map (
            O => \N__47515\,
            I => \N__47468\
        );

    \I__11251\ : LocalMux
    port map (
            O => \N__47512\,
            I => \N__47468\
        );

    \I__11250\ : LocalMux
    port map (
            O => \N__47507\,
            I => \N__47465\
        );

    \I__11249\ : InMux
    port map (
            O => \N__47506\,
            I => \N__47462\
        );

    \I__11248\ : InMux
    port map (
            O => \N__47505\,
            I => \N__47459\
        );

    \I__11247\ : InMux
    port map (
            O => \N__47504\,
            I => \N__47455\
        );

    \I__11246\ : InMux
    port map (
            O => \N__47503\,
            I => \N__47448\
        );

    \I__11245\ : InMux
    port map (
            O => \N__47502\,
            I => \N__47448\
        );

    \I__11244\ : InMux
    port map (
            O => \N__47501\,
            I => \N__47448\
        );

    \I__11243\ : InMux
    port map (
            O => \N__47498\,
            I => \N__47445\
        );

    \I__11242\ : InMux
    port map (
            O => \N__47497\,
            I => \N__47442\
        );

    \I__11241\ : InMux
    port map (
            O => \N__47496\,
            I => \N__47437\
        );

    \I__11240\ : InMux
    port map (
            O => \N__47495\,
            I => \N__47437\
        );

    \I__11239\ : InMux
    port map (
            O => \N__47494\,
            I => \N__47432\
        );

    \I__11238\ : InMux
    port map (
            O => \N__47493\,
            I => \N__47432\
        );

    \I__11237\ : LocalMux
    port map (
            O => \N__47490\,
            I => \N__47423\
        );

    \I__11236\ : LocalMux
    port map (
            O => \N__47487\,
            I => \N__47423\
        );

    \I__11235\ : LocalMux
    port map (
            O => \N__47484\,
            I => \N__47423\
        );

    \I__11234\ : LocalMux
    port map (
            O => \N__47477\,
            I => \N__47423\
        );

    \I__11233\ : InMux
    port map (
            O => \N__47476\,
            I => \N__47419\
        );

    \I__11232\ : LocalMux
    port map (
            O => \N__47473\,
            I => \N__47416\
        );

    \I__11231\ : Span4Mux_v
    port map (
            O => \N__47468\,
            I => \N__47409\
        );

    \I__11230\ : Span4Mux_h
    port map (
            O => \N__47465\,
            I => \N__47409\
        );

    \I__11229\ : LocalMux
    port map (
            O => \N__47462\,
            I => \N__47409\
        );

    \I__11228\ : LocalMux
    port map (
            O => \N__47459\,
            I => \N__47406\
        );

    \I__11227\ : InMux
    port map (
            O => \N__47458\,
            I => \N__47403\
        );

    \I__11226\ : LocalMux
    port map (
            O => \N__47455\,
            I => \N__47398\
        );

    \I__11225\ : LocalMux
    port map (
            O => \N__47448\,
            I => \N__47398\
        );

    \I__11224\ : LocalMux
    port map (
            O => \N__47445\,
            I => \N__47395\
        );

    \I__11223\ : LocalMux
    port map (
            O => \N__47442\,
            I => \N__47390\
        );

    \I__11222\ : LocalMux
    port map (
            O => \N__47437\,
            I => \N__47390\
        );

    \I__11221\ : LocalMux
    port map (
            O => \N__47432\,
            I => \N__47385\
        );

    \I__11220\ : Span4Mux_v
    port map (
            O => \N__47423\,
            I => \N__47385\
        );

    \I__11219\ : InMux
    port map (
            O => \N__47422\,
            I => \N__47382\
        );

    \I__11218\ : LocalMux
    port map (
            O => \N__47419\,
            I => \N__47379\
        );

    \I__11217\ : Span4Mux_h
    port map (
            O => \N__47416\,
            I => \N__47374\
        );

    \I__11216\ : Span4Mux_h
    port map (
            O => \N__47409\,
            I => \N__47374\
        );

    \I__11215\ : Span4Mux_v
    port map (
            O => \N__47406\,
            I => \N__47369\
        );

    \I__11214\ : LocalMux
    port map (
            O => \N__47403\,
            I => \N__47369\
        );

    \I__11213\ : Span4Mux_v
    port map (
            O => \N__47398\,
            I => \N__47366\
        );

    \I__11212\ : Span4Mux_v
    port map (
            O => \N__47395\,
            I => \N__47359\
        );

    \I__11211\ : Span4Mux_v
    port map (
            O => \N__47390\,
            I => \N__47359\
        );

    \I__11210\ : Span4Mux_h
    port map (
            O => \N__47385\,
            I => \N__47359\
        );

    \I__11209\ : LocalMux
    port map (
            O => \N__47382\,
            I => n7231
        );

    \I__11208\ : Odrv4
    port map (
            O => \N__47379\,
            I => n7231
        );

    \I__11207\ : Odrv4
    port map (
            O => \N__47374\,
            I => n7231
        );

    \I__11206\ : Odrv4
    port map (
            O => \N__47369\,
            I => n7231
        );

    \I__11205\ : Odrv4
    port map (
            O => \N__47366\,
            I => n7231
        );

    \I__11204\ : Odrv4
    port map (
            O => \N__47359\,
            I => n7231
        );

    \I__11203\ : InMux
    port map (
            O => \N__47346\,
            I => \N__47343\
        );

    \I__11202\ : LocalMux
    port map (
            O => \N__47343\,
            I => n12208
        );

    \I__11201\ : CascadeMux
    port map (
            O => \N__47340\,
            I => \n7500_cascade_\
        );

    \I__11200\ : IoInMux
    port map (
            O => \N__47337\,
            I => \N__47334\
        );

    \I__11199\ : LocalMux
    port map (
            O => \N__47334\,
            I => \N__47331\
        );

    \I__11198\ : Span4Mux_s3_v
    port map (
            O => \N__47331\,
            I => \N__47328\
        );

    \I__11197\ : Sp12to4
    port map (
            O => \N__47328\,
            I => \N__47325\
        );

    \I__11196\ : Span12Mux_h
    port map (
            O => \N__47325\,
            I => \N__47320\
        );

    \I__11195\ : CascadeMux
    port map (
            O => \N__47324\,
            I => \N__47317\
        );

    \I__11194\ : InMux
    port map (
            O => \N__47323\,
            I => \N__47314\
        );

    \I__11193\ : Span12Mux_v
    port map (
            O => \N__47320\,
            I => \N__47311\
        );

    \I__11192\ : InMux
    port map (
            O => \N__47317\,
            I => \N__47308\
        );

    \I__11191\ : LocalMux
    port map (
            O => \N__47314\,
            I => \N__47305\
        );

    \I__11190\ : Odrv12
    port map (
            O => \N__47311\,
            I => pin_out_22
        );

    \I__11189\ : LocalMux
    port map (
            O => \N__47308\,
            I => pin_out_22
        );

    \I__11188\ : Odrv4
    port map (
            O => \N__47305\,
            I => pin_out_22
        );

    \I__11187\ : InMux
    port map (
            O => \N__47298\,
            I => \N__47295\
        );

    \I__11186\ : LocalMux
    port map (
            O => \N__47295\,
            I => \N__47291\
        );

    \I__11185\ : InMux
    port map (
            O => \N__47294\,
            I => \N__47287\
        );

    \I__11184\ : Span4Mux_v
    port map (
            O => \N__47291\,
            I => \N__47284\
        );

    \I__11183\ : InMux
    port map (
            O => \N__47290\,
            I => \N__47281\
        );

    \I__11182\ : LocalMux
    port map (
            O => \N__47287\,
            I => \N__47278\
        );

    \I__11181\ : Odrv4
    port map (
            O => \N__47284\,
            I => n8_adj_723
        );

    \I__11180\ : LocalMux
    port map (
            O => \N__47281\,
            I => n8_adj_723
        );

    \I__11179\ : Odrv4
    port map (
            O => \N__47278\,
            I => n8_adj_723
        );

    \I__11178\ : InMux
    port map (
            O => \N__47271\,
            I => \N__47268\
        );

    \I__11177\ : LocalMux
    port map (
            O => \N__47268\,
            I => n4_adj_778
        );

    \I__11176\ : InMux
    port map (
            O => \N__47265\,
            I => \N__47260\
        );

    \I__11175\ : InMux
    port map (
            O => \N__47264\,
            I => \N__47255\
        );

    \I__11174\ : InMux
    port map (
            O => \N__47263\,
            I => \N__47255\
        );

    \I__11173\ : LocalMux
    port map (
            O => \N__47260\,
            I => \N__47252\
        );

    \I__11172\ : LocalMux
    port map (
            O => \N__47255\,
            I => \N__47249\
        );

    \I__11171\ : Span4Mux_h
    port map (
            O => \N__47252\,
            I => \N__47246\
        );

    \I__11170\ : Odrv4
    port map (
            O => \N__47249\,
            I => n7142
        );

    \I__11169\ : Odrv4
    port map (
            O => \N__47246\,
            I => n7142
        );

    \I__11168\ : CascadeMux
    port map (
            O => \N__47241\,
            I => \n7142_cascade_\
        );

    \I__11167\ : InMux
    port map (
            O => \N__47238\,
            I => \N__47232\
        );

    \I__11166\ : InMux
    port map (
            O => \N__47237\,
            I => \N__47226\
        );

    \I__11165\ : InMux
    port map (
            O => \N__47236\,
            I => \N__47220\
        );

    \I__11164\ : InMux
    port map (
            O => \N__47235\,
            I => \N__47220\
        );

    \I__11163\ : LocalMux
    port map (
            O => \N__47232\,
            I => \N__47217\
        );

    \I__11162\ : InMux
    port map (
            O => \N__47231\,
            I => \N__47212\
        );

    \I__11161\ : InMux
    port map (
            O => \N__47230\,
            I => \N__47212\
        );

    \I__11160\ : InMux
    port map (
            O => \N__47229\,
            I => \N__47209\
        );

    \I__11159\ : LocalMux
    port map (
            O => \N__47226\,
            I => \N__47206\
        );

    \I__11158\ : InMux
    port map (
            O => \N__47225\,
            I => \N__47203\
        );

    \I__11157\ : LocalMux
    port map (
            O => \N__47220\,
            I => \N__47200\
        );

    \I__11156\ : Span4Mux_h
    port map (
            O => \N__47217\,
            I => \N__47197\
        );

    \I__11155\ : LocalMux
    port map (
            O => \N__47212\,
            I => \N__47194\
        );

    \I__11154\ : LocalMux
    port map (
            O => \N__47209\,
            I => counter_7
        );

    \I__11153\ : Odrv4
    port map (
            O => \N__47206\,
            I => counter_7
        );

    \I__11152\ : LocalMux
    port map (
            O => \N__47203\,
            I => counter_7
        );

    \I__11151\ : Odrv4
    port map (
            O => \N__47200\,
            I => counter_7
        );

    \I__11150\ : Odrv4
    port map (
            O => \N__47197\,
            I => counter_7
        );

    \I__11149\ : Odrv12
    port map (
            O => \N__47194\,
            I => counter_7
        );

    \I__11148\ : CascadeMux
    port map (
            O => \N__47181\,
            I => \N__47177\
        );

    \I__11147\ : CascadeMux
    port map (
            O => \N__47180\,
            I => \N__47173\
        );

    \I__11146\ : InMux
    port map (
            O => \N__47177\,
            I => \N__47169\
        );

    \I__11145\ : CascadeMux
    port map (
            O => \N__47176\,
            I => \N__47165\
        );

    \I__11144\ : InMux
    port map (
            O => \N__47173\,
            I => \N__47160\
        );

    \I__11143\ : CascadeMux
    port map (
            O => \N__47172\,
            I => \N__47157\
        );

    \I__11142\ : LocalMux
    port map (
            O => \N__47169\,
            I => \N__47153\
        );

    \I__11141\ : InMux
    port map (
            O => \N__47168\,
            I => \N__47148\
        );

    \I__11140\ : InMux
    port map (
            O => \N__47165\,
            I => \N__47148\
        );

    \I__11139\ : InMux
    port map (
            O => \N__47164\,
            I => \N__47143\
        );

    \I__11138\ : InMux
    port map (
            O => \N__47163\,
            I => \N__47143\
        );

    \I__11137\ : LocalMux
    port map (
            O => \N__47160\,
            I => \N__47140\
        );

    \I__11136\ : InMux
    port map (
            O => \N__47157\,
            I => \N__47137\
        );

    \I__11135\ : InMux
    port map (
            O => \N__47156\,
            I => \N__47134\
        );

    \I__11134\ : Span4Mux_v
    port map (
            O => \N__47153\,
            I => \N__47129\
        );

    \I__11133\ : LocalMux
    port map (
            O => \N__47148\,
            I => \N__47129\
        );

    \I__11132\ : LocalMux
    port map (
            O => \N__47143\,
            I => \N__47126\
        );

    \I__11131\ : Odrv4
    port map (
            O => \N__47140\,
            I => counter_6
        );

    \I__11130\ : LocalMux
    port map (
            O => \N__47137\,
            I => counter_6
        );

    \I__11129\ : LocalMux
    port map (
            O => \N__47134\,
            I => counter_6
        );

    \I__11128\ : Odrv4
    port map (
            O => \N__47129\,
            I => counter_6
        );

    \I__11127\ : Odrv12
    port map (
            O => \N__47126\,
            I => counter_6
        );

    \I__11126\ : SRMux
    port map (
            O => \N__47115\,
            I => \N__47112\
        );

    \I__11125\ : LocalMux
    port map (
            O => \N__47112\,
            I => \N__47109\
        );

    \I__11124\ : Span4Mux_v
    port map (
            O => \N__47109\,
            I => \N__47106\
        );

    \I__11123\ : Sp12to4
    port map (
            O => \N__47106\,
            I => \N__47102\
        );

    \I__11122\ : InMux
    port map (
            O => \N__47105\,
            I => \N__47099\
        );

    \I__11121\ : Span12Mux_s6_h
    port map (
            O => \N__47102\,
            I => \N__47096\
        );

    \I__11120\ : LocalMux
    port map (
            O => \N__47099\,
            I => \N__47093\
        );

    \I__11119\ : Odrv12
    port map (
            O => \N__47096\,
            I => n73
        );

    \I__11118\ : Odrv12
    port map (
            O => \N__47093\,
            I => n73
        );

    \I__11117\ : InMux
    port map (
            O => \N__47088\,
            I => \N__47085\
        );

    \I__11116\ : LocalMux
    port map (
            O => \N__47085\,
            I => \N__47081\
        );

    \I__11115\ : InMux
    port map (
            O => \N__47084\,
            I => \N__47078\
        );

    \I__11114\ : Span4Mux_v
    port map (
            O => \N__47081\,
            I => \N__47075\
        );

    \I__11113\ : LocalMux
    port map (
            O => \N__47078\,
            I => \N__47072\
        );

    \I__11112\ : Span4Mux_v
    port map (
            O => \N__47075\,
            I => \N__47069\
        );

    \I__11111\ : Span4Mux_v
    port map (
            O => \N__47072\,
            I => \N__47066\
        );

    \I__11110\ : Span4Mux_v
    port map (
            O => \N__47069\,
            I => \N__47063\
        );

    \I__11109\ : Span4Mux_v
    port map (
            O => \N__47066\,
            I => \N__47060\
        );

    \I__11108\ : Sp12to4
    port map (
            O => \N__47063\,
            I => \N__47057\
        );

    \I__11107\ : Span4Mux_v
    port map (
            O => \N__47060\,
            I => \N__47054\
        );

    \I__11106\ : Span12Mux_h
    port map (
            O => \N__47057\,
            I => \N__47051\
        );

    \I__11105\ : Span4Mux_h
    port map (
            O => \N__47054\,
            I => \N__47048\
        );

    \I__11104\ : Odrv12
    port map (
            O => \N__47051\,
            I => pin_in_7
        );

    \I__11103\ : Odrv4
    port map (
            O => \N__47048\,
            I => pin_in_7
        );

    \I__11102\ : InMux
    port map (
            O => \N__47043\,
            I => \N__47040\
        );

    \I__11101\ : LocalMux
    port map (
            O => \N__47040\,
            I => n2385
        );

    \I__11100\ : CascadeMux
    port map (
            O => \N__47037\,
            I => \n12123_cascade_\
        );

    \I__11099\ : InMux
    port map (
            O => \N__47034\,
            I => \N__47031\
        );

    \I__11098\ : LocalMux
    port map (
            O => \N__47031\,
            I => \N__47028\
        );

    \I__11097\ : Span4Mux_v
    port map (
            O => \N__47028\,
            I => \N__47025\
        );

    \I__11096\ : Odrv4
    port map (
            O => \N__47025\,
            I => n48_adj_771
        );

    \I__11095\ : InMux
    port map (
            O => \N__47022\,
            I => \N__47019\
        );

    \I__11094\ : LocalMux
    port map (
            O => \N__47019\,
            I => \N__47016\
        );

    \I__11093\ : Span4Mux_v
    port map (
            O => \N__47016\,
            I => \N__47012\
        );

    \I__11092\ : InMux
    port map (
            O => \N__47015\,
            I => \N__47009\
        );

    \I__11091\ : Sp12to4
    port map (
            O => \N__47012\,
            I => \N__47006\
        );

    \I__11090\ : LocalMux
    port map (
            O => \N__47009\,
            I => \N__47003\
        );

    \I__11089\ : Span12Mux_h
    port map (
            O => \N__47006\,
            I => \N__46998\
        );

    \I__11088\ : Span12Mux_s7_h
    port map (
            O => \N__47003\,
            I => \N__46998\
        );

    \I__11087\ : Span12Mux_v
    port map (
            O => \N__46998\,
            I => \N__46995\
        );

    \I__11086\ : Odrv12
    port map (
            O => \N__46995\,
            I => pin_in_4
        );

    \I__11085\ : InMux
    port map (
            O => \N__46992\,
            I => \N__46989\
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__46989\,
            I => n2313
        );

    \I__11083\ : InMux
    port map (
            O => \N__46986\,
            I => n10516
        );

    \I__11082\ : CascadeMux
    port map (
            O => \N__46983\,
            I => \n8_adj_763_cascade_\
        );

    \I__11081\ : InMux
    port map (
            O => \N__46980\,
            I => \N__46974\
        );

    \I__11080\ : CascadeMux
    port map (
            O => \N__46979\,
            I => \N__46971\
        );

    \I__11079\ : CascadeMux
    port map (
            O => \N__46978\,
            I => \N__46966\
        );

    \I__11078\ : InMux
    port map (
            O => \N__46977\,
            I => \N__46960\
        );

    \I__11077\ : LocalMux
    port map (
            O => \N__46974\,
            I => \N__46955\
        );

    \I__11076\ : InMux
    port map (
            O => \N__46971\,
            I => \N__46950\
        );

    \I__11075\ : InMux
    port map (
            O => \N__46970\,
            I => \N__46950\
        );

    \I__11074\ : InMux
    port map (
            O => \N__46969\,
            I => \N__46945\
        );

    \I__11073\ : InMux
    port map (
            O => \N__46966\,
            I => \N__46945\
        );

    \I__11072\ : InMux
    port map (
            O => \N__46965\,
            I => \N__46937\
        );

    \I__11071\ : InMux
    port map (
            O => \N__46964\,
            I => \N__46932\
        );

    \I__11070\ : InMux
    port map (
            O => \N__46963\,
            I => \N__46932\
        );

    \I__11069\ : LocalMux
    port map (
            O => \N__46960\,
            I => \N__46924\
        );

    \I__11068\ : CascadeMux
    port map (
            O => \N__46959\,
            I => \N__46920\
        );

    \I__11067\ : CascadeMux
    port map (
            O => \N__46958\,
            I => \N__46917\
        );

    \I__11066\ : Span4Mux_v
    port map (
            O => \N__46955\,
            I => \N__46908\
        );

    \I__11065\ : LocalMux
    port map (
            O => \N__46950\,
            I => \N__46908\
        );

    \I__11064\ : LocalMux
    port map (
            O => \N__46945\,
            I => \N__46908\
        );

    \I__11063\ : InMux
    port map (
            O => \N__46944\,
            I => \N__46905\
        );

    \I__11062\ : InMux
    port map (
            O => \N__46943\,
            I => \N__46898\
        );

    \I__11061\ : InMux
    port map (
            O => \N__46942\,
            I => \N__46898\
        );

    \I__11060\ : InMux
    port map (
            O => \N__46941\,
            I => \N__46898\
        );

    \I__11059\ : InMux
    port map (
            O => \N__46940\,
            I => \N__46895\
        );

    \I__11058\ : LocalMux
    port map (
            O => \N__46937\,
            I => \N__46890\
        );

    \I__11057\ : LocalMux
    port map (
            O => \N__46932\,
            I => \N__46890\
        );

    \I__11056\ : CascadeMux
    port map (
            O => \N__46931\,
            I => \N__46887\
        );

    \I__11055\ : CascadeMux
    port map (
            O => \N__46930\,
            I => \N__46883\
        );

    \I__11054\ : CascadeMux
    port map (
            O => \N__46929\,
            I => \N__46879\
        );

    \I__11053\ : CascadeMux
    port map (
            O => \N__46928\,
            I => \N__46875\
        );

    \I__11052\ : CascadeMux
    port map (
            O => \N__46927\,
            I => \N__46872\
        );

    \I__11051\ : Sp12to4
    port map (
            O => \N__46924\,
            I => \N__46868\
        );

    \I__11050\ : InMux
    port map (
            O => \N__46923\,
            I => \N__46865\
        );

    \I__11049\ : InMux
    port map (
            O => \N__46920\,
            I => \N__46862\
        );

    \I__11048\ : InMux
    port map (
            O => \N__46917\,
            I => \N__46859\
        );

    \I__11047\ : InMux
    port map (
            O => \N__46916\,
            I => \N__46856\
        );

    \I__11046\ : InMux
    port map (
            O => \N__46915\,
            I => \N__46853\
        );

    \I__11045\ : Span4Mux_v
    port map (
            O => \N__46908\,
            I => \N__46850\
        );

    \I__11044\ : LocalMux
    port map (
            O => \N__46905\,
            I => \N__46841\
        );

    \I__11043\ : LocalMux
    port map (
            O => \N__46898\,
            I => \N__46841\
        );

    \I__11042\ : LocalMux
    port map (
            O => \N__46895\,
            I => \N__46841\
        );

    \I__11041\ : Span4Mux_h
    port map (
            O => \N__46890\,
            I => \N__46841\
        );

    \I__11040\ : InMux
    port map (
            O => \N__46887\,
            I => \N__46826\
        );

    \I__11039\ : InMux
    port map (
            O => \N__46886\,
            I => \N__46826\
        );

    \I__11038\ : InMux
    port map (
            O => \N__46883\,
            I => \N__46826\
        );

    \I__11037\ : InMux
    port map (
            O => \N__46882\,
            I => \N__46826\
        );

    \I__11036\ : InMux
    port map (
            O => \N__46879\,
            I => \N__46826\
        );

    \I__11035\ : InMux
    port map (
            O => \N__46878\,
            I => \N__46826\
        );

    \I__11034\ : InMux
    port map (
            O => \N__46875\,
            I => \N__46826\
        );

    \I__11033\ : InMux
    port map (
            O => \N__46872\,
            I => \N__46821\
        );

    \I__11032\ : InMux
    port map (
            O => \N__46871\,
            I => \N__46821\
        );

    \I__11031\ : Span12Mux_v
    port map (
            O => \N__46868\,
            I => \N__46818\
        );

    \I__11030\ : LocalMux
    port map (
            O => \N__46865\,
            I => \N__46807\
        );

    \I__11029\ : LocalMux
    port map (
            O => \N__46862\,
            I => \N__46807\
        );

    \I__11028\ : LocalMux
    port map (
            O => \N__46859\,
            I => \N__46807\
        );

    \I__11027\ : LocalMux
    port map (
            O => \N__46856\,
            I => \N__46807\
        );

    \I__11026\ : LocalMux
    port map (
            O => \N__46853\,
            I => \N__46807\
        );

    \I__11025\ : Span4Mux_h
    port map (
            O => \N__46850\,
            I => \N__46804\
        );

    \I__11024\ : Span4Mux_h
    port map (
            O => \N__46841\,
            I => \N__46801\
        );

    \I__11023\ : LocalMux
    port map (
            O => \N__46826\,
            I => \current_pin_7__N_155\
        );

    \I__11022\ : LocalMux
    port map (
            O => \N__46821\,
            I => \current_pin_7__N_155\
        );

    \I__11021\ : Odrv12
    port map (
            O => \N__46818\,
            I => \current_pin_7__N_155\
        );

    \I__11020\ : Odrv12
    port map (
            O => \N__46807\,
            I => \current_pin_7__N_155\
        );

    \I__11019\ : Odrv4
    port map (
            O => \N__46804\,
            I => \current_pin_7__N_155\
        );

    \I__11018\ : Odrv4
    port map (
            O => \N__46801\,
            I => \current_pin_7__N_155\
        );

    \I__11017\ : InMux
    port map (
            O => \N__46788\,
            I => \N__46783\
        );

    \I__11016\ : InMux
    port map (
            O => \N__46787\,
            I => \N__46778\
        );

    \I__11015\ : InMux
    port map (
            O => \N__46786\,
            I => \N__46778\
        );

    \I__11014\ : LocalMux
    port map (
            O => \N__46783\,
            I => \N__46769\
        );

    \I__11013\ : LocalMux
    port map (
            O => \N__46778\,
            I => \N__46769\
        );

    \I__11012\ : InMux
    port map (
            O => \N__46777\,
            I => \N__46766\
        );

    \I__11011\ : InMux
    port map (
            O => \N__46776\,
            I => \N__46763\
        );

    \I__11010\ : InMux
    port map (
            O => \N__46775\,
            I => \N__46758\
        );

    \I__11009\ : InMux
    port map (
            O => \N__46774\,
            I => \N__46758\
        );

    \I__11008\ : Span4Mux_h
    port map (
            O => \N__46769\,
            I => \N__46755\
        );

    \I__11007\ : LocalMux
    port map (
            O => \N__46766\,
            I => n7_adj_719
        );

    \I__11006\ : LocalMux
    port map (
            O => \N__46763\,
            I => n7_adj_719
        );

    \I__11005\ : LocalMux
    port map (
            O => \N__46758\,
            I => n7_adj_719
        );

    \I__11004\ : Odrv4
    port map (
            O => \N__46755\,
            I => n7_adj_719
        );

    \I__11003\ : CascadeMux
    port map (
            O => \N__46746\,
            I => \N__46740\
        );

    \I__11002\ : CascadeMux
    port map (
            O => \N__46745\,
            I => \N__46737\
        );

    \I__11001\ : InMux
    port map (
            O => \N__46744\,
            I => \N__46734\
        );

    \I__11000\ : InMux
    port map (
            O => \N__46743\,
            I => \N__46729\
        );

    \I__10999\ : InMux
    port map (
            O => \N__46740\,
            I => \N__46729\
        );

    \I__10998\ : InMux
    port map (
            O => \N__46737\,
            I => \N__46726\
        );

    \I__10997\ : LocalMux
    port map (
            O => \N__46734\,
            I => \N__46723\
        );

    \I__10996\ : LocalMux
    port map (
            O => \N__46729\,
            I => \N__46719\
        );

    \I__10995\ : LocalMux
    port map (
            O => \N__46726\,
            I => \N__46716\
        );

    \I__10994\ : Span4Mux_h
    port map (
            O => \N__46723\,
            I => \N__46713\
        );

    \I__10993\ : InMux
    port map (
            O => \N__46722\,
            I => \N__46710\
        );

    \I__10992\ : Span4Mux_h
    port map (
            O => \N__46719\,
            I => \N__46705\
        );

    \I__10991\ : Span4Mux_v
    port map (
            O => \N__46716\,
            I => \N__46705\
        );

    \I__10990\ : Span4Mux_h
    port map (
            O => \N__46713\,
            I => \N__46702\
        );

    \I__10989\ : LocalMux
    port map (
            O => \N__46710\,
            I => n21
        );

    \I__10988\ : Odrv4
    port map (
            O => \N__46705\,
            I => n21
        );

    \I__10987\ : Odrv4
    port map (
            O => \N__46702\,
            I => n21
        );

    \I__10986\ : CascadeMux
    port map (
            O => \N__46695\,
            I => \current_pin_7__N_155_cascade_\
        );

    \I__10985\ : CascadeMux
    port map (
            O => \N__46692\,
            I => \N__46689\
        );

    \I__10984\ : InMux
    port map (
            O => \N__46689\,
            I => \N__46684\
        );

    \I__10983\ : CascadeMux
    port map (
            O => \N__46688\,
            I => \N__46680\
        );

    \I__10982\ : InMux
    port map (
            O => \N__46687\,
            I => \N__46674\
        );

    \I__10981\ : LocalMux
    port map (
            O => \N__46684\,
            I => \N__46671\
        );

    \I__10980\ : InMux
    port map (
            O => \N__46683\,
            I => \N__46666\
        );

    \I__10979\ : InMux
    port map (
            O => \N__46680\,
            I => \N__46663\
        );

    \I__10978\ : InMux
    port map (
            O => \N__46679\,
            I => \N__46658\
        );

    \I__10977\ : InMux
    port map (
            O => \N__46678\,
            I => \N__46658\
        );

    \I__10976\ : InMux
    port map (
            O => \N__46677\,
            I => \N__46654\
        );

    \I__10975\ : LocalMux
    port map (
            O => \N__46674\,
            I => \N__46651\
        );

    \I__10974\ : Span4Mux_v
    port map (
            O => \N__46671\,
            I => \N__46648\
        );

    \I__10973\ : InMux
    port map (
            O => \N__46670\,
            I => \N__46643\
        );

    \I__10972\ : InMux
    port map (
            O => \N__46669\,
            I => \N__46643\
        );

    \I__10971\ : LocalMux
    port map (
            O => \N__46666\,
            I => \N__46639\
        );

    \I__10970\ : LocalMux
    port map (
            O => \N__46663\,
            I => \N__46634\
        );

    \I__10969\ : LocalMux
    port map (
            O => \N__46658\,
            I => \N__46634\
        );

    \I__10968\ : InMux
    port map (
            O => \N__46657\,
            I => \N__46631\
        );

    \I__10967\ : LocalMux
    port map (
            O => \N__46654\,
            I => \N__46626\
        );

    \I__10966\ : Span4Mux_v
    port map (
            O => \N__46651\,
            I => \N__46626\
        );

    \I__10965\ : Span4Mux_h
    port map (
            O => \N__46648\,
            I => \N__46621\
        );

    \I__10964\ : LocalMux
    port map (
            O => \N__46643\,
            I => \N__46621\
        );

    \I__10963\ : InMux
    port map (
            O => \N__46642\,
            I => \N__46618\
        );

    \I__10962\ : Span4Mux_h
    port map (
            O => \N__46639\,
            I => \N__46613\
        );

    \I__10961\ : Span4Mux_h
    port map (
            O => \N__46634\,
            I => \N__46613\
        );

    \I__10960\ : LocalMux
    port map (
            O => \N__46631\,
            I => n7166
        );

    \I__10959\ : Odrv4
    port map (
            O => \N__46626\,
            I => n7166
        );

    \I__10958\ : Odrv4
    port map (
            O => \N__46621\,
            I => n7166
        );

    \I__10957\ : LocalMux
    port map (
            O => \N__46618\,
            I => n7166
        );

    \I__10956\ : Odrv4
    port map (
            O => \N__46613\,
            I => n7166
        );

    \I__10955\ : CascadeMux
    port map (
            O => \N__46602\,
            I => \N__46599\
        );

    \I__10954\ : InMux
    port map (
            O => \N__46599\,
            I => \N__46596\
        );

    \I__10953\ : LocalMux
    port map (
            O => \N__46596\,
            I => \N__46593\
        );

    \I__10952\ : Span4Mux_h
    port map (
            O => \N__46593\,
            I => \N__46589\
        );

    \I__10951\ : InMux
    port map (
            O => \N__46592\,
            I => \N__46586\
        );

    \I__10950\ : Odrv4
    port map (
            O => \N__46589\,
            I => n6180
        );

    \I__10949\ : LocalMux
    port map (
            O => \N__46586\,
            I => n6180
        );

    \I__10948\ : InMux
    port map (
            O => \N__46581\,
            I => \N__46571\
        );

    \I__10947\ : InMux
    port map (
            O => \N__46580\,
            I => \N__46571\
        );

    \I__10946\ : InMux
    port map (
            O => \N__46579\,
            I => \N__46571\
        );

    \I__10945\ : InMux
    port map (
            O => \N__46578\,
            I => \N__46564\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__46571\,
            I => \N__46561\
        );

    \I__10943\ : InMux
    port map (
            O => \N__46570\,
            I => \N__46552\
        );

    \I__10942\ : InMux
    port map (
            O => \N__46569\,
            I => \N__46552\
        );

    \I__10941\ : InMux
    port map (
            O => \N__46568\,
            I => \N__46552\
        );

    \I__10940\ : InMux
    port map (
            O => \N__46567\,
            I => \N__46552\
        );

    \I__10939\ : LocalMux
    port map (
            O => \N__46564\,
            I => \N__46549\
        );

    \I__10938\ : Odrv4
    port map (
            O => \N__46561\,
            I => n6971
        );

    \I__10937\ : LocalMux
    port map (
            O => \N__46552\,
            I => n6971
        );

    \I__10936\ : Odrv4
    port map (
            O => \N__46549\,
            I => n6971
        );

    \I__10935\ : InMux
    port map (
            O => \N__46542\,
            I => \N__46539\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__46539\,
            I => n12135
        );

    \I__10933\ : InMux
    port map (
            O => \N__46536\,
            I => \N__46531\
        );

    \I__10932\ : InMux
    port map (
            O => \N__46535\,
            I => \N__46525\
        );

    \I__10931\ : InMux
    port map (
            O => \N__46534\,
            I => \N__46520\
        );

    \I__10930\ : LocalMux
    port map (
            O => \N__46531\,
            I => \N__46512\
        );

    \I__10929\ : InMux
    port map (
            O => \N__46530\,
            I => \N__46509\
        );

    \I__10928\ : InMux
    port map (
            O => \N__46529\,
            I => \N__46506\
        );

    \I__10927\ : InMux
    port map (
            O => \N__46528\,
            I => \N__46503\
        );

    \I__10926\ : LocalMux
    port map (
            O => \N__46525\,
            I => \N__46500\
        );

    \I__10925\ : InMux
    port map (
            O => \N__46524\,
            I => \N__46495\
        );

    \I__10924\ : InMux
    port map (
            O => \N__46523\,
            I => \N__46495\
        );

    \I__10923\ : LocalMux
    port map (
            O => \N__46520\,
            I => \N__46492\
        );

    \I__10922\ : InMux
    port map (
            O => \N__46519\,
            I => \N__46489\
        );

    \I__10921\ : InMux
    port map (
            O => \N__46518\,
            I => \N__46484\
        );

    \I__10920\ : InMux
    port map (
            O => \N__46517\,
            I => \N__46476\
        );

    \I__10919\ : InMux
    port map (
            O => \N__46516\,
            I => \N__46476\
        );

    \I__10918\ : InMux
    port map (
            O => \N__46515\,
            I => \N__46472\
        );

    \I__10917\ : Span4Mux_v
    port map (
            O => \N__46512\,
            I => \N__46467\
        );

    \I__10916\ : LocalMux
    port map (
            O => \N__46509\,
            I => \N__46467\
        );

    \I__10915\ : LocalMux
    port map (
            O => \N__46506\,
            I => \N__46464\
        );

    \I__10914\ : LocalMux
    port map (
            O => \N__46503\,
            I => \N__46457\
        );

    \I__10913\ : Span4Mux_h
    port map (
            O => \N__46500\,
            I => \N__46457\
        );

    \I__10912\ : LocalMux
    port map (
            O => \N__46495\,
            I => \N__46457\
        );

    \I__10911\ : Span4Mux_h
    port map (
            O => \N__46492\,
            I => \N__46452\
        );

    \I__10910\ : LocalMux
    port map (
            O => \N__46489\,
            I => \N__46452\
        );

    \I__10909\ : InMux
    port map (
            O => \N__46488\,
            I => \N__46445\
        );

    \I__10908\ : InMux
    port map (
            O => \N__46487\,
            I => \N__46442\
        );

    \I__10907\ : LocalMux
    port map (
            O => \N__46484\,
            I => \N__46439\
        );

    \I__10906\ : InMux
    port map (
            O => \N__46483\,
            I => \N__46436\
        );

    \I__10905\ : InMux
    port map (
            O => \N__46482\,
            I => \N__46431\
        );

    \I__10904\ : InMux
    port map (
            O => \N__46481\,
            I => \N__46431\
        );

    \I__10903\ : LocalMux
    port map (
            O => \N__46476\,
            I => \N__46428\
        );

    \I__10902\ : InMux
    port map (
            O => \N__46475\,
            I => \N__46425\
        );

    \I__10901\ : LocalMux
    port map (
            O => \N__46472\,
            I => \N__46422\
        );

    \I__10900\ : Span4Mux_h
    port map (
            O => \N__46467\,
            I => \N__46417\
        );

    \I__10899\ : Span4Mux_v
    port map (
            O => \N__46464\,
            I => \N__46417\
        );

    \I__10898\ : Span4Mux_v
    port map (
            O => \N__46457\,
            I => \N__46414\
        );

    \I__10897\ : Span4Mux_v
    port map (
            O => \N__46452\,
            I => \N__46411\
        );

    \I__10896\ : InMux
    port map (
            O => \N__46451\,
            I => \N__46408\
        );

    \I__10895\ : InMux
    port map (
            O => \N__46450\,
            I => \N__46401\
        );

    \I__10894\ : InMux
    port map (
            O => \N__46449\,
            I => \N__46401\
        );

    \I__10893\ : InMux
    port map (
            O => \N__46448\,
            I => \N__46401\
        );

    \I__10892\ : LocalMux
    port map (
            O => \N__46445\,
            I => \N__46396\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__46442\,
            I => \N__46396\
        );

    \I__10890\ : Span4Mux_v
    port map (
            O => \N__46439\,
            I => \N__46393\
        );

    \I__10889\ : LocalMux
    port map (
            O => \N__46436\,
            I => \N__46384\
        );

    \I__10888\ : LocalMux
    port map (
            O => \N__46431\,
            I => \N__46384\
        );

    \I__10887\ : Span4Mux_h
    port map (
            O => \N__46428\,
            I => \N__46384\
        );

    \I__10886\ : LocalMux
    port map (
            O => \N__46425\,
            I => \N__46384\
        );

    \I__10885\ : Span12Mux_v
    port map (
            O => \N__46422\,
            I => \N__46381\
        );

    \I__10884\ : Span4Mux_h
    port map (
            O => \N__46417\,
            I => \N__46376\
        );

    \I__10883\ : Span4Mux_h
    port map (
            O => \N__46414\,
            I => \N__46376\
        );

    \I__10882\ : Span4Mux_h
    port map (
            O => \N__46411\,
            I => \N__46371\
        );

    \I__10881\ : LocalMux
    port map (
            O => \N__46408\,
            I => \N__46371\
        );

    \I__10880\ : LocalMux
    port map (
            O => \N__46401\,
            I => n149
        );

    \I__10879\ : Odrv12
    port map (
            O => \N__46396\,
            I => n149
        );

    \I__10878\ : Odrv4
    port map (
            O => \N__46393\,
            I => n149
        );

    \I__10877\ : Odrv4
    port map (
            O => \N__46384\,
            I => n149
        );

    \I__10876\ : Odrv12
    port map (
            O => \N__46381\,
            I => n149
        );

    \I__10875\ : Odrv4
    port map (
            O => \N__46376\,
            I => n149
        );

    \I__10874\ : Odrv4
    port map (
            O => \N__46371\,
            I => n149
        );

    \I__10873\ : InMux
    port map (
            O => \N__46356\,
            I => n10572
        );

    \I__10872\ : InMux
    port map (
            O => \N__46353\,
            I => \N__46349\
        );

    \I__10871\ : InMux
    port map (
            O => \N__46352\,
            I => \N__46346\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__46349\,
            I => blink_counter_25
        );

    \I__10869\ : LocalMux
    port map (
            O => \N__46346\,
            I => blink_counter_25
        );

    \I__10868\ : InMux
    port map (
            O => \N__46341\,
            I => \N__46338\
        );

    \I__10867\ : LocalMux
    port map (
            O => \N__46338\,
            I => n45
        );

    \I__10866\ : InMux
    port map (
            O => \N__46335\,
            I => \bfn_16_15_0_\
        );

    \I__10865\ : InMux
    port map (
            O => \N__46332\,
            I => n10510
        );

    \I__10864\ : InMux
    port map (
            O => \N__46329\,
            I => n10511
        );

    \I__10863\ : InMux
    port map (
            O => \N__46326\,
            I => n10512
        );

    \I__10862\ : InMux
    port map (
            O => \N__46323\,
            I => n10513
        );

    \I__10861\ : InMux
    port map (
            O => \N__46320\,
            I => n10514
        );

    \I__10860\ : InMux
    port map (
            O => \N__46317\,
            I => n10515
        );

    \I__10859\ : InMux
    port map (
            O => \N__46314\,
            I => \N__46311\
        );

    \I__10858\ : LocalMux
    port map (
            O => \N__46311\,
            I => n9
        );

    \I__10857\ : InMux
    port map (
            O => \N__46308\,
            I => n10564
        );

    \I__10856\ : InMux
    port map (
            O => \N__46305\,
            I => \N__46302\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__46302\,
            I => n8_adj_755
        );

    \I__10854\ : InMux
    port map (
            O => \N__46299\,
            I => n10565
        );

    \I__10853\ : InMux
    port map (
            O => \N__46296\,
            I => \N__46293\
        );

    \I__10852\ : LocalMux
    port map (
            O => \N__46293\,
            I => n7
        );

    \I__10851\ : InMux
    port map (
            O => \N__46290\,
            I => n10566
        );

    \I__10850\ : InMux
    port map (
            O => \N__46287\,
            I => \N__46284\
        );

    \I__10849\ : LocalMux
    port map (
            O => \N__46284\,
            I => n6_adj_756
        );

    \I__10848\ : InMux
    port map (
            O => \N__46281\,
            I => n10567
        );

    \I__10847\ : CascadeMux
    port map (
            O => \N__46278\,
            I => \N__46275\
        );

    \I__10846\ : InMux
    port map (
            O => \N__46275\,
            I => \N__46268\
        );

    \I__10845\ : InMux
    port map (
            O => \N__46274\,
            I => \N__46268\
        );

    \I__10844\ : InMux
    port map (
            O => \N__46273\,
            I => \N__46265\
        );

    \I__10843\ : LocalMux
    port map (
            O => \N__46268\,
            I => blink_counter_21
        );

    \I__10842\ : LocalMux
    port map (
            O => \N__46265\,
            I => blink_counter_21
        );

    \I__10841\ : InMux
    port map (
            O => \N__46260\,
            I => n10568
        );

    \I__10840\ : InMux
    port map (
            O => \N__46257\,
            I => \N__46250\
        );

    \I__10839\ : InMux
    port map (
            O => \N__46256\,
            I => \N__46250\
        );

    \I__10838\ : InMux
    port map (
            O => \N__46255\,
            I => \N__46247\
        );

    \I__10837\ : LocalMux
    port map (
            O => \N__46250\,
            I => blink_counter_22
        );

    \I__10836\ : LocalMux
    port map (
            O => \N__46247\,
            I => blink_counter_22
        );

    \I__10835\ : InMux
    port map (
            O => \N__46242\,
            I => n10569
        );

    \I__10834\ : CascadeMux
    port map (
            O => \N__46239\,
            I => \N__46235\
        );

    \I__10833\ : InMux
    port map (
            O => \N__46238\,
            I => \N__46229\
        );

    \I__10832\ : InMux
    port map (
            O => \N__46235\,
            I => \N__46229\
        );

    \I__10831\ : InMux
    port map (
            O => \N__46234\,
            I => \N__46226\
        );

    \I__10830\ : LocalMux
    port map (
            O => \N__46229\,
            I => blink_counter_23
        );

    \I__10829\ : LocalMux
    port map (
            O => \N__46226\,
            I => blink_counter_23
        );

    \I__10828\ : InMux
    port map (
            O => \N__46221\,
            I => n10570
        );

    \I__10827\ : InMux
    port map (
            O => \N__46218\,
            I => \N__46211\
        );

    \I__10826\ : InMux
    port map (
            O => \N__46217\,
            I => \N__46211\
        );

    \I__10825\ : InMux
    port map (
            O => \N__46216\,
            I => \N__46208\
        );

    \I__10824\ : LocalMux
    port map (
            O => \N__46211\,
            I => blink_counter_24
        );

    \I__10823\ : LocalMux
    port map (
            O => \N__46208\,
            I => blink_counter_24
        );

    \I__10822\ : InMux
    port map (
            O => \N__46203\,
            I => \bfn_15_29_0_\
        );

    \I__10821\ : InMux
    port map (
            O => \N__46200\,
            I => \N__46197\
        );

    \I__10820\ : LocalMux
    port map (
            O => \N__46197\,
            I => n18
        );

    \I__10819\ : InMux
    port map (
            O => \N__46194\,
            I => \bfn_15_27_0_\
        );

    \I__10818\ : InMux
    port map (
            O => \N__46191\,
            I => \N__46188\
        );

    \I__10817\ : LocalMux
    port map (
            O => \N__46188\,
            I => n17
        );

    \I__10816\ : InMux
    port map (
            O => \N__46185\,
            I => n10556
        );

    \I__10815\ : InMux
    port map (
            O => \N__46182\,
            I => \N__46179\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__46179\,
            I => n16
        );

    \I__10813\ : InMux
    port map (
            O => \N__46176\,
            I => n10557
        );

    \I__10812\ : InMux
    port map (
            O => \N__46173\,
            I => \N__46170\
        );

    \I__10811\ : LocalMux
    port map (
            O => \N__46170\,
            I => n15_adj_759
        );

    \I__10810\ : InMux
    port map (
            O => \N__46167\,
            I => n10558
        );

    \I__10809\ : InMux
    port map (
            O => \N__46164\,
            I => \N__46161\
        );

    \I__10808\ : LocalMux
    port map (
            O => \N__46161\,
            I => n14_adj_745
        );

    \I__10807\ : InMux
    port map (
            O => \N__46158\,
            I => n10559
        );

    \I__10806\ : InMux
    port map (
            O => \N__46155\,
            I => \N__46152\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__46152\,
            I => n13
        );

    \I__10804\ : InMux
    port map (
            O => \N__46149\,
            I => n10560
        );

    \I__10803\ : InMux
    port map (
            O => \N__46146\,
            I => \N__46143\
        );

    \I__10802\ : LocalMux
    port map (
            O => \N__46143\,
            I => n12
        );

    \I__10801\ : InMux
    port map (
            O => \N__46140\,
            I => n10561
        );

    \I__10800\ : InMux
    port map (
            O => \N__46137\,
            I => \N__46134\
        );

    \I__10799\ : LocalMux
    port map (
            O => \N__46134\,
            I => n11_adj_758
        );

    \I__10798\ : InMux
    port map (
            O => \N__46131\,
            I => n10562
        );

    \I__10797\ : InMux
    port map (
            O => \N__46128\,
            I => \N__46125\
        );

    \I__10796\ : LocalMux
    port map (
            O => \N__46125\,
            I => n10_adj_757
        );

    \I__10795\ : InMux
    port map (
            O => \N__46122\,
            I => \bfn_15_28_0_\
        );

    \I__10794\ : InMux
    port map (
            O => \N__46119\,
            I => \N__46116\
        );

    \I__10793\ : LocalMux
    port map (
            O => \N__46116\,
            I => n26
        );

    \I__10792\ : InMux
    port map (
            O => \N__46113\,
            I => \bfn_15_26_0_\
        );

    \I__10791\ : InMux
    port map (
            O => \N__46110\,
            I => \N__46107\
        );

    \I__10790\ : LocalMux
    port map (
            O => \N__46107\,
            I => n25
        );

    \I__10789\ : InMux
    port map (
            O => \N__46104\,
            I => n10548
        );

    \I__10788\ : InMux
    port map (
            O => \N__46101\,
            I => \N__46098\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__46098\,
            I => n24
        );

    \I__10786\ : InMux
    port map (
            O => \N__46095\,
            I => n10549
        );

    \I__10785\ : InMux
    port map (
            O => \N__46092\,
            I => \N__46089\
        );

    \I__10784\ : LocalMux
    port map (
            O => \N__46089\,
            I => n23
        );

    \I__10783\ : InMux
    port map (
            O => \N__46086\,
            I => n10550
        );

    \I__10782\ : InMux
    port map (
            O => \N__46083\,
            I => \N__46080\
        );

    \I__10781\ : LocalMux
    port map (
            O => \N__46080\,
            I => n22
        );

    \I__10780\ : InMux
    port map (
            O => \N__46077\,
            I => n10551
        );

    \I__10779\ : InMux
    port map (
            O => \N__46074\,
            I => \N__46071\
        );

    \I__10778\ : LocalMux
    port map (
            O => \N__46071\,
            I => n21_adj_737
        );

    \I__10777\ : InMux
    port map (
            O => \N__46068\,
            I => n10552
        );

    \I__10776\ : InMux
    port map (
            O => \N__46065\,
            I => \N__46062\
        );

    \I__10775\ : LocalMux
    port map (
            O => \N__46062\,
            I => n20
        );

    \I__10774\ : InMux
    port map (
            O => \N__46059\,
            I => n10553
        );

    \I__10773\ : InMux
    port map (
            O => \N__46056\,
            I => \N__46053\
        );

    \I__10772\ : LocalMux
    port map (
            O => \N__46053\,
            I => n19_adj_718
        );

    \I__10771\ : InMux
    port map (
            O => \N__46050\,
            I => n10554
        );

    \I__10770\ : InMux
    port map (
            O => \N__46047\,
            I => \N__46043\
        );

    \I__10769\ : CascadeMux
    port map (
            O => \N__46046\,
            I => \N__46040\
        );

    \I__10768\ : LocalMux
    port map (
            O => \N__46043\,
            I => \N__46036\
        );

    \I__10767\ : InMux
    port map (
            O => \N__46040\,
            I => \N__46033\
        );

    \I__10766\ : InMux
    port map (
            O => \N__46039\,
            I => \N__46030\
        );

    \I__10765\ : Odrv4
    port map (
            O => \N__46036\,
            I => \nx.n2298\
        );

    \I__10764\ : LocalMux
    port map (
            O => \N__46033\,
            I => \nx.n2298\
        );

    \I__10763\ : LocalMux
    port map (
            O => \N__46030\,
            I => \nx.n2298\
        );

    \I__10762\ : CascadeMux
    port map (
            O => \N__46023\,
            I => \N__46020\
        );

    \I__10761\ : InMux
    port map (
            O => \N__46020\,
            I => \N__46017\
        );

    \I__10760\ : LocalMux
    port map (
            O => \N__46017\,
            I => \N__46014\
        );

    \I__10759\ : Odrv4
    port map (
            O => \N__46014\,
            I => \nx.n2365\
        );

    \I__10758\ : InMux
    port map (
            O => \N__46011\,
            I => \nx.n10719\
        );

    \I__10757\ : CascadeMux
    port map (
            O => \N__46008\,
            I => \N__46004\
        );

    \I__10756\ : CascadeMux
    port map (
            O => \N__46007\,
            I => \N__46001\
        );

    \I__10755\ : InMux
    port map (
            O => \N__46004\,
            I => \N__45998\
        );

    \I__10754\ : InMux
    port map (
            O => \N__46001\,
            I => \N__45995\
        );

    \I__10753\ : LocalMux
    port map (
            O => \N__45998\,
            I => \nx.n2297\
        );

    \I__10752\ : LocalMux
    port map (
            O => \N__45995\,
            I => \nx.n2297\
        );

    \I__10751\ : InMux
    port map (
            O => \N__45990\,
            I => \N__45987\
        );

    \I__10750\ : LocalMux
    port map (
            O => \N__45987\,
            I => \nx.n2364\
        );

    \I__10749\ : InMux
    port map (
            O => \N__45984\,
            I => \nx.n10720\
        );

    \I__10748\ : CascadeMux
    port map (
            O => \N__45981\,
            I => \N__45978\
        );

    \I__10747\ : InMux
    port map (
            O => \N__45978\,
            I => \N__45975\
        );

    \I__10746\ : LocalMux
    port map (
            O => \N__45975\,
            I => \N__45972\
        );

    \I__10745\ : Span4Mux_v
    port map (
            O => \N__45972\,
            I => \N__45968\
        );

    \I__10744\ : InMux
    port map (
            O => \N__45971\,
            I => \N__45965\
        );

    \I__10743\ : Odrv4
    port map (
            O => \N__45968\,
            I => \nx.n2296\
        );

    \I__10742\ : LocalMux
    port map (
            O => \N__45965\,
            I => \nx.n2296\
        );

    \I__10741\ : InMux
    port map (
            O => \N__45960\,
            I => \N__45957\
        );

    \I__10740\ : LocalMux
    port map (
            O => \N__45957\,
            I => \N__45954\
        );

    \I__10739\ : Span4Mux_h
    port map (
            O => \N__45954\,
            I => \N__45951\
        );

    \I__10738\ : Odrv4
    port map (
            O => \N__45951\,
            I => \nx.n2363\
        );

    \I__10737\ : InMux
    port map (
            O => \N__45948\,
            I => \nx.n10721\
        );

    \I__10736\ : CascadeMux
    port map (
            O => \N__45945\,
            I => \N__45942\
        );

    \I__10735\ : InMux
    port map (
            O => \N__45942\,
            I => \N__45939\
        );

    \I__10734\ : LocalMux
    port map (
            O => \N__45939\,
            I => \N__45935\
        );

    \I__10733\ : InMux
    port map (
            O => \N__45938\,
            I => \N__45931\
        );

    \I__10732\ : Span4Mux_h
    port map (
            O => \N__45935\,
            I => \N__45928\
        );

    \I__10731\ : InMux
    port map (
            O => \N__45934\,
            I => \N__45925\
        );

    \I__10730\ : LocalMux
    port map (
            O => \N__45931\,
            I => \nx.n2295\
        );

    \I__10729\ : Odrv4
    port map (
            O => \N__45928\,
            I => \nx.n2295\
        );

    \I__10728\ : LocalMux
    port map (
            O => \N__45925\,
            I => \nx.n2295\
        );

    \I__10727\ : CascadeMux
    port map (
            O => \N__45918\,
            I => \N__45915\
        );

    \I__10726\ : InMux
    port map (
            O => \N__45915\,
            I => \N__45912\
        );

    \I__10725\ : LocalMux
    port map (
            O => \N__45912\,
            I => \N__45909\
        );

    \I__10724\ : Span4Mux_h
    port map (
            O => \N__45909\,
            I => \N__45906\
        );

    \I__10723\ : Span4Mux_h
    port map (
            O => \N__45906\,
            I => \N__45903\
        );

    \I__10722\ : Odrv4
    port map (
            O => \N__45903\,
            I => \nx.n2362\
        );

    \I__10721\ : InMux
    port map (
            O => \N__45900\,
            I => \nx.n10722\
        );

    \I__10720\ : CascadeMux
    port map (
            O => \N__45897\,
            I => \N__45894\
        );

    \I__10719\ : InMux
    port map (
            O => \N__45894\,
            I => \N__45891\
        );

    \I__10718\ : LocalMux
    port map (
            O => \N__45891\,
            I => \N__45887\
        );

    \I__10717\ : InMux
    port map (
            O => \N__45890\,
            I => \N__45883\
        );

    \I__10716\ : Span4Mux_h
    port map (
            O => \N__45887\,
            I => \N__45880\
        );

    \I__10715\ : InMux
    port map (
            O => \N__45886\,
            I => \N__45877\
        );

    \I__10714\ : LocalMux
    port map (
            O => \N__45883\,
            I => \nx.n2294\
        );

    \I__10713\ : Odrv4
    port map (
            O => \N__45880\,
            I => \nx.n2294\
        );

    \I__10712\ : LocalMux
    port map (
            O => \N__45877\,
            I => \nx.n2294\
        );

    \I__10711\ : InMux
    port map (
            O => \N__45870\,
            I => \N__45867\
        );

    \I__10710\ : LocalMux
    port map (
            O => \N__45867\,
            I => \N__45864\
        );

    \I__10709\ : Span4Mux_h
    port map (
            O => \N__45864\,
            I => \N__45861\
        );

    \I__10708\ : Span4Mux_h
    port map (
            O => \N__45861\,
            I => \N__45858\
        );

    \I__10707\ : Odrv4
    port map (
            O => \N__45858\,
            I => \nx.n2361\
        );

    \I__10706\ : InMux
    port map (
            O => \N__45855\,
            I => \bfn_15_25_0_\
        );

    \I__10705\ : CascadeMux
    port map (
            O => \N__45852\,
            I => \N__45849\
        );

    \I__10704\ : InMux
    port map (
            O => \N__45849\,
            I => \N__45845\
        );

    \I__10703\ : CascadeMux
    port map (
            O => \N__45848\,
            I => \N__45842\
        );

    \I__10702\ : LocalMux
    port map (
            O => \N__45845\,
            I => \N__45839\
        );

    \I__10701\ : InMux
    port map (
            O => \N__45842\,
            I => \N__45836\
        );

    \I__10700\ : Span4Mux_h
    port map (
            O => \N__45839\,
            I => \N__45833\
        );

    \I__10699\ : LocalMux
    port map (
            O => \N__45836\,
            I => \nx.n2293\
        );

    \I__10698\ : Odrv4
    port map (
            O => \N__45833\,
            I => \nx.n2293\
        );

    \I__10697\ : InMux
    port map (
            O => \N__45828\,
            I => \N__45825\
        );

    \I__10696\ : LocalMux
    port map (
            O => \N__45825\,
            I => \N__45822\
        );

    \I__10695\ : Span4Mux_h
    port map (
            O => \N__45822\,
            I => \N__45819\
        );

    \I__10694\ : Span4Mux_h
    port map (
            O => \N__45819\,
            I => \N__45816\
        );

    \I__10693\ : Odrv4
    port map (
            O => \N__45816\,
            I => \nx.n2360\
        );

    \I__10692\ : InMux
    port map (
            O => \N__45813\,
            I => \nx.n10724\
        );

    \I__10691\ : CascadeMux
    port map (
            O => \N__45810\,
            I => \N__45807\
        );

    \I__10690\ : InMux
    port map (
            O => \N__45807\,
            I => \N__45802\
        );

    \I__10689\ : CascadeMux
    port map (
            O => \N__45806\,
            I => \N__45799\
        );

    \I__10688\ : CascadeMux
    port map (
            O => \N__45805\,
            I => \N__45796\
        );

    \I__10687\ : LocalMux
    port map (
            O => \N__45802\,
            I => \N__45793\
        );

    \I__10686\ : InMux
    port map (
            O => \N__45799\,
            I => \N__45790\
        );

    \I__10685\ : InMux
    port map (
            O => \N__45796\,
            I => \N__45787\
        );

    \I__10684\ : Span4Mux_h
    port map (
            O => \N__45793\,
            I => \N__45784\
        );

    \I__10683\ : LocalMux
    port map (
            O => \N__45790\,
            I => \nx.n2292\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__45787\,
            I => \nx.n2292\
        );

    \I__10681\ : Odrv4
    port map (
            O => \N__45784\,
            I => \nx.n2292\
        );

    \I__10680\ : InMux
    port map (
            O => \N__45777\,
            I => \N__45774\
        );

    \I__10679\ : LocalMux
    port map (
            O => \N__45774\,
            I => \N__45771\
        );

    \I__10678\ : Odrv4
    port map (
            O => \N__45771\,
            I => \nx.n2359\
        );

    \I__10677\ : InMux
    port map (
            O => \N__45768\,
            I => \nx.n10725\
        );

    \I__10676\ : CascadeMux
    port map (
            O => \N__45765\,
            I => \N__45734\
        );

    \I__10675\ : CascadeMux
    port map (
            O => \N__45764\,
            I => \N__45724\
        );

    \I__10674\ : CascadeMux
    port map (
            O => \N__45763\,
            I => \N__45721\
        );

    \I__10673\ : CascadeMux
    port map (
            O => \N__45762\,
            I => \N__45717\
        );

    \I__10672\ : CascadeMux
    port map (
            O => \N__45761\,
            I => \N__45714\
        );

    \I__10671\ : CascadeMux
    port map (
            O => \N__45760\,
            I => \N__45711\
        );

    \I__10670\ : CascadeMux
    port map (
            O => \N__45759\,
            I => \N__45708\
        );

    \I__10669\ : CascadeMux
    port map (
            O => \N__45758\,
            I => \N__45705\
        );

    \I__10668\ : InMux
    port map (
            O => \N__45757\,
            I => \N__45701\
        );

    \I__10667\ : CascadeMux
    port map (
            O => \N__45756\,
            I => \N__45681\
        );

    \I__10666\ : CascadeMux
    port map (
            O => \N__45755\,
            I => \N__45673\
        );

    \I__10665\ : CascadeMux
    port map (
            O => \N__45754\,
            I => \N__45667\
        );

    \I__10664\ : CascadeMux
    port map (
            O => \N__45753\,
            I => \N__45662\
        );

    \I__10663\ : CascadeMux
    port map (
            O => \N__45752\,
            I => \N__45651\
        );

    \I__10662\ : CascadeMux
    port map (
            O => \N__45751\,
            I => \N__45639\
        );

    \I__10661\ : CascadeMux
    port map (
            O => \N__45750\,
            I => \N__45636\
        );

    \I__10660\ : InMux
    port map (
            O => \N__45749\,
            I => \N__45616\
        );

    \I__10659\ : InMux
    port map (
            O => \N__45748\,
            I => \N__45616\
        );

    \I__10658\ : InMux
    port map (
            O => \N__45747\,
            I => \N__45616\
        );

    \I__10657\ : InMux
    port map (
            O => \N__45746\,
            I => \N__45616\
        );

    \I__10656\ : InMux
    port map (
            O => \N__45745\,
            I => \N__45607\
        );

    \I__10655\ : InMux
    port map (
            O => \N__45744\,
            I => \N__45607\
        );

    \I__10654\ : InMux
    port map (
            O => \N__45743\,
            I => \N__45607\
        );

    \I__10653\ : InMux
    port map (
            O => \N__45742\,
            I => \N__45607\
        );

    \I__10652\ : InMux
    port map (
            O => \N__45741\,
            I => \N__45600\
        );

    \I__10651\ : InMux
    port map (
            O => \N__45740\,
            I => \N__45600\
        );

    \I__10650\ : InMux
    port map (
            O => \N__45739\,
            I => \N__45600\
        );

    \I__10649\ : InMux
    port map (
            O => \N__45738\,
            I => \N__45591\
        );

    \I__10648\ : InMux
    port map (
            O => \N__45737\,
            I => \N__45591\
        );

    \I__10647\ : InMux
    port map (
            O => \N__45734\,
            I => \N__45591\
        );

    \I__10646\ : InMux
    port map (
            O => \N__45733\,
            I => \N__45591\
        );

    \I__10645\ : CascadeMux
    port map (
            O => \N__45732\,
            I => \N__45581\
        );

    \I__10644\ : CascadeMux
    port map (
            O => \N__45731\,
            I => \N__45573\
        );

    \I__10643\ : CascadeMux
    port map (
            O => \N__45730\,
            I => \N__45559\
        );

    \I__10642\ : CascadeMux
    port map (
            O => \N__45729\,
            I => \N__45544\
        );

    \I__10641\ : CascadeMux
    port map (
            O => \N__45728\,
            I => \N__45536\
        );

    \I__10640\ : CascadeMux
    port map (
            O => \N__45727\,
            I => \N__45527\
        );

    \I__10639\ : InMux
    port map (
            O => \N__45724\,
            I => \N__45514\
        );

    \I__10638\ : InMux
    port map (
            O => \N__45721\,
            I => \N__45514\
        );

    \I__10637\ : InMux
    port map (
            O => \N__45720\,
            I => \N__45514\
        );

    \I__10636\ : InMux
    port map (
            O => \N__45717\,
            I => \N__45514\
        );

    \I__10635\ : InMux
    port map (
            O => \N__45714\,
            I => \N__45514\
        );

    \I__10634\ : InMux
    port map (
            O => \N__45711\,
            I => \N__45507\
        );

    \I__10633\ : InMux
    port map (
            O => \N__45708\,
            I => \N__45507\
        );

    \I__10632\ : InMux
    port map (
            O => \N__45705\,
            I => \N__45507\
        );

    \I__10631\ : CascadeMux
    port map (
            O => \N__45704\,
            I => \N__45498\
        );

    \I__10630\ : LocalMux
    port map (
            O => \N__45701\,
            I => \N__45493\
        );

    \I__10629\ : InMux
    port map (
            O => \N__45700\,
            I => \N__45486\
        );

    \I__10628\ : InMux
    port map (
            O => \N__45699\,
            I => \N__45486\
        );

    \I__10627\ : InMux
    port map (
            O => \N__45698\,
            I => \N__45486\
        );

    \I__10626\ : InMux
    port map (
            O => \N__45697\,
            I => \N__45479\
        );

    \I__10625\ : InMux
    port map (
            O => \N__45696\,
            I => \N__45479\
        );

    \I__10624\ : InMux
    port map (
            O => \N__45695\,
            I => \N__45479\
        );

    \I__10623\ : InMux
    port map (
            O => \N__45694\,
            I => \N__45470\
        );

    \I__10622\ : InMux
    port map (
            O => \N__45693\,
            I => \N__45470\
        );

    \I__10621\ : InMux
    port map (
            O => \N__45692\,
            I => \N__45470\
        );

    \I__10620\ : InMux
    port map (
            O => \N__45691\,
            I => \N__45470\
        );

    \I__10619\ : InMux
    port map (
            O => \N__45690\,
            I => \N__45463\
        );

    \I__10618\ : InMux
    port map (
            O => \N__45689\,
            I => \N__45463\
        );

    \I__10617\ : InMux
    port map (
            O => \N__45688\,
            I => \N__45463\
        );

    \I__10616\ : InMux
    port map (
            O => \N__45687\,
            I => \N__45456\
        );

    \I__10615\ : InMux
    port map (
            O => \N__45686\,
            I => \N__45456\
        );

    \I__10614\ : InMux
    port map (
            O => \N__45685\,
            I => \N__45456\
        );

    \I__10613\ : InMux
    port map (
            O => \N__45684\,
            I => \N__45423\
        );

    \I__10612\ : InMux
    port map (
            O => \N__45681\,
            I => \N__45423\
        );

    \I__10611\ : InMux
    port map (
            O => \N__45680\,
            I => \N__45423\
        );

    \I__10610\ : InMux
    port map (
            O => \N__45679\,
            I => \N__45423\
        );

    \I__10609\ : InMux
    port map (
            O => \N__45678\,
            I => \N__45418\
        );

    \I__10608\ : InMux
    port map (
            O => \N__45677\,
            I => \N__45418\
        );

    \I__10607\ : InMux
    port map (
            O => \N__45676\,
            I => \N__45402\
        );

    \I__10606\ : InMux
    port map (
            O => \N__45673\,
            I => \N__45402\
        );

    \I__10605\ : InMux
    port map (
            O => \N__45672\,
            I => \N__45402\
        );

    \I__10604\ : InMux
    port map (
            O => \N__45671\,
            I => \N__45402\
        );

    \I__10603\ : CascadeMux
    port map (
            O => \N__45670\,
            I => \N__45396\
        );

    \I__10602\ : InMux
    port map (
            O => \N__45667\,
            I => \N__45386\
        );

    \I__10601\ : InMux
    port map (
            O => \N__45666\,
            I => \N__45386\
        );

    \I__10600\ : InMux
    port map (
            O => \N__45665\,
            I => \N__45375\
        );

    \I__10599\ : InMux
    port map (
            O => \N__45662\,
            I => \N__45375\
        );

    \I__10598\ : InMux
    port map (
            O => \N__45661\,
            I => \N__45375\
        );

    \I__10597\ : InMux
    port map (
            O => \N__45660\,
            I => \N__45375\
        );

    \I__10596\ : InMux
    port map (
            O => \N__45659\,
            I => \N__45375\
        );

    \I__10595\ : InMux
    port map (
            O => \N__45658\,
            I => \N__45368\
        );

    \I__10594\ : InMux
    port map (
            O => \N__45657\,
            I => \N__45368\
        );

    \I__10593\ : InMux
    port map (
            O => \N__45656\,
            I => \N__45368\
        );

    \I__10592\ : InMux
    port map (
            O => \N__45655\,
            I => \N__45357\
        );

    \I__10591\ : InMux
    port map (
            O => \N__45654\,
            I => \N__45357\
        );

    \I__10590\ : InMux
    port map (
            O => \N__45651\,
            I => \N__45357\
        );

    \I__10589\ : InMux
    port map (
            O => \N__45650\,
            I => \N__45357\
        );

    \I__10588\ : InMux
    port map (
            O => \N__45649\,
            I => \N__45357\
        );

    \I__10587\ : InMux
    port map (
            O => \N__45648\,
            I => \N__45348\
        );

    \I__10586\ : InMux
    port map (
            O => \N__45647\,
            I => \N__45348\
        );

    \I__10585\ : InMux
    port map (
            O => \N__45646\,
            I => \N__45348\
        );

    \I__10584\ : InMux
    port map (
            O => \N__45645\,
            I => \N__45348\
        );

    \I__10583\ : InMux
    port map (
            O => \N__45644\,
            I => \N__45339\
        );

    \I__10582\ : InMux
    port map (
            O => \N__45643\,
            I => \N__45339\
        );

    \I__10581\ : InMux
    port map (
            O => \N__45642\,
            I => \N__45339\
        );

    \I__10580\ : InMux
    port map (
            O => \N__45639\,
            I => \N__45339\
        );

    \I__10579\ : InMux
    port map (
            O => \N__45636\,
            I => \N__45333\
        );

    \I__10578\ : InMux
    port map (
            O => \N__45635\,
            I => \N__45333\
        );

    \I__10577\ : InMux
    port map (
            O => \N__45634\,
            I => \N__45326\
        );

    \I__10576\ : InMux
    port map (
            O => \N__45633\,
            I => \N__45326\
        );

    \I__10575\ : InMux
    port map (
            O => \N__45632\,
            I => \N__45326\
        );

    \I__10574\ : CascadeMux
    port map (
            O => \N__45631\,
            I => \N__45319\
        );

    \I__10573\ : CascadeMux
    port map (
            O => \N__45630\,
            I => \N__45314\
        );

    \I__10572\ : CascadeMux
    port map (
            O => \N__45629\,
            I => \N__45304\
        );

    \I__10571\ : CascadeMux
    port map (
            O => \N__45628\,
            I => \N__45299\
        );

    \I__10570\ : CascadeMux
    port map (
            O => \N__45627\,
            I => \N__45293\
        );

    \I__10569\ : CascadeMux
    port map (
            O => \N__45626\,
            I => \N__45289\
        );

    \I__10568\ : CascadeMux
    port map (
            O => \N__45625\,
            I => \N__45286\
        );

    \I__10567\ : LocalMux
    port map (
            O => \N__45616\,
            I => \N__45276\
        );

    \I__10566\ : LocalMux
    port map (
            O => \N__45607\,
            I => \N__45269\
        );

    \I__10565\ : LocalMux
    port map (
            O => \N__45600\,
            I => \N__45269\
        );

    \I__10564\ : LocalMux
    port map (
            O => \N__45591\,
            I => \N__45269\
        );

    \I__10563\ : InMux
    port map (
            O => \N__45590\,
            I => \N__45262\
        );

    \I__10562\ : InMux
    port map (
            O => \N__45589\,
            I => \N__45262\
        );

    \I__10561\ : InMux
    port map (
            O => \N__45588\,
            I => \N__45262\
        );

    \I__10560\ : InMux
    port map (
            O => \N__45587\,
            I => \N__45251\
        );

    \I__10559\ : InMux
    port map (
            O => \N__45586\,
            I => \N__45251\
        );

    \I__10558\ : InMux
    port map (
            O => \N__45585\,
            I => \N__45251\
        );

    \I__10557\ : InMux
    port map (
            O => \N__45584\,
            I => \N__45251\
        );

    \I__10556\ : InMux
    port map (
            O => \N__45581\,
            I => \N__45251\
        );

    \I__10555\ : InMux
    port map (
            O => \N__45580\,
            I => \N__45244\
        );

    \I__10554\ : InMux
    port map (
            O => \N__45579\,
            I => \N__45244\
        );

    \I__10553\ : InMux
    port map (
            O => \N__45578\,
            I => \N__45244\
        );

    \I__10552\ : InMux
    port map (
            O => \N__45577\,
            I => \N__45239\
        );

    \I__10551\ : InMux
    port map (
            O => \N__45576\,
            I => \N__45239\
        );

    \I__10550\ : InMux
    port map (
            O => \N__45573\,
            I => \N__45232\
        );

    \I__10549\ : InMux
    port map (
            O => \N__45572\,
            I => \N__45232\
        );

    \I__10548\ : InMux
    port map (
            O => \N__45571\,
            I => \N__45232\
        );

    \I__10547\ : CascadeMux
    port map (
            O => \N__45570\,
            I => \N__45228\
        );

    \I__10546\ : CascadeMux
    port map (
            O => \N__45569\,
            I => \N__45224\
        );

    \I__10545\ : CascadeMux
    port map (
            O => \N__45568\,
            I => \N__45220\
        );

    \I__10544\ : InMux
    port map (
            O => \N__45567\,
            I => \N__45211\
        );

    \I__10543\ : InMux
    port map (
            O => \N__45566\,
            I => \N__45211\
        );

    \I__10542\ : InMux
    port map (
            O => \N__45565\,
            I => \N__45211\
        );

    \I__10541\ : InMux
    port map (
            O => \N__45564\,
            I => \N__45206\
        );

    \I__10540\ : InMux
    port map (
            O => \N__45563\,
            I => \N__45206\
        );

    \I__10539\ : InMux
    port map (
            O => \N__45562\,
            I => \N__45197\
        );

    \I__10538\ : InMux
    port map (
            O => \N__45559\,
            I => \N__45197\
        );

    \I__10537\ : InMux
    port map (
            O => \N__45558\,
            I => \N__45197\
        );

    \I__10536\ : InMux
    port map (
            O => \N__45557\,
            I => \N__45197\
        );

    \I__10535\ : InMux
    port map (
            O => \N__45556\,
            I => \N__45190\
        );

    \I__10534\ : InMux
    port map (
            O => \N__45555\,
            I => \N__45190\
        );

    \I__10533\ : InMux
    port map (
            O => \N__45554\,
            I => \N__45190\
        );

    \I__10532\ : InMux
    port map (
            O => \N__45553\,
            I => \N__45183\
        );

    \I__10531\ : InMux
    port map (
            O => \N__45552\,
            I => \N__45183\
        );

    \I__10530\ : InMux
    port map (
            O => \N__45551\,
            I => \N__45183\
        );

    \I__10529\ : InMux
    port map (
            O => \N__45550\,
            I => \N__45174\
        );

    \I__10528\ : InMux
    port map (
            O => \N__45549\,
            I => \N__45174\
        );

    \I__10527\ : InMux
    port map (
            O => \N__45548\,
            I => \N__45174\
        );

    \I__10526\ : InMux
    port map (
            O => \N__45547\,
            I => \N__45174\
        );

    \I__10525\ : InMux
    port map (
            O => \N__45544\,
            I => \N__45163\
        );

    \I__10524\ : InMux
    port map (
            O => \N__45543\,
            I => \N__45163\
        );

    \I__10523\ : InMux
    port map (
            O => \N__45542\,
            I => \N__45163\
        );

    \I__10522\ : InMux
    port map (
            O => \N__45541\,
            I => \N__45163\
        );

    \I__10521\ : InMux
    port map (
            O => \N__45540\,
            I => \N__45163\
        );

    \I__10520\ : InMux
    port map (
            O => \N__45539\,
            I => \N__45152\
        );

    \I__10519\ : InMux
    port map (
            O => \N__45536\,
            I => \N__45152\
        );

    \I__10518\ : InMux
    port map (
            O => \N__45535\,
            I => \N__45152\
        );

    \I__10517\ : InMux
    port map (
            O => \N__45534\,
            I => \N__45152\
        );

    \I__10516\ : InMux
    port map (
            O => \N__45533\,
            I => \N__45152\
        );

    \I__10515\ : InMux
    port map (
            O => \N__45532\,
            I => \N__45145\
        );

    \I__10514\ : InMux
    port map (
            O => \N__45531\,
            I => \N__45145\
        );

    \I__10513\ : InMux
    port map (
            O => \N__45530\,
            I => \N__45145\
        );

    \I__10512\ : InMux
    port map (
            O => \N__45527\,
            I => \N__45142\
        );

    \I__10511\ : InMux
    port map (
            O => \N__45526\,
            I => \N__45131\
        );

    \I__10510\ : InMux
    port map (
            O => \N__45525\,
            I => \N__45128\
        );

    \I__10509\ : LocalMux
    port map (
            O => \N__45514\,
            I => \N__45123\
        );

    \I__10508\ : LocalMux
    port map (
            O => \N__45507\,
            I => \N__45123\
        );

    \I__10507\ : InMux
    port map (
            O => \N__45506\,
            I => \N__45116\
        );

    \I__10506\ : InMux
    port map (
            O => \N__45505\,
            I => \N__45116\
        );

    \I__10505\ : InMux
    port map (
            O => \N__45504\,
            I => \N__45116\
        );

    \I__10504\ : InMux
    port map (
            O => \N__45503\,
            I => \N__45105\
        );

    \I__10503\ : InMux
    port map (
            O => \N__45502\,
            I => \N__45105\
        );

    \I__10502\ : InMux
    port map (
            O => \N__45501\,
            I => \N__45105\
        );

    \I__10501\ : InMux
    port map (
            O => \N__45498\,
            I => \N__45105\
        );

    \I__10500\ : InMux
    port map (
            O => \N__45497\,
            I => \N__45105\
        );

    \I__10499\ : CascadeMux
    port map (
            O => \N__45496\,
            I => \N__45101\
        );

    \I__10498\ : Span4Mux_v
    port map (
            O => \N__45493\,
            I => \N__45087\
        );

    \I__10497\ : LocalMux
    port map (
            O => \N__45486\,
            I => \N__45082\
        );

    \I__10496\ : LocalMux
    port map (
            O => \N__45479\,
            I => \N__45082\
        );

    \I__10495\ : LocalMux
    port map (
            O => \N__45470\,
            I => \N__45079\
        );

    \I__10494\ : LocalMux
    port map (
            O => \N__45463\,
            I => \N__45074\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__45456\,
            I => \N__45074\
        );

    \I__10492\ : InMux
    port map (
            O => \N__45455\,
            I => \N__45067\
        );

    \I__10491\ : InMux
    port map (
            O => \N__45454\,
            I => \N__45067\
        );

    \I__10490\ : InMux
    port map (
            O => \N__45453\,
            I => \N__45067\
        );

    \I__10489\ : InMux
    port map (
            O => \N__45452\,
            I => \N__45060\
        );

    \I__10488\ : InMux
    port map (
            O => \N__45451\,
            I => \N__45060\
        );

    \I__10487\ : InMux
    port map (
            O => \N__45450\,
            I => \N__45060\
        );

    \I__10486\ : InMux
    port map (
            O => \N__45449\,
            I => \N__45053\
        );

    \I__10485\ : InMux
    port map (
            O => \N__45448\,
            I => \N__45053\
        );

    \I__10484\ : InMux
    port map (
            O => \N__45447\,
            I => \N__45053\
        );

    \I__10483\ : InMux
    port map (
            O => \N__45446\,
            I => \N__45046\
        );

    \I__10482\ : InMux
    port map (
            O => \N__45445\,
            I => \N__45046\
        );

    \I__10481\ : InMux
    port map (
            O => \N__45444\,
            I => \N__45046\
        );

    \I__10480\ : InMux
    port map (
            O => \N__45443\,
            I => \N__45037\
        );

    \I__10479\ : InMux
    port map (
            O => \N__45442\,
            I => \N__45037\
        );

    \I__10478\ : InMux
    port map (
            O => \N__45441\,
            I => \N__45037\
        );

    \I__10477\ : InMux
    port map (
            O => \N__45440\,
            I => \N__45037\
        );

    \I__10476\ : CascadeMux
    port map (
            O => \N__45439\,
            I => \N__45033\
        );

    \I__10475\ : CascadeMux
    port map (
            O => \N__45438\,
            I => \N__45030\
        );

    \I__10474\ : CascadeMux
    port map (
            O => \N__45437\,
            I => \N__45020\
        );

    \I__10473\ : InMux
    port map (
            O => \N__45436\,
            I => \N__45007\
        );

    \I__10472\ : InMux
    port map (
            O => \N__45435\,
            I => \N__45007\
        );

    \I__10471\ : InMux
    port map (
            O => \N__45434\,
            I => \N__45007\
        );

    \I__10470\ : InMux
    port map (
            O => \N__45433\,
            I => \N__45007\
        );

    \I__10469\ : InMux
    port map (
            O => \N__45432\,
            I => \N__45004\
        );

    \I__10468\ : LocalMux
    port map (
            O => \N__45423\,
            I => \N__44999\
        );

    \I__10467\ : LocalMux
    port map (
            O => \N__45418\,
            I => \N__44999\
        );

    \I__10466\ : InMux
    port map (
            O => \N__45417\,
            I => \N__44990\
        );

    \I__10465\ : InMux
    port map (
            O => \N__45416\,
            I => \N__44990\
        );

    \I__10464\ : InMux
    port map (
            O => \N__45415\,
            I => \N__44990\
        );

    \I__10463\ : InMux
    port map (
            O => \N__45414\,
            I => \N__44990\
        );

    \I__10462\ : InMux
    port map (
            O => \N__45413\,
            I => \N__44983\
        );

    \I__10461\ : InMux
    port map (
            O => \N__45412\,
            I => \N__44983\
        );

    \I__10460\ : InMux
    port map (
            O => \N__45411\,
            I => \N__44983\
        );

    \I__10459\ : LocalMux
    port map (
            O => \N__45402\,
            I => \N__44980\
        );

    \I__10458\ : InMux
    port map (
            O => \N__45401\,
            I => \N__44973\
        );

    \I__10457\ : InMux
    port map (
            O => \N__45400\,
            I => \N__44973\
        );

    \I__10456\ : InMux
    port map (
            O => \N__45399\,
            I => \N__44973\
        );

    \I__10455\ : InMux
    port map (
            O => \N__45396\,
            I => \N__44962\
        );

    \I__10454\ : InMux
    port map (
            O => \N__45395\,
            I => \N__44962\
        );

    \I__10453\ : InMux
    port map (
            O => \N__45394\,
            I => \N__44962\
        );

    \I__10452\ : InMux
    port map (
            O => \N__45393\,
            I => \N__44962\
        );

    \I__10451\ : InMux
    port map (
            O => \N__45392\,
            I => \N__44962\
        );

    \I__10450\ : CascadeMux
    port map (
            O => \N__45391\,
            I => \N__44959\
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__45386\,
            I => \N__44950\
        );

    \I__10448\ : LocalMux
    port map (
            O => \N__45375\,
            I => \N__44950\
        );

    \I__10447\ : LocalMux
    port map (
            O => \N__45368\,
            I => \N__44941\
        );

    \I__10446\ : LocalMux
    port map (
            O => \N__45357\,
            I => \N__44941\
        );

    \I__10445\ : LocalMux
    port map (
            O => \N__45348\,
            I => \N__44941\
        );

    \I__10444\ : LocalMux
    port map (
            O => \N__45339\,
            I => \N__44941\
        );

    \I__10443\ : InMux
    port map (
            O => \N__45338\,
            I => \N__44938\
        );

    \I__10442\ : LocalMux
    port map (
            O => \N__45333\,
            I => \N__44918\
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__45326\,
            I => \N__44918\
        );

    \I__10440\ : InMux
    port map (
            O => \N__45325\,
            I => \N__44907\
        );

    \I__10439\ : InMux
    port map (
            O => \N__45324\,
            I => \N__44907\
        );

    \I__10438\ : InMux
    port map (
            O => \N__45323\,
            I => \N__44907\
        );

    \I__10437\ : InMux
    port map (
            O => \N__45322\,
            I => \N__44907\
        );

    \I__10436\ : InMux
    port map (
            O => \N__45319\,
            I => \N__44907\
        );

    \I__10435\ : InMux
    port map (
            O => \N__45318\,
            I => \N__44900\
        );

    \I__10434\ : InMux
    port map (
            O => \N__45317\,
            I => \N__44900\
        );

    \I__10433\ : InMux
    port map (
            O => \N__45314\,
            I => \N__44900\
        );

    \I__10432\ : InMux
    port map (
            O => \N__45313\,
            I => \N__44893\
        );

    \I__10431\ : InMux
    port map (
            O => \N__45312\,
            I => \N__44893\
        );

    \I__10430\ : InMux
    port map (
            O => \N__45311\,
            I => \N__44893\
        );

    \I__10429\ : InMux
    port map (
            O => \N__45310\,
            I => \N__44886\
        );

    \I__10428\ : InMux
    port map (
            O => \N__45309\,
            I => \N__44886\
        );

    \I__10427\ : InMux
    port map (
            O => \N__45308\,
            I => \N__44886\
        );

    \I__10426\ : InMux
    port map (
            O => \N__45307\,
            I => \N__44879\
        );

    \I__10425\ : InMux
    port map (
            O => \N__45304\,
            I => \N__44879\
        );

    \I__10424\ : InMux
    port map (
            O => \N__45303\,
            I => \N__44879\
        );

    \I__10423\ : InMux
    port map (
            O => \N__45302\,
            I => \N__44872\
        );

    \I__10422\ : InMux
    port map (
            O => \N__45299\,
            I => \N__44872\
        );

    \I__10421\ : InMux
    port map (
            O => \N__45298\,
            I => \N__44872\
        );

    \I__10420\ : InMux
    port map (
            O => \N__45297\,
            I => \N__44864\
        );

    \I__10419\ : InMux
    port map (
            O => \N__45296\,
            I => \N__44864\
        );

    \I__10418\ : InMux
    port map (
            O => \N__45293\,
            I => \N__44856\
        );

    \I__10417\ : InMux
    port map (
            O => \N__45292\,
            I => \N__44849\
        );

    \I__10416\ : InMux
    port map (
            O => \N__45289\,
            I => \N__44849\
        );

    \I__10415\ : InMux
    port map (
            O => \N__45286\,
            I => \N__44849\
        );

    \I__10414\ : InMux
    port map (
            O => \N__45285\,
            I => \N__44844\
        );

    \I__10413\ : InMux
    port map (
            O => \N__45284\,
            I => \N__44844\
        );

    \I__10412\ : InMux
    port map (
            O => \N__45283\,
            I => \N__44835\
        );

    \I__10411\ : InMux
    port map (
            O => \N__45282\,
            I => \N__44835\
        );

    \I__10410\ : InMux
    port map (
            O => \N__45281\,
            I => \N__44835\
        );

    \I__10409\ : InMux
    port map (
            O => \N__45280\,
            I => \N__44835\
        );

    \I__10408\ : CascadeMux
    port map (
            O => \N__45279\,
            I => \N__44829\
        );

    \I__10407\ : Span4Mux_v
    port map (
            O => \N__45276\,
            I => \N__44823\
        );

    \I__10406\ : Span4Mux_v
    port map (
            O => \N__45269\,
            I => \N__44823\
        );

    \I__10405\ : LocalMux
    port map (
            O => \N__45262\,
            I => \N__44812\
        );

    \I__10404\ : LocalMux
    port map (
            O => \N__45251\,
            I => \N__44812\
        );

    \I__10403\ : LocalMux
    port map (
            O => \N__45244\,
            I => \N__44812\
        );

    \I__10402\ : LocalMux
    port map (
            O => \N__45239\,
            I => \N__44812\
        );

    \I__10401\ : LocalMux
    port map (
            O => \N__45232\,
            I => \N__44812\
        );

    \I__10400\ : InMux
    port map (
            O => \N__45231\,
            I => \N__44805\
        );

    \I__10399\ : InMux
    port map (
            O => \N__45228\,
            I => \N__44805\
        );

    \I__10398\ : InMux
    port map (
            O => \N__45227\,
            I => \N__44805\
        );

    \I__10397\ : InMux
    port map (
            O => \N__45224\,
            I => \N__44794\
        );

    \I__10396\ : InMux
    port map (
            O => \N__45223\,
            I => \N__44794\
        );

    \I__10395\ : InMux
    port map (
            O => \N__45220\,
            I => \N__44794\
        );

    \I__10394\ : InMux
    port map (
            O => \N__45219\,
            I => \N__44794\
        );

    \I__10393\ : InMux
    port map (
            O => \N__45218\,
            I => \N__44794\
        );

    \I__10392\ : LocalMux
    port map (
            O => \N__45211\,
            I => \N__44791\
        );

    \I__10391\ : LocalMux
    port map (
            O => \N__45206\,
            I => \N__44774\
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__45197\,
            I => \N__44774\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__45190\,
            I => \N__44774\
        );

    \I__10388\ : LocalMux
    port map (
            O => \N__45183\,
            I => \N__44774\
        );

    \I__10387\ : LocalMux
    port map (
            O => \N__45174\,
            I => \N__44774\
        );

    \I__10386\ : LocalMux
    port map (
            O => \N__45163\,
            I => \N__44774\
        );

    \I__10385\ : LocalMux
    port map (
            O => \N__45152\,
            I => \N__44774\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__45145\,
            I => \N__44774\
        );

    \I__10383\ : LocalMux
    port map (
            O => \N__45142\,
            I => \N__44771\
        );

    \I__10382\ : InMux
    port map (
            O => \N__45141\,
            I => \N__44762\
        );

    \I__10381\ : InMux
    port map (
            O => \N__45140\,
            I => \N__44762\
        );

    \I__10380\ : InMux
    port map (
            O => \N__45139\,
            I => \N__44762\
        );

    \I__10379\ : InMux
    port map (
            O => \N__45138\,
            I => \N__44762\
        );

    \I__10378\ : InMux
    port map (
            O => \N__45137\,
            I => \N__44753\
        );

    \I__10377\ : InMux
    port map (
            O => \N__45136\,
            I => \N__44753\
        );

    \I__10376\ : InMux
    port map (
            O => \N__45135\,
            I => \N__44753\
        );

    \I__10375\ : InMux
    port map (
            O => \N__45134\,
            I => \N__44753\
        );

    \I__10374\ : LocalMux
    port map (
            O => \N__45131\,
            I => \N__44748\
        );

    \I__10373\ : LocalMux
    port map (
            O => \N__45128\,
            I => \N__44748\
        );

    \I__10372\ : Span4Mux_s1_h
    port map (
            O => \N__45123\,
            I => \N__44743\
        );

    \I__10371\ : LocalMux
    port map (
            O => \N__45116\,
            I => \N__44743\
        );

    \I__10370\ : LocalMux
    port map (
            O => \N__45105\,
            I => \N__44740\
        );

    \I__10369\ : InMux
    port map (
            O => \N__45104\,
            I => \N__44737\
        );

    \I__10368\ : InMux
    port map (
            O => \N__45101\,
            I => \N__44730\
        );

    \I__10367\ : InMux
    port map (
            O => \N__45100\,
            I => \N__44730\
        );

    \I__10366\ : InMux
    port map (
            O => \N__45099\,
            I => \N__44730\
        );

    \I__10365\ : InMux
    port map (
            O => \N__45098\,
            I => \N__44723\
        );

    \I__10364\ : InMux
    port map (
            O => \N__45097\,
            I => \N__44723\
        );

    \I__10363\ : InMux
    port map (
            O => \N__45096\,
            I => \N__44723\
        );

    \I__10362\ : CascadeMux
    port map (
            O => \N__45095\,
            I => \N__44719\
        );

    \I__10361\ : CascadeMux
    port map (
            O => \N__45094\,
            I => \N__44711\
        );

    \I__10360\ : CascadeMux
    port map (
            O => \N__45093\,
            I => \N__44707\
        );

    \I__10359\ : InMux
    port map (
            O => \N__45092\,
            I => \N__44699\
        );

    \I__10358\ : InMux
    port map (
            O => \N__45091\,
            I => \N__44699\
        );

    \I__10357\ : InMux
    port map (
            O => \N__45090\,
            I => \N__44699\
        );

    \I__10356\ : Span4Mux_h
    port map (
            O => \N__45087\,
            I => \N__44692\
        );

    \I__10355\ : Span4Mux_v
    port map (
            O => \N__45082\,
            I => \N__44692\
        );

    \I__10354\ : Span4Mux_h
    port map (
            O => \N__45079\,
            I => \N__44692\
        );

    \I__10353\ : Span4Mux_h
    port map (
            O => \N__45074\,
            I => \N__44685\
        );

    \I__10352\ : LocalMux
    port map (
            O => \N__45067\,
            I => \N__44685\
        );

    \I__10351\ : LocalMux
    port map (
            O => \N__45060\,
            I => \N__44685\
        );

    \I__10350\ : LocalMux
    port map (
            O => \N__45053\,
            I => \N__44678\
        );

    \I__10349\ : LocalMux
    port map (
            O => \N__45046\,
            I => \N__44678\
        );

    \I__10348\ : LocalMux
    port map (
            O => \N__45037\,
            I => \N__44678\
        );

    \I__10347\ : InMux
    port map (
            O => \N__45036\,
            I => \N__44671\
        );

    \I__10346\ : InMux
    port map (
            O => \N__45033\,
            I => \N__44671\
        );

    \I__10345\ : InMux
    port map (
            O => \N__45030\,
            I => \N__44671\
        );

    \I__10344\ : CascadeMux
    port map (
            O => \N__45029\,
            I => \N__44667\
        );

    \I__10343\ : InMux
    port map (
            O => \N__45028\,
            I => \N__44656\
        );

    \I__10342\ : InMux
    port map (
            O => \N__45027\,
            I => \N__44656\
        );

    \I__10341\ : InMux
    port map (
            O => \N__45026\,
            I => \N__44656\
        );

    \I__10340\ : InMux
    port map (
            O => \N__45025\,
            I => \N__44656\
        );

    \I__10339\ : InMux
    port map (
            O => \N__45024\,
            I => \N__44649\
        );

    \I__10338\ : InMux
    port map (
            O => \N__45023\,
            I => \N__44649\
        );

    \I__10337\ : InMux
    port map (
            O => \N__45020\,
            I => \N__44649\
        );

    \I__10336\ : CascadeMux
    port map (
            O => \N__45019\,
            I => \N__44646\
        );

    \I__10335\ : InMux
    port map (
            O => \N__45018\,
            I => \N__44637\
        );

    \I__10334\ : InMux
    port map (
            O => \N__45017\,
            I => \N__44637\
        );

    \I__10333\ : InMux
    port map (
            O => \N__45016\,
            I => \N__44637\
        );

    \I__10332\ : LocalMux
    port map (
            O => \N__45007\,
            I => \N__44625\
        );

    \I__10331\ : LocalMux
    port map (
            O => \N__45004\,
            I => \N__44625\
        );

    \I__10330\ : Span4Mux_h
    port map (
            O => \N__44999\,
            I => \N__44618\
        );

    \I__10329\ : LocalMux
    port map (
            O => \N__44990\,
            I => \N__44618\
        );

    \I__10328\ : LocalMux
    port map (
            O => \N__44983\,
            I => \N__44618\
        );

    \I__10327\ : Span4Mux_s2_h
    port map (
            O => \N__44980\,
            I => \N__44611\
        );

    \I__10326\ : LocalMux
    port map (
            O => \N__44973\,
            I => \N__44611\
        );

    \I__10325\ : LocalMux
    port map (
            O => \N__44962\,
            I => \N__44611\
        );

    \I__10324\ : InMux
    port map (
            O => \N__44959\,
            I => \N__44602\
        );

    \I__10323\ : InMux
    port map (
            O => \N__44958\,
            I => \N__44602\
        );

    \I__10322\ : InMux
    port map (
            O => \N__44957\,
            I => \N__44602\
        );

    \I__10321\ : InMux
    port map (
            O => \N__44956\,
            I => \N__44602\
        );

    \I__10320\ : CascadeMux
    port map (
            O => \N__44955\,
            I => \N__44597\
        );

    \I__10319\ : Span4Mux_h
    port map (
            O => \N__44950\,
            I => \N__44589\
        );

    \I__10318\ : Span4Mux_v
    port map (
            O => \N__44941\,
            I => \N__44589\
        );

    \I__10317\ : LocalMux
    port map (
            O => \N__44938\,
            I => \N__44589\
        );

    \I__10316\ : InMux
    port map (
            O => \N__44937\,
            I => \N__44582\
        );

    \I__10315\ : InMux
    port map (
            O => \N__44936\,
            I => \N__44582\
        );

    \I__10314\ : InMux
    port map (
            O => \N__44935\,
            I => \N__44582\
        );

    \I__10313\ : InMux
    port map (
            O => \N__44934\,
            I => \N__44575\
        );

    \I__10312\ : InMux
    port map (
            O => \N__44933\,
            I => \N__44575\
        );

    \I__10311\ : InMux
    port map (
            O => \N__44932\,
            I => \N__44575\
        );

    \I__10310\ : InMux
    port map (
            O => \N__44931\,
            I => \N__44568\
        );

    \I__10309\ : InMux
    port map (
            O => \N__44930\,
            I => \N__44568\
        );

    \I__10308\ : InMux
    port map (
            O => \N__44929\,
            I => \N__44568\
        );

    \I__10307\ : InMux
    port map (
            O => \N__44928\,
            I => \N__44561\
        );

    \I__10306\ : InMux
    port map (
            O => \N__44927\,
            I => \N__44561\
        );

    \I__10305\ : InMux
    port map (
            O => \N__44926\,
            I => \N__44561\
        );

    \I__10304\ : InMux
    port map (
            O => \N__44925\,
            I => \N__44554\
        );

    \I__10303\ : InMux
    port map (
            O => \N__44924\,
            I => \N__44554\
        );

    \I__10302\ : InMux
    port map (
            O => \N__44923\,
            I => \N__44554\
        );

    \I__10301\ : Span4Mux_v
    port map (
            O => \N__44918\,
            I => \N__44547\
        );

    \I__10300\ : LocalMux
    port map (
            O => \N__44907\,
            I => \N__44547\
        );

    \I__10299\ : LocalMux
    port map (
            O => \N__44900\,
            I => \N__44547\
        );

    \I__10298\ : LocalMux
    port map (
            O => \N__44893\,
            I => \N__44538\
        );

    \I__10297\ : LocalMux
    port map (
            O => \N__44886\,
            I => \N__44538\
        );

    \I__10296\ : LocalMux
    port map (
            O => \N__44879\,
            I => \N__44538\
        );

    \I__10295\ : LocalMux
    port map (
            O => \N__44872\,
            I => \N__44538\
        );

    \I__10294\ : InMux
    port map (
            O => \N__44871\,
            I => \N__44531\
        );

    \I__10293\ : InMux
    port map (
            O => \N__44870\,
            I => \N__44531\
        );

    \I__10292\ : InMux
    port map (
            O => \N__44869\,
            I => \N__44531\
        );

    \I__10291\ : LocalMux
    port map (
            O => \N__44864\,
            I => \N__44528\
        );

    \I__10290\ : InMux
    port map (
            O => \N__44863\,
            I => \N__44523\
        );

    \I__10289\ : InMux
    port map (
            O => \N__44862\,
            I => \N__44523\
        );

    \I__10288\ : InMux
    port map (
            O => \N__44861\,
            I => \N__44513\
        );

    \I__10287\ : InMux
    port map (
            O => \N__44860\,
            I => \N__44513\
        );

    \I__10286\ : InMux
    port map (
            O => \N__44859\,
            I => \N__44510\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__44856\,
            I => \N__44507\
        );

    \I__10284\ : LocalMux
    port map (
            O => \N__44849\,
            I => \N__44500\
        );

    \I__10283\ : LocalMux
    port map (
            O => \N__44844\,
            I => \N__44500\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__44835\,
            I => \N__44500\
        );

    \I__10281\ : InMux
    port map (
            O => \N__44834\,
            I => \N__44495\
        );

    \I__10280\ : InMux
    port map (
            O => \N__44833\,
            I => \N__44495\
        );

    \I__10279\ : InMux
    port map (
            O => \N__44832\,
            I => \N__44492\
        );

    \I__10278\ : InMux
    port map (
            O => \N__44829\,
            I => \N__44487\
        );

    \I__10277\ : InMux
    port map (
            O => \N__44828\,
            I => \N__44487\
        );

    \I__10276\ : Span4Mux_v
    port map (
            O => \N__44823\,
            I => \N__44474\
        );

    \I__10275\ : Span4Mux_v
    port map (
            O => \N__44812\,
            I => \N__44474\
        );

    \I__10274\ : LocalMux
    port map (
            O => \N__44805\,
            I => \N__44474\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__44794\,
            I => \N__44474\
        );

    \I__10272\ : Span4Mux_h
    port map (
            O => \N__44791\,
            I => \N__44463\
        );

    \I__10271\ : Span4Mux_v
    port map (
            O => \N__44774\,
            I => \N__44463\
        );

    \I__10270\ : Span4Mux_v
    port map (
            O => \N__44771\,
            I => \N__44463\
        );

    \I__10269\ : LocalMux
    port map (
            O => \N__44762\,
            I => \N__44463\
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__44753\,
            I => \N__44463\
        );

    \I__10267\ : Span4Mux_v
    port map (
            O => \N__44748\,
            I => \N__44450\
        );

    \I__10266\ : Span4Mux_h
    port map (
            O => \N__44743\,
            I => \N__44450\
        );

    \I__10265\ : Span4Mux_v
    port map (
            O => \N__44740\,
            I => \N__44450\
        );

    \I__10264\ : LocalMux
    port map (
            O => \N__44737\,
            I => \N__44450\
        );

    \I__10263\ : LocalMux
    port map (
            O => \N__44730\,
            I => \N__44450\
        );

    \I__10262\ : LocalMux
    port map (
            O => \N__44723\,
            I => \N__44450\
        );

    \I__10261\ : InMux
    port map (
            O => \N__44722\,
            I => \N__44441\
        );

    \I__10260\ : InMux
    port map (
            O => \N__44719\,
            I => \N__44441\
        );

    \I__10259\ : InMux
    port map (
            O => \N__44718\,
            I => \N__44441\
        );

    \I__10258\ : InMux
    port map (
            O => \N__44717\,
            I => \N__44441\
        );

    \I__10257\ : CascadeMux
    port map (
            O => \N__44716\,
            I => \N__44437\
        );

    \I__10256\ : InMux
    port map (
            O => \N__44715\,
            I => \N__44426\
        );

    \I__10255\ : InMux
    port map (
            O => \N__44714\,
            I => \N__44426\
        );

    \I__10254\ : InMux
    port map (
            O => \N__44711\,
            I => \N__44426\
        );

    \I__10253\ : InMux
    port map (
            O => \N__44710\,
            I => \N__44419\
        );

    \I__10252\ : InMux
    port map (
            O => \N__44707\,
            I => \N__44419\
        );

    \I__10251\ : InMux
    port map (
            O => \N__44706\,
            I => \N__44419\
        );

    \I__10250\ : LocalMux
    port map (
            O => \N__44699\,
            I => \N__44416\
        );

    \I__10249\ : Span4Mux_h
    port map (
            O => \N__44692\,
            I => \N__44407\
        );

    \I__10248\ : Span4Mux_v
    port map (
            O => \N__44685\,
            I => \N__44407\
        );

    \I__10247\ : Span4Mux_h
    port map (
            O => \N__44678\,
            I => \N__44407\
        );

    \I__10246\ : LocalMux
    port map (
            O => \N__44671\,
            I => \N__44407\
        );

    \I__10245\ : InMux
    port map (
            O => \N__44670\,
            I => \N__44398\
        );

    \I__10244\ : InMux
    port map (
            O => \N__44667\,
            I => \N__44398\
        );

    \I__10243\ : InMux
    port map (
            O => \N__44666\,
            I => \N__44398\
        );

    \I__10242\ : InMux
    port map (
            O => \N__44665\,
            I => \N__44398\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__44656\,
            I => \N__44393\
        );

    \I__10240\ : LocalMux
    port map (
            O => \N__44649\,
            I => \N__44393\
        );

    \I__10239\ : InMux
    port map (
            O => \N__44646\,
            I => \N__44386\
        );

    \I__10238\ : InMux
    port map (
            O => \N__44645\,
            I => \N__44386\
        );

    \I__10237\ : InMux
    port map (
            O => \N__44644\,
            I => \N__44386\
        );

    \I__10236\ : LocalMux
    port map (
            O => \N__44637\,
            I => \N__44382\
        );

    \I__10235\ : InMux
    port map (
            O => \N__44636\,
            I => \N__44375\
        );

    \I__10234\ : InMux
    port map (
            O => \N__44635\,
            I => \N__44375\
        );

    \I__10233\ : InMux
    port map (
            O => \N__44634\,
            I => \N__44375\
        );

    \I__10232\ : InMux
    port map (
            O => \N__44633\,
            I => \N__44368\
        );

    \I__10231\ : InMux
    port map (
            O => \N__44632\,
            I => \N__44368\
        );

    \I__10230\ : InMux
    port map (
            O => \N__44631\,
            I => \N__44368\
        );

    \I__10229\ : InMux
    port map (
            O => \N__44630\,
            I => \N__44365\
        );

    \I__10228\ : Span4Mux_v
    port map (
            O => \N__44625\,
            I => \N__44360\
        );

    \I__10227\ : Span4Mux_v
    port map (
            O => \N__44618\,
            I => \N__44360\
        );

    \I__10226\ : Span4Mux_h
    port map (
            O => \N__44611\,
            I => \N__44355\
        );

    \I__10225\ : LocalMux
    port map (
            O => \N__44602\,
            I => \N__44355\
        );

    \I__10224\ : InMux
    port map (
            O => \N__44601\,
            I => \N__44346\
        );

    \I__10223\ : InMux
    port map (
            O => \N__44600\,
            I => \N__44346\
        );

    \I__10222\ : InMux
    port map (
            O => \N__44597\,
            I => \N__44346\
        );

    \I__10221\ : InMux
    port map (
            O => \N__44596\,
            I => \N__44346\
        );

    \I__10220\ : Span4Mux_v
    port map (
            O => \N__44589\,
            I => \N__44339\
        );

    \I__10219\ : LocalMux
    port map (
            O => \N__44582\,
            I => \N__44339\
        );

    \I__10218\ : LocalMux
    port map (
            O => \N__44575\,
            I => \N__44339\
        );

    \I__10217\ : LocalMux
    port map (
            O => \N__44568\,
            I => \N__44332\
        );

    \I__10216\ : LocalMux
    port map (
            O => \N__44561\,
            I => \N__44332\
        );

    \I__10215\ : LocalMux
    port map (
            O => \N__44554\,
            I => \N__44332\
        );

    \I__10214\ : Span4Mux_v
    port map (
            O => \N__44547\,
            I => \N__44325\
        );

    \I__10213\ : Span4Mux_s2_h
    port map (
            O => \N__44538\,
            I => \N__44325\
        );

    \I__10212\ : LocalMux
    port map (
            O => \N__44531\,
            I => \N__44325\
        );

    \I__10211\ : Span4Mux_h
    port map (
            O => \N__44528\,
            I => \N__44320\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__44523\,
            I => \N__44320\
        );

    \I__10209\ : InMux
    port map (
            O => \N__44522\,
            I => \N__44313\
        );

    \I__10208\ : InMux
    port map (
            O => \N__44521\,
            I => \N__44313\
        );

    \I__10207\ : InMux
    port map (
            O => \N__44520\,
            I => \N__44313\
        );

    \I__10206\ : InMux
    port map (
            O => \N__44519\,
            I => \N__44308\
        );

    \I__10205\ : InMux
    port map (
            O => \N__44518\,
            I => \N__44308\
        );

    \I__10204\ : LocalMux
    port map (
            O => \N__44513\,
            I => \N__44305\
        );

    \I__10203\ : LocalMux
    port map (
            O => \N__44510\,
            I => \N__44302\
        );

    \I__10202\ : Span4Mux_v
    port map (
            O => \N__44507\,
            I => \N__44291\
        );

    \I__10201\ : Span4Mux_v
    port map (
            O => \N__44500\,
            I => \N__44291\
        );

    \I__10200\ : LocalMux
    port map (
            O => \N__44495\,
            I => \N__44291\
        );

    \I__10199\ : LocalMux
    port map (
            O => \N__44492\,
            I => \N__44291\
        );

    \I__10198\ : LocalMux
    port map (
            O => \N__44487\,
            I => \N__44291\
        );

    \I__10197\ : InMux
    port map (
            O => \N__44486\,
            I => \N__44288\
        );

    \I__10196\ : InMux
    port map (
            O => \N__44485\,
            I => \N__44281\
        );

    \I__10195\ : InMux
    port map (
            O => \N__44484\,
            I => \N__44281\
        );

    \I__10194\ : InMux
    port map (
            O => \N__44483\,
            I => \N__44281\
        );

    \I__10193\ : Span4Mux_h
    port map (
            O => \N__44474\,
            I => \N__44272\
        );

    \I__10192\ : Span4Mux_h
    port map (
            O => \N__44463\,
            I => \N__44272\
        );

    \I__10191\ : Span4Mux_h
    port map (
            O => \N__44450\,
            I => \N__44272\
        );

    \I__10190\ : LocalMux
    port map (
            O => \N__44441\,
            I => \N__44272\
        );

    \I__10189\ : InMux
    port map (
            O => \N__44440\,
            I => \N__44265\
        );

    \I__10188\ : InMux
    port map (
            O => \N__44437\,
            I => \N__44265\
        );

    \I__10187\ : InMux
    port map (
            O => \N__44436\,
            I => \N__44265\
        );

    \I__10186\ : InMux
    port map (
            O => \N__44435\,
            I => \N__44258\
        );

    \I__10185\ : InMux
    port map (
            O => \N__44434\,
            I => \N__44258\
        );

    \I__10184\ : InMux
    port map (
            O => \N__44433\,
            I => \N__44258\
        );

    \I__10183\ : LocalMux
    port map (
            O => \N__44426\,
            I => \N__44251\
        );

    \I__10182\ : LocalMux
    port map (
            O => \N__44419\,
            I => \N__44251\
        );

    \I__10181\ : Sp12to4
    port map (
            O => \N__44416\,
            I => \N__44251\
        );

    \I__10180\ : Span4Mux_v
    port map (
            O => \N__44407\,
            I => \N__44248\
        );

    \I__10179\ : LocalMux
    port map (
            O => \N__44398\,
            I => \N__44245\
        );

    \I__10178\ : Sp12to4
    port map (
            O => \N__44393\,
            I => \N__44240\
        );

    \I__10177\ : LocalMux
    port map (
            O => \N__44386\,
            I => \N__44240\
        );

    \I__10176\ : InMux
    port map (
            O => \N__44385\,
            I => \N__44237\
        );

    \I__10175\ : Span12Mux_s8_h
    port map (
            O => \N__44382\,
            I => \N__44228\
        );

    \I__10174\ : LocalMux
    port map (
            O => \N__44375\,
            I => \N__44228\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__44368\,
            I => \N__44228\
        );

    \I__10172\ : LocalMux
    port map (
            O => \N__44365\,
            I => \N__44228\
        );

    \I__10171\ : Span4Mux_h
    port map (
            O => \N__44360\,
            I => \N__44221\
        );

    \I__10170\ : Span4Mux_h
    port map (
            O => \N__44355\,
            I => \N__44221\
        );

    \I__10169\ : LocalMux
    port map (
            O => \N__44346\,
            I => \N__44221\
        );

    \I__10168\ : Span4Mux_v
    port map (
            O => \N__44339\,
            I => \N__44208\
        );

    \I__10167\ : Span4Mux_h
    port map (
            O => \N__44332\,
            I => \N__44208\
        );

    \I__10166\ : Span4Mux_h
    port map (
            O => \N__44325\,
            I => \N__44208\
        );

    \I__10165\ : Span4Mux_v
    port map (
            O => \N__44320\,
            I => \N__44208\
        );

    \I__10164\ : LocalMux
    port map (
            O => \N__44313\,
            I => \N__44208\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__44308\,
            I => \N__44208\
        );

    \I__10162\ : Span4Mux_v
    port map (
            O => \N__44305\,
            I => \N__44203\
        );

    \I__10161\ : Span4Mux_v
    port map (
            O => \N__44302\,
            I => \N__44203\
        );

    \I__10160\ : Span4Mux_h
    port map (
            O => \N__44291\,
            I => \N__44196\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__44288\,
            I => \N__44196\
        );

    \I__10158\ : LocalMux
    port map (
            O => \N__44281\,
            I => \N__44196\
        );

    \I__10157\ : Span4Mux_v
    port map (
            O => \N__44272\,
            I => \N__44189\
        );

    \I__10156\ : LocalMux
    port map (
            O => \N__44265\,
            I => \N__44189\
        );

    \I__10155\ : LocalMux
    port map (
            O => \N__44258\,
            I => \N__44189\
        );

    \I__10154\ : Span12Mux_s10_h
    port map (
            O => \N__44251\,
            I => \N__44186\
        );

    \I__10153\ : Span4Mux_v
    port map (
            O => \N__44248\,
            I => \N__44183\
        );

    \I__10152\ : Span12Mux_v
    port map (
            O => \N__44245\,
            I => \N__44176\
        );

    \I__10151\ : Span12Mux_v
    port map (
            O => \N__44240\,
            I => \N__44176\
        );

    \I__10150\ : LocalMux
    port map (
            O => \N__44237\,
            I => \N__44176\
        );

    \I__10149\ : Span12Mux_v
    port map (
            O => \N__44228\,
            I => \N__44173\
        );

    \I__10148\ : Span4Mux_v
    port map (
            O => \N__44221\,
            I => \N__44168\
        );

    \I__10147\ : Span4Mux_h
    port map (
            O => \N__44208\,
            I => \N__44168\
        );

    \I__10146\ : Span4Mux_v
    port map (
            O => \N__44203\,
            I => \N__44161\
        );

    \I__10145\ : Span4Mux_h
    port map (
            O => \N__44196\,
            I => \N__44161\
        );

    \I__10144\ : Span4Mux_v
    port map (
            O => \N__44189\,
            I => \N__44161\
        );

    \I__10143\ : Odrv12
    port map (
            O => \N__44186\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10142\ : Odrv4
    port map (
            O => \N__44183\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10141\ : Odrv12
    port map (
            O => \N__44176\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10140\ : Odrv12
    port map (
            O => \N__44173\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10139\ : Odrv4
    port map (
            O => \N__44168\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10138\ : Odrv4
    port map (
            O => \N__44161\,
            I => \CONSTANT_ONE_NET\
        );

    \I__10137\ : InMux
    port map (
            O => \N__44148\,
            I => \N__44144\
        );

    \I__10136\ : InMux
    port map (
            O => \N__44147\,
            I => \N__44141\
        );

    \I__10135\ : LocalMux
    port map (
            O => \N__44144\,
            I => \N__44138\
        );

    \I__10134\ : LocalMux
    port map (
            O => \N__44141\,
            I => \N__44135\
        );

    \I__10133\ : Odrv4
    port map (
            O => \N__44138\,
            I => \nx.n2291\
        );

    \I__10132\ : Odrv4
    port map (
            O => \N__44135\,
            I => \nx.n2291\
        );

    \I__10131\ : CascadeMux
    port map (
            O => \N__44130\,
            I => \N__44124\
        );

    \I__10130\ : CascadeMux
    port map (
            O => \N__44129\,
            I => \N__44119\
        );

    \I__10129\ : CascadeMux
    port map (
            O => \N__44128\,
            I => \N__44110\
        );

    \I__10128\ : InMux
    port map (
            O => \N__44127\,
            I => \N__44106\
        );

    \I__10127\ : InMux
    port map (
            O => \N__44124\,
            I => \N__44103\
        );

    \I__10126\ : CascadeMux
    port map (
            O => \N__44123\,
            I => \N__44100\
        );

    \I__10125\ : InMux
    port map (
            O => \N__44122\,
            I => \N__44091\
        );

    \I__10124\ : InMux
    port map (
            O => \N__44119\,
            I => \N__44091\
        );

    \I__10123\ : InMux
    port map (
            O => \N__44118\,
            I => \N__44091\
        );

    \I__10122\ : CascadeMux
    port map (
            O => \N__44117\,
            I => \N__44087\
        );

    \I__10121\ : CascadeMux
    port map (
            O => \N__44116\,
            I => \N__44083\
        );

    \I__10120\ : InMux
    port map (
            O => \N__44115\,
            I => \N__44070\
        );

    \I__10119\ : InMux
    port map (
            O => \N__44114\,
            I => \N__44070\
        );

    \I__10118\ : InMux
    port map (
            O => \N__44113\,
            I => \N__44070\
        );

    \I__10117\ : InMux
    port map (
            O => \N__44110\,
            I => \N__44070\
        );

    \I__10116\ : InMux
    port map (
            O => \N__44109\,
            I => \N__44070\
        );

    \I__10115\ : LocalMux
    port map (
            O => \N__44106\,
            I => \N__44067\
        );

    \I__10114\ : LocalMux
    port map (
            O => \N__44103\,
            I => \N__44064\
        );

    \I__10113\ : InMux
    port map (
            O => \N__44100\,
            I => \N__44061\
        );

    \I__10112\ : InMux
    port map (
            O => \N__44099\,
            I => \N__44058\
        );

    \I__10111\ : InMux
    port map (
            O => \N__44098\,
            I => \N__44055\
        );

    \I__10110\ : LocalMux
    port map (
            O => \N__44091\,
            I => \N__44052\
        );

    \I__10109\ : InMux
    port map (
            O => \N__44090\,
            I => \N__44045\
        );

    \I__10108\ : InMux
    port map (
            O => \N__44087\,
            I => \N__44045\
        );

    \I__10107\ : InMux
    port map (
            O => \N__44086\,
            I => \N__44045\
        );

    \I__10106\ : InMux
    port map (
            O => \N__44083\,
            I => \N__44038\
        );

    \I__10105\ : InMux
    port map (
            O => \N__44082\,
            I => \N__44038\
        );

    \I__10104\ : InMux
    port map (
            O => \N__44081\,
            I => \N__44038\
        );

    \I__10103\ : LocalMux
    port map (
            O => \N__44070\,
            I => \N__44035\
        );

    \I__10102\ : Span4Mux_h
    port map (
            O => \N__44067\,
            I => \N__44026\
        );

    \I__10101\ : Span4Mux_h
    port map (
            O => \N__44064\,
            I => \N__44026\
        );

    \I__10100\ : LocalMux
    port map (
            O => \N__44061\,
            I => \N__44026\
        );

    \I__10099\ : LocalMux
    port map (
            O => \N__44058\,
            I => \N__44026\
        );

    \I__10098\ : LocalMux
    port map (
            O => \N__44055\,
            I => \nx.n2324\
        );

    \I__10097\ : Odrv4
    port map (
            O => \N__44052\,
            I => \nx.n2324\
        );

    \I__10096\ : LocalMux
    port map (
            O => \N__44045\,
            I => \nx.n2324\
        );

    \I__10095\ : LocalMux
    port map (
            O => \N__44038\,
            I => \nx.n2324\
        );

    \I__10094\ : Odrv4
    port map (
            O => \N__44035\,
            I => \nx.n2324\
        );

    \I__10093\ : Odrv4
    port map (
            O => \N__44026\,
            I => \nx.n2324\
        );

    \I__10092\ : InMux
    port map (
            O => \N__44013\,
            I => \nx.n10726\
        );

    \I__10091\ : InMux
    port map (
            O => \N__44010\,
            I => \N__44007\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__44007\,
            I => \N__44003\
        );

    \I__10089\ : InMux
    port map (
            O => \N__44006\,
            I => \N__44000\
        );

    \I__10088\ : Span4Mux_h
    port map (
            O => \N__44003\,
            I => \N__43997\
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__44000\,
            I => \N__43992\
        );

    \I__10086\ : Span4Mux_h
    port map (
            O => \N__43997\,
            I => \N__43992\
        );

    \I__10085\ : Odrv4
    port map (
            O => \N__43992\,
            I => \nx.n2390\
        );

    \I__10084\ : InMux
    port map (
            O => \N__43989\,
            I => \nx.n10711\
        );

    \I__10083\ : CascadeMux
    port map (
            O => \N__43986\,
            I => \N__43982\
        );

    \I__10082\ : CascadeMux
    port map (
            O => \N__43985\,
            I => \N__43979\
        );

    \I__10081\ : InMux
    port map (
            O => \N__43982\,
            I => \N__43976\
        );

    \I__10080\ : InMux
    port map (
            O => \N__43979\,
            I => \N__43972\
        );

    \I__10079\ : LocalMux
    port map (
            O => \N__43976\,
            I => \N__43969\
        );

    \I__10078\ : InMux
    port map (
            O => \N__43975\,
            I => \N__43966\
        );

    \I__10077\ : LocalMux
    port map (
            O => \N__43972\,
            I => \N__43963\
        );

    \I__10076\ : Odrv4
    port map (
            O => \N__43969\,
            I => \nx.n2305\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__43966\,
            I => \nx.n2305\
        );

    \I__10074\ : Odrv4
    port map (
            O => \N__43963\,
            I => \nx.n2305\
        );

    \I__10073\ : InMux
    port map (
            O => \N__43956\,
            I => \N__43953\
        );

    \I__10072\ : LocalMux
    port map (
            O => \N__43953\,
            I => \N__43950\
        );

    \I__10071\ : Span4Mux_h
    port map (
            O => \N__43950\,
            I => \N__43947\
        );

    \I__10070\ : Odrv4
    port map (
            O => \N__43947\,
            I => \nx.n2372\
        );

    \I__10069\ : InMux
    port map (
            O => \N__43944\,
            I => \nx.n10712\
        );

    \I__10068\ : InMux
    port map (
            O => \N__43941\,
            I => \N__43937\
        );

    \I__10067\ : InMux
    port map (
            O => \N__43940\,
            I => \N__43933\
        );

    \I__10066\ : LocalMux
    port map (
            O => \N__43937\,
            I => \N__43930\
        );

    \I__10065\ : InMux
    port map (
            O => \N__43936\,
            I => \N__43927\
        );

    \I__10064\ : LocalMux
    port map (
            O => \N__43933\,
            I => \N__43924\
        );

    \I__10063\ : Odrv4
    port map (
            O => \N__43930\,
            I => \nx.n2304\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__43927\,
            I => \nx.n2304\
        );

    \I__10061\ : Odrv12
    port map (
            O => \N__43924\,
            I => \nx.n2304\
        );

    \I__10060\ : CascadeMux
    port map (
            O => \N__43917\,
            I => \N__43914\
        );

    \I__10059\ : InMux
    port map (
            O => \N__43914\,
            I => \N__43911\
        );

    \I__10058\ : LocalMux
    port map (
            O => \N__43911\,
            I => \N__43908\
        );

    \I__10057\ : Span4Mux_h
    port map (
            O => \N__43908\,
            I => \N__43905\
        );

    \I__10056\ : Odrv4
    port map (
            O => \N__43905\,
            I => \nx.n2371\
        );

    \I__10055\ : InMux
    port map (
            O => \N__43902\,
            I => \nx.n10713\
        );

    \I__10054\ : InMux
    port map (
            O => \N__43899\,
            I => \N__43895\
        );

    \I__10053\ : CascadeMux
    port map (
            O => \N__43898\,
            I => \N__43891\
        );

    \I__10052\ : LocalMux
    port map (
            O => \N__43895\,
            I => \N__43888\
        );

    \I__10051\ : InMux
    port map (
            O => \N__43894\,
            I => \N__43885\
        );

    \I__10050\ : InMux
    port map (
            O => \N__43891\,
            I => \N__43882\
        );

    \I__10049\ : Span4Mux_h
    port map (
            O => \N__43888\,
            I => \N__43879\
        );

    \I__10048\ : LocalMux
    port map (
            O => \N__43885\,
            I => \nx.n2303\
        );

    \I__10047\ : LocalMux
    port map (
            O => \N__43882\,
            I => \nx.n2303\
        );

    \I__10046\ : Odrv4
    port map (
            O => \N__43879\,
            I => \nx.n2303\
        );

    \I__10045\ : CascadeMux
    port map (
            O => \N__43872\,
            I => \N__43869\
        );

    \I__10044\ : InMux
    port map (
            O => \N__43869\,
            I => \N__43866\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__43866\,
            I => \nx.n2370\
        );

    \I__10042\ : InMux
    port map (
            O => \N__43863\,
            I => \nx.n10714\
        );

    \I__10041\ : CascadeMux
    port map (
            O => \N__43860\,
            I => \N__43857\
        );

    \I__10040\ : InMux
    port map (
            O => \N__43857\,
            I => \N__43854\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__43854\,
            I => \N__43849\
        );

    \I__10038\ : InMux
    port map (
            O => \N__43853\,
            I => \N__43846\
        );

    \I__10037\ : InMux
    port map (
            O => \N__43852\,
            I => \N__43843\
        );

    \I__10036\ : Span4Mux_v
    port map (
            O => \N__43849\,
            I => \N__43840\
        );

    \I__10035\ : LocalMux
    port map (
            O => \N__43846\,
            I => \nx.n2302\
        );

    \I__10034\ : LocalMux
    port map (
            O => \N__43843\,
            I => \nx.n2302\
        );

    \I__10033\ : Odrv4
    port map (
            O => \N__43840\,
            I => \nx.n2302\
        );

    \I__10032\ : CascadeMux
    port map (
            O => \N__43833\,
            I => \N__43830\
        );

    \I__10031\ : InMux
    port map (
            O => \N__43830\,
            I => \N__43827\
        );

    \I__10030\ : LocalMux
    port map (
            O => \N__43827\,
            I => \N__43824\
        );

    \I__10029\ : Span4Mux_h
    port map (
            O => \N__43824\,
            I => \N__43821\
        );

    \I__10028\ : Odrv4
    port map (
            O => \N__43821\,
            I => \nx.n2369\
        );

    \I__10027\ : InMux
    port map (
            O => \N__43818\,
            I => \bfn_15_24_0_\
        );

    \I__10026\ : CascadeMux
    port map (
            O => \N__43815\,
            I => \N__43812\
        );

    \I__10025\ : InMux
    port map (
            O => \N__43812\,
            I => \N__43807\
        );

    \I__10024\ : CascadeMux
    port map (
            O => \N__43811\,
            I => \N__43804\
        );

    \I__10023\ : InMux
    port map (
            O => \N__43810\,
            I => \N__43801\
        );

    \I__10022\ : LocalMux
    port map (
            O => \N__43807\,
            I => \N__43798\
        );

    \I__10021\ : InMux
    port map (
            O => \N__43804\,
            I => \N__43795\
        );

    \I__10020\ : LocalMux
    port map (
            O => \N__43801\,
            I => \N__43792\
        );

    \I__10019\ : Odrv4
    port map (
            O => \N__43798\,
            I => \nx.n2301\
        );

    \I__10018\ : LocalMux
    port map (
            O => \N__43795\,
            I => \nx.n2301\
        );

    \I__10017\ : Odrv4
    port map (
            O => \N__43792\,
            I => \nx.n2301\
        );

    \I__10016\ : InMux
    port map (
            O => \N__43785\,
            I => \N__43782\
        );

    \I__10015\ : LocalMux
    port map (
            O => \N__43782\,
            I => \N__43779\
        );

    \I__10014\ : Odrv4
    port map (
            O => \N__43779\,
            I => \nx.n2368\
        );

    \I__10013\ : InMux
    port map (
            O => \N__43776\,
            I => \nx.n10716\
        );

    \I__10012\ : CascadeMux
    port map (
            O => \N__43773\,
            I => \N__43770\
        );

    \I__10011\ : InMux
    port map (
            O => \N__43770\,
            I => \N__43767\
        );

    \I__10010\ : LocalMux
    port map (
            O => \N__43767\,
            I => \N__43763\
        );

    \I__10009\ : InMux
    port map (
            O => \N__43766\,
            I => \N__43760\
        );

    \I__10008\ : Span4Mux_v
    port map (
            O => \N__43763\,
            I => \N__43757\
        );

    \I__10007\ : LocalMux
    port map (
            O => \N__43760\,
            I => \nx.n2300\
        );

    \I__10006\ : Odrv4
    port map (
            O => \N__43757\,
            I => \nx.n2300\
        );

    \I__10005\ : InMux
    port map (
            O => \N__43752\,
            I => \N__43749\
        );

    \I__10004\ : LocalMux
    port map (
            O => \N__43749\,
            I => \N__43746\
        );

    \I__10003\ : Span4Mux_h
    port map (
            O => \N__43746\,
            I => \N__43743\
        );

    \I__10002\ : Odrv4
    port map (
            O => \N__43743\,
            I => \nx.n2367\
        );

    \I__10001\ : InMux
    port map (
            O => \N__43740\,
            I => \nx.n10717\
        );

    \I__10000\ : CascadeMux
    port map (
            O => \N__43737\,
            I => \N__43734\
        );

    \I__9999\ : InMux
    port map (
            O => \N__43734\,
            I => \N__43730\
        );

    \I__9998\ : CascadeMux
    port map (
            O => \N__43733\,
            I => \N__43727\
        );

    \I__9997\ : LocalMux
    port map (
            O => \N__43730\,
            I => \N__43723\
        );

    \I__9996\ : InMux
    port map (
            O => \N__43727\,
            I => \N__43720\
        );

    \I__9995\ : InMux
    port map (
            O => \N__43726\,
            I => \N__43717\
        );

    \I__9994\ : Odrv4
    port map (
            O => \N__43723\,
            I => \nx.n2299\
        );

    \I__9993\ : LocalMux
    port map (
            O => \N__43720\,
            I => \nx.n2299\
        );

    \I__9992\ : LocalMux
    port map (
            O => \N__43717\,
            I => \nx.n2299\
        );

    \I__9991\ : InMux
    port map (
            O => \N__43710\,
            I => \N__43707\
        );

    \I__9990\ : LocalMux
    port map (
            O => \N__43707\,
            I => \N__43704\
        );

    \I__9989\ : Odrv4
    port map (
            O => \N__43704\,
            I => \nx.n2366\
        );

    \I__9988\ : InMux
    port map (
            O => \N__43701\,
            I => \nx.n10718\
        );

    \I__9987\ : CascadeMux
    port map (
            O => \N__43698\,
            I => \N__43695\
        );

    \I__9986\ : InMux
    port map (
            O => \N__43695\,
            I => \N__43692\
        );

    \I__9985\ : LocalMux
    port map (
            O => \N__43692\,
            I => \N__43689\
        );

    \I__9984\ : Span4Mux_h
    port map (
            O => \N__43689\,
            I => \N__43685\
        );

    \I__9983\ : CascadeMux
    port map (
            O => \N__43688\,
            I => \N__43682\
        );

    \I__9982\ : Span4Mux_h
    port map (
            O => \N__43685\,
            I => \N__43679\
        );

    \I__9981\ : InMux
    port map (
            O => \N__43682\,
            I => \N__43676\
        );

    \I__9980\ : Odrv4
    port map (
            O => \N__43679\,
            I => \nx.n2400\
        );

    \I__9979\ : LocalMux
    port map (
            O => \N__43676\,
            I => \nx.n2400\
        );

    \I__9978\ : CascadeMux
    port map (
            O => \N__43671\,
            I => \nx.n2400_cascade_\
        );

    \I__9977\ : InMux
    port map (
            O => \N__43668\,
            I => \N__43664\
        );

    \I__9976\ : CascadeMux
    port map (
            O => \N__43667\,
            I => \N__43660\
        );

    \I__9975\ : LocalMux
    port map (
            O => \N__43664\,
            I => \N__43657\
        );

    \I__9974\ : InMux
    port map (
            O => \N__43663\,
            I => \N__43654\
        );

    \I__9973\ : InMux
    port map (
            O => \N__43660\,
            I => \N__43651\
        );

    \I__9972\ : Span4Mux_h
    port map (
            O => \N__43657\,
            I => \N__43648\
        );

    \I__9971\ : LocalMux
    port map (
            O => \N__43654\,
            I => \nx.n2403\
        );

    \I__9970\ : LocalMux
    port map (
            O => \N__43651\,
            I => \nx.n2403\
        );

    \I__9969\ : Odrv4
    port map (
            O => \N__43648\,
            I => \nx.n2403\
        );

    \I__9968\ : InMux
    port map (
            O => \N__43641\,
            I => \N__43638\
        );

    \I__9967\ : LocalMux
    port map (
            O => \N__43638\,
            I => \N__43635\
        );

    \I__9966\ : Span4Mux_h
    port map (
            O => \N__43635\,
            I => \N__43632\
        );

    \I__9965\ : Span4Mux_h
    port map (
            O => \N__43632\,
            I => \N__43629\
        );

    \I__9964\ : Odrv4
    port map (
            O => \N__43629\,
            I => \nx.n35_adj_658\
        );

    \I__9963\ : CascadeMux
    port map (
            O => \N__43626\,
            I => \N__43623\
        );

    \I__9962\ : InMux
    port map (
            O => \N__43623\,
            I => \N__43620\
        );

    \I__9961\ : LocalMux
    port map (
            O => \N__43620\,
            I => \N__43617\
        );

    \I__9960\ : Span4Mux_h
    port map (
            O => \N__43617\,
            I => \N__43612\
        );

    \I__9959\ : InMux
    port map (
            O => \N__43616\,
            I => \N__43609\
        );

    \I__9958\ : InMux
    port map (
            O => \N__43615\,
            I => \N__43606\
        );

    \I__9957\ : Odrv4
    port map (
            O => \N__43612\,
            I => \nx.n2402\
        );

    \I__9956\ : LocalMux
    port map (
            O => \N__43609\,
            I => \nx.n2402\
        );

    \I__9955\ : LocalMux
    port map (
            O => \N__43606\,
            I => \nx.n2402\
        );

    \I__9954\ : InMux
    port map (
            O => \N__43599\,
            I => \N__43596\
        );

    \I__9953\ : LocalMux
    port map (
            O => \N__43596\,
            I => \N__43592\
        );

    \I__9952\ : CascadeMux
    port map (
            O => \N__43595\,
            I => \N__43588\
        );

    \I__9951\ : Span4Mux_h
    port map (
            O => \N__43592\,
            I => \N__43585\
        );

    \I__9950\ : InMux
    port map (
            O => \N__43591\,
            I => \N__43582\
        );

    \I__9949\ : InMux
    port map (
            O => \N__43588\,
            I => \N__43579\
        );

    \I__9948\ : Odrv4
    port map (
            O => \N__43585\,
            I => \nx.n2406\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__43582\,
            I => \nx.n2406\
        );

    \I__9946\ : LocalMux
    port map (
            O => \N__43579\,
            I => \nx.n2406\
        );

    \I__9945\ : InMux
    port map (
            O => \N__43572\,
            I => \N__43568\
        );

    \I__9944\ : InMux
    port map (
            O => \N__43571\,
            I => \N__43564\
        );

    \I__9943\ : LocalMux
    port map (
            O => \N__43568\,
            I => \N__43561\
        );

    \I__9942\ : InMux
    port map (
            O => \N__43567\,
            I => \N__43558\
        );

    \I__9941\ : LocalMux
    port map (
            O => \N__43564\,
            I => \N__43555\
        );

    \I__9940\ : Span4Mux_v
    port map (
            O => \N__43561\,
            I => \N__43552\
        );

    \I__9939\ : LocalMux
    port map (
            O => \N__43558\,
            I => \N__43549\
        );

    \I__9938\ : Span4Mux_v
    port map (
            O => \N__43555\,
            I => \N__43545\
        );

    \I__9937\ : Span4Mux_h
    port map (
            O => \N__43552\,
            I => \N__43540\
        );

    \I__9936\ : Span4Mux_h
    port map (
            O => \N__43549\,
            I => \N__43540\
        );

    \I__9935\ : InMux
    port map (
            O => \N__43548\,
            I => \N__43536\
        );

    \I__9934\ : Span4Mux_h
    port map (
            O => \N__43545\,
            I => \N__43533\
        );

    \I__9933\ : Span4Mux_h
    port map (
            O => \N__43540\,
            I => \N__43530\
        );

    \I__9932\ : InMux
    port map (
            O => \N__43539\,
            I => \N__43527\
        );

    \I__9931\ : LocalMux
    port map (
            O => \N__43536\,
            I => \N__43524\
        );

    \I__9930\ : Span4Mux_h
    port map (
            O => \N__43533\,
            I => \N__43521\
        );

    \I__9929\ : Span4Mux_h
    port map (
            O => \N__43530\,
            I => \N__43518\
        );

    \I__9928\ : LocalMux
    port map (
            O => \N__43527\,
            I => \nx.bit_ctr_12\
        );

    \I__9927\ : Odrv4
    port map (
            O => \N__43524\,
            I => \nx.bit_ctr_12\
        );

    \I__9926\ : Odrv4
    port map (
            O => \N__43521\,
            I => \nx.bit_ctr_12\
        );

    \I__9925\ : Odrv4
    port map (
            O => \N__43518\,
            I => \nx.bit_ctr_12\
        );

    \I__9924\ : InMux
    port map (
            O => \N__43509\,
            I => \N__43506\
        );

    \I__9923\ : LocalMux
    port map (
            O => \N__43506\,
            I => \N__43503\
        );

    \I__9922\ : Span4Mux_h
    port map (
            O => \N__43503\,
            I => \N__43500\
        );

    \I__9921\ : Odrv4
    port map (
            O => \N__43500\,
            I => \nx.n2377\
        );

    \I__9920\ : InMux
    port map (
            O => \N__43497\,
            I => \bfn_15_23_0_\
        );

    \I__9919\ : CascadeMux
    port map (
            O => \N__43494\,
            I => \N__43491\
        );

    \I__9918\ : InMux
    port map (
            O => \N__43491\,
            I => \N__43487\
        );

    \I__9917\ : InMux
    port map (
            O => \N__43490\,
            I => \N__43483\
        );

    \I__9916\ : LocalMux
    port map (
            O => \N__43487\,
            I => \N__43480\
        );

    \I__9915\ : InMux
    port map (
            O => \N__43486\,
            I => \N__43477\
        );

    \I__9914\ : LocalMux
    port map (
            O => \N__43483\,
            I => \nx.n2309\
        );

    \I__9913\ : Odrv4
    port map (
            O => \N__43480\,
            I => \nx.n2309\
        );

    \I__9912\ : LocalMux
    port map (
            O => \N__43477\,
            I => \nx.n2309\
        );

    \I__9911\ : CascadeMux
    port map (
            O => \N__43470\,
            I => \N__43467\
        );

    \I__9910\ : InMux
    port map (
            O => \N__43467\,
            I => \N__43464\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__43464\,
            I => \N__43461\
        );

    \I__9908\ : Span4Mux_v
    port map (
            O => \N__43461\,
            I => \N__43458\
        );

    \I__9907\ : Odrv4
    port map (
            O => \N__43458\,
            I => \nx.n2376\
        );

    \I__9906\ : InMux
    port map (
            O => \N__43455\,
            I => \nx.n10708\
        );

    \I__9905\ : CascadeMux
    port map (
            O => \N__43452\,
            I => \N__43448\
        );

    \I__9904\ : CascadeMux
    port map (
            O => \N__43451\,
            I => \N__43444\
        );

    \I__9903\ : InMux
    port map (
            O => \N__43448\,
            I => \N__43441\
        );

    \I__9902\ : InMux
    port map (
            O => \N__43447\,
            I => \N__43438\
        );

    \I__9901\ : InMux
    port map (
            O => \N__43444\,
            I => \N__43435\
        );

    \I__9900\ : LocalMux
    port map (
            O => \N__43441\,
            I => \N__43432\
        );

    \I__9899\ : LocalMux
    port map (
            O => \N__43438\,
            I => \nx.n2308\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__43435\,
            I => \nx.n2308\
        );

    \I__9897\ : Odrv4
    port map (
            O => \N__43432\,
            I => \nx.n2308\
        );

    \I__9896\ : InMux
    port map (
            O => \N__43425\,
            I => \N__43422\
        );

    \I__9895\ : LocalMux
    port map (
            O => \N__43422\,
            I => \N__43419\
        );

    \I__9894\ : Span4Mux_h
    port map (
            O => \N__43419\,
            I => \N__43416\
        );

    \I__9893\ : Odrv4
    port map (
            O => \N__43416\,
            I => \nx.n2375\
        );

    \I__9892\ : InMux
    port map (
            O => \N__43413\,
            I => \nx.n10709\
        );

    \I__9891\ : InMux
    port map (
            O => \N__43410\,
            I => \N__43406\
        );

    \I__9890\ : CascadeMux
    port map (
            O => \N__43409\,
            I => \N__43403\
        );

    \I__9889\ : LocalMux
    port map (
            O => \N__43406\,
            I => \N__43400\
        );

    \I__9888\ : InMux
    port map (
            O => \N__43403\,
            I => \N__43396\
        );

    \I__9887\ : Span4Mux_h
    port map (
            O => \N__43400\,
            I => \N__43393\
        );

    \I__9886\ : InMux
    port map (
            O => \N__43399\,
            I => \N__43390\
        );

    \I__9885\ : LocalMux
    port map (
            O => \N__43396\,
            I => \N__43387\
        );

    \I__9884\ : Odrv4
    port map (
            O => \N__43393\,
            I => \nx.n2307\
        );

    \I__9883\ : LocalMux
    port map (
            O => \N__43390\,
            I => \nx.n2307\
        );

    \I__9882\ : Odrv12
    port map (
            O => \N__43387\,
            I => \nx.n2307\
        );

    \I__9881\ : InMux
    port map (
            O => \N__43380\,
            I => \N__43377\
        );

    \I__9880\ : LocalMux
    port map (
            O => \N__43377\,
            I => \nx.n2374\
        );

    \I__9879\ : InMux
    port map (
            O => \N__43374\,
            I => \nx.n10710\
        );

    \I__9878\ : CascadeMux
    port map (
            O => \N__43371\,
            I => \N__43366\
        );

    \I__9877\ : InMux
    port map (
            O => \N__43370\,
            I => \N__43361\
        );

    \I__9876\ : InMux
    port map (
            O => \N__43369\,
            I => \N__43361\
        );

    \I__9875\ : InMux
    port map (
            O => \N__43366\,
            I => \N__43358\
        );

    \I__9874\ : LocalMux
    port map (
            O => \N__43361\,
            I => \nx.n2306\
        );

    \I__9873\ : LocalMux
    port map (
            O => \N__43358\,
            I => \nx.n2306\
        );

    \I__9872\ : InMux
    port map (
            O => \N__43353\,
            I => \N__43350\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__43350\,
            I => \N__43347\
        );

    \I__9870\ : Span4Mux_h
    port map (
            O => \N__43347\,
            I => \N__43344\
        );

    \I__9869\ : Odrv4
    port map (
            O => \N__43344\,
            I => \nx.n2373\
        );

    \I__9868\ : CascadeMux
    port map (
            O => \N__43341\,
            I => \n19_adj_735_cascade_\
        );

    \I__9867\ : InMux
    port map (
            O => \N__43338\,
            I => \N__43335\
        );

    \I__9866\ : LocalMux
    port map (
            O => \N__43335\,
            I => n13141
        );

    \I__9865\ : CascadeMux
    port map (
            O => \N__43332\,
            I => \N__43329\
        );

    \I__9864\ : InMux
    port map (
            O => \N__43329\,
            I => \N__43326\
        );

    \I__9863\ : LocalMux
    port map (
            O => \N__43326\,
            I => n1
        );

    \I__9862\ : InMux
    port map (
            O => \N__43323\,
            I => \N__43320\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__43320\,
            I => \N__43315\
        );

    \I__9860\ : InMux
    port map (
            O => \N__43319\,
            I => \N__43312\
        );

    \I__9859\ : InMux
    port map (
            O => \N__43318\,
            I => \N__43309\
        );

    \I__9858\ : Span4Mux_v
    port map (
            O => \N__43315\,
            I => \N__43304\
        );

    \I__9857\ : LocalMux
    port map (
            O => \N__43312\,
            I => \N__43304\
        );

    \I__9856\ : LocalMux
    port map (
            O => \N__43309\,
            I => n8_adj_747
        );

    \I__9855\ : Odrv4
    port map (
            O => \N__43304\,
            I => n8_adj_747
        );

    \I__9854\ : CascadeMux
    port map (
            O => \N__43299\,
            I => \N__43296\
        );

    \I__9853\ : InMux
    port map (
            O => \N__43296\,
            I => \N__43290\
        );

    \I__9852\ : InMux
    port map (
            O => \N__43295\,
            I => \N__43286\
        );

    \I__9851\ : InMux
    port map (
            O => \N__43294\,
            I => \N__43283\
        );

    \I__9850\ : InMux
    port map (
            O => \N__43293\,
            I => \N__43280\
        );

    \I__9849\ : LocalMux
    port map (
            O => \N__43290\,
            I => \N__43277\
        );

    \I__9848\ : InMux
    port map (
            O => \N__43289\,
            I => \N__43274\
        );

    \I__9847\ : LocalMux
    port map (
            O => \N__43286\,
            I => \N__43269\
        );

    \I__9846\ : LocalMux
    port map (
            O => \N__43283\,
            I => \N__43269\
        );

    \I__9845\ : LocalMux
    port map (
            O => \N__43280\,
            I => \N__43266\
        );

    \I__9844\ : Span4Mux_v
    port map (
            O => \N__43277\,
            I => \N__43259\
        );

    \I__9843\ : LocalMux
    port map (
            O => \N__43274\,
            I => \N__43259\
        );

    \I__9842\ : Span4Mux_v
    port map (
            O => \N__43269\,
            I => \N__43259\
        );

    \I__9841\ : Span4Mux_v
    port map (
            O => \N__43266\,
            I => \N__43256\
        );

    \I__9840\ : Odrv4
    port map (
            O => \N__43259\,
            I => n9426
        );

    \I__9839\ : Odrv4
    port map (
            O => \N__43256\,
            I => n9426
        );

    \I__9838\ : InMux
    port map (
            O => \N__43251\,
            I => \N__43245\
        );

    \I__9837\ : InMux
    port map (
            O => \N__43250\,
            I => \N__43245\
        );

    \I__9836\ : LocalMux
    port map (
            O => \N__43245\,
            I => \N__43242\
        );

    \I__9835\ : Span4Mux_v
    port map (
            O => \N__43242\,
            I => \N__43239\
        );

    \I__9834\ : Odrv4
    port map (
            O => \N__43239\,
            I => n6178
        );

    \I__9833\ : CascadeMux
    port map (
            O => \N__43236\,
            I => \n7310_cascade_\
        );

    \I__9832\ : InMux
    port map (
            O => \N__43233\,
            I => \N__43229\
        );

    \I__9831\ : InMux
    port map (
            O => \N__43232\,
            I => \N__43225\
        );

    \I__9830\ : LocalMux
    port map (
            O => \N__43229\,
            I => \N__43222\
        );

    \I__9829\ : CascadeMux
    port map (
            O => \N__43228\,
            I => \N__43219\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__43225\,
            I => \N__43216\
        );

    \I__9827\ : Span4Mux_h
    port map (
            O => \N__43222\,
            I => \N__43213\
        );

    \I__9826\ : InMux
    port map (
            O => \N__43219\,
            I => \N__43210\
        );

    \I__9825\ : Span4Mux_v
    port map (
            O => \N__43216\,
            I => \N__43207\
        );

    \I__9824\ : Odrv4
    port map (
            O => \N__43213\,
            I => \nx.n2398\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__43210\,
            I => \nx.n2398\
        );

    \I__9822\ : Odrv4
    port map (
            O => \N__43207\,
            I => \nx.n2398\
        );

    \I__9821\ : InMux
    port map (
            O => \N__43200\,
            I => \N__43195\
        );

    \I__9820\ : InMux
    port map (
            O => \N__43199\,
            I => \N__43192\
        );

    \I__9819\ : CascadeMux
    port map (
            O => \N__43198\,
            I => \N__43189\
        );

    \I__9818\ : LocalMux
    port map (
            O => \N__43195\,
            I => \N__43186\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__43192\,
            I => \N__43183\
        );

    \I__9816\ : InMux
    port map (
            O => \N__43189\,
            I => \N__43180\
        );

    \I__9815\ : Span4Mux_v
    port map (
            O => \N__43186\,
            I => \N__43175\
        );

    \I__9814\ : Span4Mux_h
    port map (
            O => \N__43183\,
            I => \N__43175\
        );

    \I__9813\ : LocalMux
    port map (
            O => \N__43180\,
            I => \N__43170\
        );

    \I__9812\ : Span4Mux_h
    port map (
            O => \N__43175\,
            I => \N__43170\
        );

    \I__9811\ : Odrv4
    port map (
            O => \N__43170\,
            I => \nx.n2397\
        );

    \I__9810\ : InMux
    port map (
            O => \N__43167\,
            I => \N__43164\
        );

    \I__9809\ : LocalMux
    port map (
            O => \N__43164\,
            I => \N__43161\
        );

    \I__9808\ : Span4Mux_v
    port map (
            O => \N__43161\,
            I => \N__43156\
        );

    \I__9807\ : InMux
    port map (
            O => \N__43160\,
            I => \N__43153\
        );

    \I__9806\ : InMux
    port map (
            O => \N__43159\,
            I => \N__43150\
        );

    \I__9805\ : Span4Mux_h
    port map (
            O => \N__43156\,
            I => \N__43146\
        );

    \I__9804\ : LocalMux
    port map (
            O => \N__43153\,
            I => \N__43143\
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__43150\,
            I => \N__43140\
        );

    \I__9802\ : InMux
    port map (
            O => \N__43149\,
            I => \N__43137\
        );

    \I__9801\ : Sp12to4
    port map (
            O => \N__43146\,
            I => \N__43132\
        );

    \I__9800\ : Span12Mux_v
    port map (
            O => \N__43143\,
            I => \N__43132\
        );

    \I__9799\ : Odrv12
    port map (
            O => \N__43140\,
            I => neopxl_color_14
        );

    \I__9798\ : LocalMux
    port map (
            O => \N__43137\,
            I => neopxl_color_14
        );

    \I__9797\ : Odrv12
    port map (
            O => \N__43132\,
            I => neopxl_color_14
        );

    \I__9796\ : CascadeMux
    port map (
            O => \N__43125\,
            I => \N__43122\
        );

    \I__9795\ : InMux
    port map (
            O => \N__43122\,
            I => \N__43119\
        );

    \I__9794\ : LocalMux
    port map (
            O => \N__43119\,
            I => \N__43116\
        );

    \I__9793\ : Span4Mux_v
    port map (
            O => \N__43116\,
            I => \N__43113\
        );

    \I__9792\ : Span4Mux_h
    port map (
            O => \N__43113\,
            I => \N__43110\
        );

    \I__9791\ : Span4Mux_h
    port map (
            O => \N__43110\,
            I => \N__43107\
        );

    \I__9790\ : Span4Mux_h
    port map (
            O => \N__43107\,
            I => \N__43104\
        );

    \I__9789\ : Odrv4
    port map (
            O => \N__43104\,
            I => neopxl_color_prev_14
        );

    \I__9788\ : IoInMux
    port map (
            O => \N__43101\,
            I => \N__43098\
        );

    \I__9787\ : LocalMux
    port map (
            O => \N__43098\,
            I => \N__43095\
        );

    \I__9786\ : Span4Mux_s1_h
    port map (
            O => \N__43095\,
            I => \N__43092\
        );

    \I__9785\ : Sp12to4
    port map (
            O => \N__43092\,
            I => \N__43089\
        );

    \I__9784\ : Span12Mux_v
    port map (
            O => \N__43089\,
            I => \N__43086\
        );

    \I__9783\ : Span12Mux_h
    port map (
            O => \N__43086\,
            I => \N__43081\
        );

    \I__9782\ : InMux
    port map (
            O => \N__43085\,
            I => \N__43078\
        );

    \I__9781\ : InMux
    port map (
            O => \N__43084\,
            I => \N__43075\
        );

    \I__9780\ : Odrv12
    port map (
            O => \N__43081\,
            I => pin_out_16
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__43078\,
            I => pin_out_16
        );

    \I__9778\ : LocalMux
    port map (
            O => \N__43075\,
            I => pin_out_16
        );

    \I__9777\ : CascadeMux
    port map (
            O => \N__43068\,
            I => \n13438_cascade_\
        );

    \I__9776\ : IoInMux
    port map (
            O => \N__43065\,
            I => \N__43062\
        );

    \I__9775\ : LocalMux
    port map (
            O => \N__43062\,
            I => \N__43059\
        );

    \I__9774\ : Span4Mux_s2_v
    port map (
            O => \N__43059\,
            I => \N__43056\
        );

    \I__9773\ : Sp12to4
    port map (
            O => \N__43056\,
            I => \N__43053\
        );

    \I__9772\ : Span12Mux_s7_h
    port map (
            O => \N__43053\,
            I => \N__43049\
        );

    \I__9771\ : InMux
    port map (
            O => \N__43052\,
            I => \N__43045\
        );

    \I__9770\ : Span12Mux_v
    port map (
            O => \N__43049\,
            I => \N__43042\
        );

    \I__9769\ : InMux
    port map (
            O => \N__43048\,
            I => \N__43039\
        );

    \I__9768\ : LocalMux
    port map (
            O => \N__43045\,
            I => \N__43036\
        );

    \I__9767\ : Odrv12
    port map (
            O => \N__43042\,
            I => pin_out_17
        );

    \I__9766\ : LocalMux
    port map (
            O => \N__43039\,
            I => pin_out_17
        );

    \I__9765\ : Odrv4
    port map (
            O => \N__43036\,
            I => pin_out_17
        );

    \I__9764\ : CascadeMux
    port map (
            O => \N__43029\,
            I => \n13441_cascade_\
        );

    \I__9763\ : CascadeMux
    port map (
            O => \N__43026\,
            I => \n13142_cascade_\
        );

    \I__9762\ : InMux
    port map (
            O => \N__43023\,
            I => \N__43020\
        );

    \I__9761\ : LocalMux
    port map (
            O => \N__43020\,
            I => \N__43017\
        );

    \I__9760\ : Odrv4
    port map (
            O => \N__43017\,
            I => n13362
        );

    \I__9759\ : CascadeMux
    port map (
            O => \N__43014\,
            I => \n149_cascade_\
        );

    \I__9758\ : IoInMux
    port map (
            O => \N__43011\,
            I => \N__43008\
        );

    \I__9757\ : LocalMux
    port map (
            O => \N__43008\,
            I => \N__43005\
        );

    \I__9756\ : IoSpan4Mux
    port map (
            O => \N__43005\,
            I => \N__43002\
        );

    \I__9755\ : Span4Mux_s2_v
    port map (
            O => \N__43002\,
            I => \N__42999\
        );

    \I__9754\ : Sp12to4
    port map (
            O => \N__42999\,
            I => \N__42995\
        );

    \I__9753\ : CascadeMux
    port map (
            O => \N__42998\,
            I => \N__42991\
        );

    \I__9752\ : Span12Mux_v
    port map (
            O => \N__42995\,
            I => \N__42988\
        );

    \I__9751\ : InMux
    port map (
            O => \N__42994\,
            I => \N__42983\
        );

    \I__9750\ : InMux
    port map (
            O => \N__42991\,
            I => \N__42983\
        );

    \I__9749\ : Odrv12
    port map (
            O => \N__42988\,
            I => pin_out_19
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__42983\,
            I => pin_out_19
        );

    \I__9747\ : InMux
    port map (
            O => \N__42978\,
            I => \N__42975\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__42975\,
            I => \N__42969\
        );

    \I__9745\ : InMux
    port map (
            O => \N__42974\,
            I => \N__42966\
        );

    \I__9744\ : InMux
    port map (
            O => \N__42973\,
            I => \N__42963\
        );

    \I__9743\ : InMux
    port map (
            O => \N__42972\,
            I => \N__42960\
        );

    \I__9742\ : Span4Mux_v
    port map (
            O => \N__42969\,
            I => \N__42955\
        );

    \I__9741\ : LocalMux
    port map (
            O => \N__42966\,
            I => \N__42955\
        );

    \I__9740\ : LocalMux
    port map (
            O => \N__42963\,
            I => n8_adj_746
        );

    \I__9739\ : LocalMux
    port map (
            O => \N__42960\,
            I => n8_adj_746
        );

    \I__9738\ : Odrv4
    port map (
            O => \N__42955\,
            I => n8_adj_746
        );

    \I__9737\ : InMux
    port map (
            O => \N__42948\,
            I => \N__42942\
        );

    \I__9736\ : InMux
    port map (
            O => \N__42947\,
            I => \N__42942\
        );

    \I__9735\ : LocalMux
    port map (
            O => \N__42942\,
            I => \N__42939\
        );

    \I__9734\ : Span4Mux_h
    port map (
            O => \N__42939\,
            I => \N__42936\
        );

    \I__9733\ : Odrv4
    port map (
            O => \N__42936\,
            I => n6186
        );

    \I__9732\ : InMux
    port map (
            O => \N__42933\,
            I => \N__42930\
        );

    \I__9731\ : LocalMux
    port map (
            O => \N__42930\,
            I => n7326
        );

    \I__9730\ : InMux
    port map (
            O => \N__42927\,
            I => \N__42924\
        );

    \I__9729\ : LocalMux
    port map (
            O => \N__42924\,
            I => n11_adj_734
        );

    \I__9728\ : CascadeMux
    port map (
            O => \N__42921\,
            I => \n11_adj_734_cascade_\
        );

    \I__9727\ : InMux
    port map (
            O => \N__42918\,
            I => \N__42915\
        );

    \I__9726\ : LocalMux
    port map (
            O => \N__42915\,
            I => \N__42912\
        );

    \I__9725\ : Odrv4
    port map (
            O => \N__42912\,
            I => n36_adj_773
        );

    \I__9724\ : IoInMux
    port map (
            O => \N__42909\,
            I => \N__42906\
        );

    \I__9723\ : LocalMux
    port map (
            O => \N__42906\,
            I => \N__42903\
        );

    \I__9722\ : Span4Mux_s2_v
    port map (
            O => \N__42903\,
            I => \N__42900\
        );

    \I__9721\ : Span4Mux_v
    port map (
            O => \N__42900\,
            I => \N__42895\
        );

    \I__9720\ : CascadeMux
    port map (
            O => \N__42899\,
            I => \N__42892\
        );

    \I__9719\ : InMux
    port map (
            O => \N__42898\,
            I => \N__42889\
        );

    \I__9718\ : Sp12to4
    port map (
            O => \N__42895\,
            I => \N__42886\
        );

    \I__9717\ : InMux
    port map (
            O => \N__42892\,
            I => \N__42883\
        );

    \I__9716\ : LocalMux
    port map (
            O => \N__42889\,
            I => \N__42880\
        );

    \I__9715\ : Span12Mux_h
    port map (
            O => \N__42886\,
            I => \N__42877\
        );

    \I__9714\ : LocalMux
    port map (
            O => \N__42883\,
            I => \N__42872\
        );

    \I__9713\ : Span4Mux_v
    port map (
            O => \N__42880\,
            I => \N__42872\
        );

    \I__9712\ : Odrv12
    port map (
            O => \N__42877\,
            I => pin_out_21
        );

    \I__9711\ : Odrv4
    port map (
            O => \N__42872\,
            I => pin_out_21
        );

    \I__9710\ : IoInMux
    port map (
            O => \N__42867\,
            I => \N__42864\
        );

    \I__9709\ : LocalMux
    port map (
            O => \N__42864\,
            I => \N__42860\
        );

    \I__9708\ : CascadeMux
    port map (
            O => \N__42863\,
            I => \N__42857\
        );

    \I__9707\ : Span12Mux_s6_v
    port map (
            O => \N__42860\,
            I => \N__42853\
        );

    \I__9706\ : InMux
    port map (
            O => \N__42857\,
            I => \N__42850\
        );

    \I__9705\ : InMux
    port map (
            O => \N__42856\,
            I => \N__42847\
        );

    \I__9704\ : Span12Mux_h
    port map (
            O => \N__42853\,
            I => \N__42844\
        );

    \I__9703\ : LocalMux
    port map (
            O => \N__42850\,
            I => \N__42841\
        );

    \I__9702\ : LocalMux
    port map (
            O => \N__42847\,
            I => \N__42838\
        );

    \I__9701\ : Odrv12
    port map (
            O => \N__42844\,
            I => pin_out_20
        );

    \I__9700\ : Odrv4
    port map (
            O => \N__42841\,
            I => pin_out_20
        );

    \I__9699\ : Odrv4
    port map (
            O => \N__42838\,
            I => pin_out_20
        );

    \I__9698\ : InMux
    port map (
            O => \N__42831\,
            I => \N__42827\
        );

    \I__9697\ : InMux
    port map (
            O => \N__42830\,
            I => \N__42824\
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__42827\,
            I => \N__42821\
        );

    \I__9695\ : LocalMux
    port map (
            O => \N__42824\,
            I => \N__42818\
        );

    \I__9694\ : Span4Mux_v
    port map (
            O => \N__42821\,
            I => \N__42815\
        );

    \I__9693\ : Span4Mux_v
    port map (
            O => \N__42818\,
            I => \N__42812\
        );

    \I__9692\ : Odrv4
    port map (
            O => \N__42815\,
            I => n10_adj_736
        );

    \I__9691\ : Odrv4
    port map (
            O => \N__42812\,
            I => n10_adj_736
        );

    \I__9690\ : InMux
    port map (
            O => \N__42807\,
            I => \N__42804\
        );

    \I__9689\ : LocalMux
    port map (
            O => \N__42804\,
            I => \N__42801\
        );

    \I__9688\ : Span4Mux_v
    port map (
            O => \N__42801\,
            I => \N__42797\
        );

    \I__9687\ : InMux
    port map (
            O => \N__42800\,
            I => \N__42794\
        );

    \I__9686\ : Span4Mux_h
    port map (
            O => \N__42797\,
            I => \N__42791\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__42794\,
            I => \N__42788\
        );

    \I__9684\ : Sp12to4
    port map (
            O => \N__42791\,
            I => \N__42785\
        );

    \I__9683\ : Span12Mux_h
    port map (
            O => \N__42788\,
            I => \N__42782\
        );

    \I__9682\ : Span12Mux_h
    port map (
            O => \N__42785\,
            I => \N__42779\
        );

    \I__9681\ : Span12Mux_v
    port map (
            O => \N__42782\,
            I => \N__42776\
        );

    \I__9680\ : Span12Mux_v
    port map (
            O => \N__42779\,
            I => \N__42771\
        );

    \I__9679\ : Span12Mux_h
    port map (
            O => \N__42776\,
            I => \N__42771\
        );

    \I__9678\ : Odrv12
    port map (
            O => \N__42771\,
            I => pin_in_14
        );

    \I__9677\ : CascadeMux
    port map (
            O => \N__42768\,
            I => \N__42762\
        );

    \I__9676\ : InMux
    port map (
            O => \N__42767\,
            I => \N__42759\
        );

    \I__9675\ : InMux
    port map (
            O => \N__42766\,
            I => \N__42756\
        );

    \I__9674\ : InMux
    port map (
            O => \N__42765\,
            I => \N__42753\
        );

    \I__9673\ : InMux
    port map (
            O => \N__42762\,
            I => \N__42750\
        );

    \I__9672\ : LocalMux
    port map (
            O => \N__42759\,
            I => \N__42747\
        );

    \I__9671\ : LocalMux
    port map (
            O => \N__42756\,
            I => \N__42742\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__42753\,
            I => \N__42742\
        );

    \I__9669\ : LocalMux
    port map (
            O => \N__42750\,
            I => n7145
        );

    \I__9668\ : Odrv4
    port map (
            O => \N__42747\,
            I => n7145
        );

    \I__9667\ : Odrv4
    port map (
            O => \N__42742\,
            I => n7145
        );

    \I__9666\ : InMux
    port map (
            O => \N__42735\,
            I => \N__42732\
        );

    \I__9665\ : LocalMux
    port map (
            O => \N__42732\,
            I => \N__42729\
        );

    \I__9664\ : Odrv4
    port map (
            O => \N__42729\,
            I => n7314
        );

    \I__9663\ : InMux
    port map (
            O => \N__42726\,
            I => \N__42722\
        );

    \I__9662\ : CascadeMux
    port map (
            O => \N__42725\,
            I => \N__42719\
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__42722\,
            I => \N__42716\
        );

    \I__9660\ : InMux
    port map (
            O => \N__42719\,
            I => \N__42712\
        );

    \I__9659\ : Span4Mux_h
    port map (
            O => \N__42716\,
            I => \N__42709\
        );

    \I__9658\ : InMux
    port map (
            O => \N__42715\,
            I => \N__42706\
        );

    \I__9657\ : LocalMux
    port map (
            O => \N__42712\,
            I => \N__42703\
        );

    \I__9656\ : Span4Mux_h
    port map (
            O => \N__42709\,
            I => \N__42696\
        );

    \I__9655\ : LocalMux
    port map (
            O => \N__42706\,
            I => \N__42696\
        );

    \I__9654\ : Span4Mux_h
    port map (
            O => \N__42703\,
            I => \N__42693\
        );

    \I__9653\ : CascadeMux
    port map (
            O => \N__42702\,
            I => \N__42690\
        );

    \I__9652\ : CascadeMux
    port map (
            O => \N__42701\,
            I => \N__42687\
        );

    \I__9651\ : Span4Mux_v
    port map (
            O => \N__42696\,
            I => \N__42684\
        );

    \I__9650\ : Span4Mux_h
    port map (
            O => \N__42693\,
            I => \N__42681\
        );

    \I__9649\ : InMux
    port map (
            O => \N__42690\,
            I => \N__42676\
        );

    \I__9648\ : InMux
    port map (
            O => \N__42687\,
            I => \N__42676\
        );

    \I__9647\ : Span4Mux_h
    port map (
            O => \N__42684\,
            I => \N__42673\
        );

    \I__9646\ : Odrv4
    port map (
            O => \N__42681\,
            I => n6
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__42676\,
            I => n6
        );

    \I__9644\ : Odrv4
    port map (
            O => \N__42673\,
            I => n6
        );

    \I__9643\ : InMux
    port map (
            O => \N__42666\,
            I => \N__42660\
        );

    \I__9642\ : InMux
    port map (
            O => \N__42665\,
            I => \N__42660\
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__42660\,
            I => \N__42657\
        );

    \I__9640\ : Span4Mux_v
    port map (
            O => \N__42657\,
            I => \N__42654\
        );

    \I__9639\ : Span4Mux_h
    port map (
            O => \N__42654\,
            I => \N__42651\
        );

    \I__9638\ : Odrv4
    port map (
            O => \N__42651\,
            I => n6182
        );

    \I__9637\ : CascadeMux
    port map (
            O => \N__42648\,
            I => \n7318_cascade_\
        );

    \I__9636\ : CascadeMux
    port map (
            O => \N__42645\,
            I => \N__42642\
        );

    \I__9635\ : InMux
    port map (
            O => \N__42642\,
            I => \N__42637\
        );

    \I__9634\ : CascadeMux
    port map (
            O => \N__42641\,
            I => \N__42634\
        );

    \I__9633\ : InMux
    port map (
            O => \N__42640\,
            I => \N__42630\
        );

    \I__9632\ : LocalMux
    port map (
            O => \N__42637\,
            I => \N__42627\
        );

    \I__9631\ : InMux
    port map (
            O => \N__42634\,
            I => \N__42622\
        );

    \I__9630\ : CascadeMux
    port map (
            O => \N__42633\,
            I => \N__42619\
        );

    \I__9629\ : LocalMux
    port map (
            O => \N__42630\,
            I => \N__42614\
        );

    \I__9628\ : Span4Mux_v
    port map (
            O => \N__42627\,
            I => \N__42614\
        );

    \I__9627\ : CascadeMux
    port map (
            O => \N__42626\,
            I => \N__42611\
        );

    \I__9626\ : InMux
    port map (
            O => \N__42625\,
            I => \N__42606\
        );

    \I__9625\ : LocalMux
    port map (
            O => \N__42622\,
            I => \N__42603\
        );

    \I__9624\ : InMux
    port map (
            O => \N__42619\,
            I => \N__42600\
        );

    \I__9623\ : Span4Mux_h
    port map (
            O => \N__42614\,
            I => \N__42597\
        );

    \I__9622\ : InMux
    port map (
            O => \N__42611\,
            I => \N__42594\
        );

    \I__9621\ : InMux
    port map (
            O => \N__42610\,
            I => \N__42589\
        );

    \I__9620\ : InMux
    port map (
            O => \N__42609\,
            I => \N__42589\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__42606\,
            I => n9_adj_733
        );

    \I__9618\ : Odrv4
    port map (
            O => \N__42603\,
            I => n9_adj_733
        );

    \I__9617\ : LocalMux
    port map (
            O => \N__42600\,
            I => n9_adj_733
        );

    \I__9616\ : Odrv4
    port map (
            O => \N__42597\,
            I => n9_adj_733
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__42594\,
            I => n9_adj_733
        );

    \I__9614\ : LocalMux
    port map (
            O => \N__42589\,
            I => n9_adj_733
        );

    \I__9613\ : CascadeMux
    port map (
            O => \N__42576\,
            I => \N__42572\
        );

    \I__9612\ : InMux
    port map (
            O => \N__42575\,
            I => \N__42567\
        );

    \I__9611\ : InMux
    port map (
            O => \N__42572\,
            I => \N__42567\
        );

    \I__9610\ : LocalMux
    port map (
            O => \N__42567\,
            I => \N__42564\
        );

    \I__9609\ : Odrv4
    port map (
            O => \N__42564\,
            I => n6188
        );

    \I__9608\ : InMux
    port map (
            O => \N__42561\,
            I => \N__42558\
        );

    \I__9607\ : LocalMux
    port map (
            O => \N__42558\,
            I => n7330
        );

    \I__9606\ : IoInMux
    port map (
            O => \N__42555\,
            I => \N__42552\
        );

    \I__9605\ : LocalMux
    port map (
            O => \N__42552\,
            I => \N__42549\
        );

    \I__9604\ : IoSpan4Mux
    port map (
            O => \N__42549\,
            I => \N__42546\
        );

    \I__9603\ : Sp12to4
    port map (
            O => \N__42546\,
            I => \N__42543\
        );

    \I__9602\ : Span12Mux_v
    port map (
            O => \N__42543\,
            I => \N__42539\
        );

    \I__9601\ : InMux
    port map (
            O => \N__42542\,
            I => \N__42535\
        );

    \I__9600\ : Span12Mux_h
    port map (
            O => \N__42539\,
            I => \N__42532\
        );

    \I__9599\ : InMux
    port map (
            O => \N__42538\,
            I => \N__42529\
        );

    \I__9598\ : LocalMux
    port map (
            O => \N__42535\,
            I => \N__42526\
        );

    \I__9597\ : Odrv12
    port map (
            O => \N__42532\,
            I => pin_out_18
        );

    \I__9596\ : LocalMux
    port map (
            O => \N__42529\,
            I => pin_out_18
        );

    \I__9595\ : Odrv4
    port map (
            O => \N__42526\,
            I => pin_out_18
        );

    \I__9594\ : InMux
    port map (
            O => \N__42519\,
            I => \N__42513\
        );

    \I__9593\ : InMux
    port map (
            O => \N__42518\,
            I => \N__42513\
        );

    \I__9592\ : LocalMux
    port map (
            O => \N__42513\,
            I => n6176
        );

    \I__9591\ : CascadeMux
    port map (
            O => \N__42510\,
            I => \n7306_cascade_\
        );

    \I__9590\ : IoInMux
    port map (
            O => \N__42507\,
            I => \N__42504\
        );

    \I__9589\ : LocalMux
    port map (
            O => \N__42504\,
            I => \N__42501\
        );

    \I__9588\ : Span4Mux_s2_v
    port map (
            O => \N__42501\,
            I => \N__42498\
        );

    \I__9587\ : Sp12to4
    port map (
            O => \N__42498\,
            I => \N__42495\
        );

    \I__9586\ : Span12Mux_s8_h
    port map (
            O => \N__42495\,
            I => \N__42491\
        );

    \I__9585\ : CascadeMux
    port map (
            O => \N__42494\,
            I => \N__42488\
        );

    \I__9584\ : Span12Mux_v
    port map (
            O => \N__42491\,
            I => \N__42484\
        );

    \I__9583\ : InMux
    port map (
            O => \N__42488\,
            I => \N__42481\
        );

    \I__9582\ : InMux
    port map (
            O => \N__42487\,
            I => \N__42478\
        );

    \I__9581\ : Odrv12
    port map (
            O => \N__42484\,
            I => pin_out_9
        );

    \I__9580\ : LocalMux
    port map (
            O => \N__42481\,
            I => pin_out_9
        );

    \I__9579\ : LocalMux
    port map (
            O => \N__42478\,
            I => pin_out_9
        );

    \I__9578\ : InMux
    port map (
            O => \N__42471\,
            I => \N__42468\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__42468\,
            I => \N__42465\
        );

    \I__9576\ : Span4Mux_v
    port map (
            O => \N__42465\,
            I => \N__42462\
        );

    \I__9575\ : Odrv4
    port map (
            O => \N__42462\,
            I => n13162
        );

    \I__9574\ : CascadeMux
    port map (
            O => \N__42459\,
            I => \n13161_cascade_\
        );

    \I__9573\ : InMux
    port map (
            O => \N__42456\,
            I => \N__42451\
        );

    \I__9572\ : InMux
    port map (
            O => \N__42455\,
            I => \N__42448\
        );

    \I__9571\ : InMux
    port map (
            O => \N__42454\,
            I => \N__42445\
        );

    \I__9570\ : LocalMux
    port map (
            O => \N__42451\,
            I => \N__42442\
        );

    \I__9569\ : LocalMux
    port map (
            O => \N__42448\,
            I => \N__42439\
        );

    \I__9568\ : LocalMux
    port map (
            O => \N__42445\,
            I => \N__42436\
        );

    \I__9567\ : Span4Mux_h
    port map (
            O => \N__42442\,
            I => \N__42433\
        );

    \I__9566\ : Odrv4
    port map (
            O => \N__42439\,
            I => n8_adj_751
        );

    \I__9565\ : Odrv4
    port map (
            O => \N__42436\,
            I => n8_adj_751
        );

    \I__9564\ : Odrv4
    port map (
            O => \N__42433\,
            I => n8_adj_751
        );

    \I__9563\ : InMux
    port map (
            O => \N__42426\,
            I => \N__42422\
        );

    \I__9562\ : InMux
    port map (
            O => \N__42425\,
            I => \N__42419\
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__42422\,
            I => n6164
        );

    \I__9560\ : LocalMux
    port map (
            O => \N__42419\,
            I => n6164
        );

    \I__9559\ : CascadeMux
    port map (
            O => \N__42414\,
            I => \n7282_cascade_\
        );

    \I__9558\ : IoInMux
    port map (
            O => \N__42411\,
            I => \N__42408\
        );

    \I__9557\ : LocalMux
    port map (
            O => \N__42408\,
            I => \N__42405\
        );

    \I__9556\ : Span12Mux_s4_v
    port map (
            O => \N__42405\,
            I => \N__42402\
        );

    \I__9555\ : Span12Mux_v
    port map (
            O => \N__42402\,
            I => \N__42397\
        );

    \I__9554\ : InMux
    port map (
            O => \N__42401\,
            I => \N__42392\
        );

    \I__9553\ : InMux
    port map (
            O => \N__42400\,
            I => \N__42392\
        );

    \I__9552\ : Odrv12
    port map (
            O => \N__42397\,
            I => pin_out_8
        );

    \I__9551\ : LocalMux
    port map (
            O => \N__42392\,
            I => pin_out_8
        );

    \I__9550\ : CascadeMux
    port map (
            O => \N__42387\,
            I => \N__42383\
        );

    \I__9549\ : InMux
    port map (
            O => \N__42386\,
            I => \N__42380\
        );

    \I__9548\ : InMux
    port map (
            O => \N__42383\,
            I => \N__42377\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__42380\,
            I => n6184
        );

    \I__9546\ : LocalMux
    port map (
            O => \N__42377\,
            I => n6184
        );

    \I__9545\ : CascadeMux
    port map (
            O => \N__42372\,
            I => \n7322_cascade_\
        );

    \I__9544\ : InMux
    port map (
            O => \N__42369\,
            I => \N__42366\
        );

    \I__9543\ : LocalMux
    port map (
            O => \N__42366\,
            I => n13471
        );

    \I__9542\ : InMux
    port map (
            O => \N__42363\,
            I => \N__42360\
        );

    \I__9541\ : LocalMux
    port map (
            O => \N__42360\,
            I => \N__42357\
        );

    \I__9540\ : Odrv12
    port map (
            O => \N__42357\,
            I => n13465
        );

    \I__9539\ : CascadeMux
    port map (
            O => \N__42354\,
            I => \n13177_cascade_\
        );

    \I__9538\ : IoInMux
    port map (
            O => \N__42351\,
            I => \N__42348\
        );

    \I__9537\ : LocalMux
    port map (
            O => \N__42348\,
            I => \N__42345\
        );

    \I__9536\ : Span4Mux_s0_v
    port map (
            O => \N__42345\,
            I => \N__42342\
        );

    \I__9535\ : Sp12to4
    port map (
            O => \N__42342\,
            I => \N__42339\
        );

    \I__9534\ : Span12Mux_h
    port map (
            O => \N__42339\,
            I => \N__42336\
        );

    \I__9533\ : Odrv12
    port map (
            O => \N__42336\,
            I => \LED_c\
        );

    \I__9532\ : InMux
    port map (
            O => \N__42333\,
            I => \N__42330\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__42330\,
            I => n13176
        );

    \I__9530\ : InMux
    port map (
            O => \N__42327\,
            I => \N__42321\
        );

    \I__9529\ : InMux
    port map (
            O => \N__42326\,
            I => \N__42318\
        );

    \I__9528\ : InMux
    port map (
            O => \N__42325\,
            I => \N__42315\
        );

    \I__9527\ : InMux
    port map (
            O => \N__42324\,
            I => \N__42312\
        );

    \I__9526\ : LocalMux
    port map (
            O => \N__42321\,
            I => n21_adj_741
        );

    \I__9525\ : LocalMux
    port map (
            O => \N__42318\,
            I => n21_adj_741
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__42315\,
            I => n21_adj_741
        );

    \I__9523\ : LocalMux
    port map (
            O => \N__42312\,
            I => n21_adj_741
        );

    \I__9522\ : InMux
    port map (
            O => \N__42303\,
            I => \N__42300\
        );

    \I__9521\ : LocalMux
    port map (
            O => \N__42300\,
            I => n6172
        );

    \I__9520\ : InMux
    port map (
            O => \N__42297\,
            I => \N__42294\
        );

    \I__9519\ : LocalMux
    port map (
            O => \N__42294\,
            I => n7298
        );

    \I__9518\ : CascadeMux
    port map (
            O => \N__42291\,
            I => \n6172_cascade_\
        );

    \I__9517\ : CascadeMux
    port map (
            O => \N__42288\,
            I => \N__42285\
        );

    \I__9516\ : InMux
    port map (
            O => \N__42285\,
            I => \N__42281\
        );

    \I__9515\ : InMux
    port map (
            O => \N__42284\,
            I => \N__42278\
        );

    \I__9514\ : LocalMux
    port map (
            O => \N__42281\,
            I => \N__42275\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__42278\,
            I => n6174
        );

    \I__9512\ : Odrv12
    port map (
            O => \N__42275\,
            I => n6174
        );

    \I__9511\ : InMux
    port map (
            O => \N__42270\,
            I => \N__42267\
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__42267\,
            I => n7302
        );

    \I__9509\ : CascadeMux
    port map (
            O => \N__42264\,
            I => \N__42257\
        );

    \I__9508\ : CascadeMux
    port map (
            O => \N__42263\,
            I => \N__42253\
        );

    \I__9507\ : InMux
    port map (
            O => \N__42262\,
            I => \N__42249\
        );

    \I__9506\ : InMux
    port map (
            O => \N__42261\,
            I => \N__42246\
        );

    \I__9505\ : InMux
    port map (
            O => \N__42260\,
            I => \N__42241\
        );

    \I__9504\ : InMux
    port map (
            O => \N__42257\,
            I => \N__42241\
        );

    \I__9503\ : InMux
    port map (
            O => \N__42256\,
            I => \N__42236\
        );

    \I__9502\ : InMux
    port map (
            O => \N__42253\,
            I => \N__42236\
        );

    \I__9501\ : InMux
    port map (
            O => \N__42252\,
            I => \N__42233\
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__42249\,
            I => n7_adj_753
        );

    \I__9499\ : LocalMux
    port map (
            O => \N__42246\,
            I => n7_adj_753
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__42241\,
            I => n7_adj_753
        );

    \I__9497\ : LocalMux
    port map (
            O => \N__42236\,
            I => n7_adj_753
        );

    \I__9496\ : LocalMux
    port map (
            O => \N__42233\,
            I => n7_adj_753
        );

    \I__9495\ : InMux
    port map (
            O => \N__42222\,
            I => \N__42219\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__42219\,
            I => \N__42216\
        );

    \I__9493\ : Odrv4
    port map (
            O => \N__42216\,
            I => \nx.n2271\
        );

    \I__9492\ : CascadeMux
    port map (
            O => \N__42213\,
            I => \N__42210\
        );

    \I__9491\ : InMux
    port map (
            O => \N__42210\,
            I => \N__42205\
        );

    \I__9490\ : InMux
    port map (
            O => \N__42209\,
            I => \N__42202\
        );

    \I__9489\ : InMux
    port map (
            O => \N__42208\,
            I => \N__42199\
        );

    \I__9488\ : LocalMux
    port map (
            O => \N__42205\,
            I => \N__42194\
        );

    \I__9487\ : LocalMux
    port map (
            O => \N__42202\,
            I => \N__42194\
        );

    \I__9486\ : LocalMux
    port map (
            O => \N__42199\,
            I => \nx.n2204\
        );

    \I__9485\ : Odrv4
    port map (
            O => \N__42194\,
            I => \nx.n2204\
        );

    \I__9484\ : InMux
    port map (
            O => \N__42189\,
            I => \N__42186\
        );

    \I__9483\ : LocalMux
    port map (
            O => \N__42186\,
            I => \nx.n2265\
        );

    \I__9482\ : InMux
    port map (
            O => \N__42183\,
            I => \N__42179\
        );

    \I__9481\ : CascadeMux
    port map (
            O => \N__42182\,
            I => \N__42176\
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__42179\,
            I => \N__42173\
        );

    \I__9479\ : InMux
    port map (
            O => \N__42176\,
            I => \N__42170\
        );

    \I__9478\ : Span4Mux_h
    port map (
            O => \N__42173\,
            I => \N__42164\
        );

    \I__9477\ : LocalMux
    port map (
            O => \N__42170\,
            I => \N__42164\
        );

    \I__9476\ : InMux
    port map (
            O => \N__42169\,
            I => \N__42161\
        );

    \I__9475\ : Odrv4
    port map (
            O => \N__42164\,
            I => \nx.n2198\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__42161\,
            I => \nx.n2198\
        );

    \I__9473\ : CascadeMux
    port map (
            O => \N__42156\,
            I => \nx.n2297_cascade_\
        );

    \I__9472\ : InMux
    port map (
            O => \N__42153\,
            I => \N__42150\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__42150\,
            I => \N__42147\
        );

    \I__9470\ : Odrv4
    port map (
            O => \N__42147\,
            I => \nx.n9650\
        );

    \I__9469\ : InMux
    port map (
            O => \N__42144\,
            I => \N__42141\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__42141\,
            I => \N__42138\
        );

    \I__9467\ : Odrv4
    port map (
            O => \N__42138\,
            I => \nx.n31_adj_645\
        );

    \I__9466\ : InMux
    port map (
            O => \N__42135\,
            I => \N__42132\
        );

    \I__9465\ : LocalMux
    port map (
            O => \N__42132\,
            I => \nx.n2269\
        );

    \I__9464\ : CascadeMux
    port map (
            O => \N__42129\,
            I => \N__42125\
        );

    \I__9463\ : InMux
    port map (
            O => \N__42128\,
            I => \N__42121\
        );

    \I__9462\ : InMux
    port map (
            O => \N__42125\,
            I => \N__42118\
        );

    \I__9461\ : CascadeMux
    port map (
            O => \N__42124\,
            I => \N__42115\
        );

    \I__9460\ : LocalMux
    port map (
            O => \N__42121\,
            I => \N__42110\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__42118\,
            I => \N__42110\
        );

    \I__9458\ : InMux
    port map (
            O => \N__42115\,
            I => \N__42107\
        );

    \I__9457\ : Span4Mux_h
    port map (
            O => \N__42110\,
            I => \N__42104\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__42107\,
            I => \nx.n2202\
        );

    \I__9455\ : Odrv4
    port map (
            O => \N__42104\,
            I => \nx.n2202\
        );

    \I__9454\ : InMux
    port map (
            O => \N__42099\,
            I => \N__42096\
        );

    \I__9453\ : LocalMux
    port map (
            O => \N__42096\,
            I => \nx.n2267\
        );

    \I__9452\ : CascadeMux
    port map (
            O => \N__42093\,
            I => \N__42090\
        );

    \I__9451\ : InMux
    port map (
            O => \N__42090\,
            I => \N__42086\
        );

    \I__9450\ : CascadeMux
    port map (
            O => \N__42089\,
            I => \N__42083\
        );

    \I__9449\ : LocalMux
    port map (
            O => \N__42086\,
            I => \N__42080\
        );

    \I__9448\ : InMux
    port map (
            O => \N__42083\,
            I => \N__42077\
        );

    \I__9447\ : Span4Mux_h
    port map (
            O => \N__42080\,
            I => \N__42071\
        );

    \I__9446\ : LocalMux
    port map (
            O => \N__42077\,
            I => \N__42071\
        );

    \I__9445\ : InMux
    port map (
            O => \N__42076\,
            I => \N__42068\
        );

    \I__9444\ : Odrv4
    port map (
            O => \N__42071\,
            I => \nx.n2200\
        );

    \I__9443\ : LocalMux
    port map (
            O => \N__42068\,
            I => \nx.n2200\
        );

    \I__9442\ : InMux
    port map (
            O => \N__42063\,
            I => \N__42060\
        );

    \I__9441\ : LocalMux
    port map (
            O => \N__42060\,
            I => \nx.n2266\
        );

    \I__9440\ : InMux
    port map (
            O => \N__42057\,
            I => \N__42053\
        );

    \I__9439\ : CascadeMux
    port map (
            O => \N__42056\,
            I => \N__42049\
        );

    \I__9438\ : LocalMux
    port map (
            O => \N__42053\,
            I => \N__42046\
        );

    \I__9437\ : InMux
    port map (
            O => \N__42052\,
            I => \N__42043\
        );

    \I__9436\ : InMux
    port map (
            O => \N__42049\,
            I => \N__42040\
        );

    \I__9435\ : Span4Mux_h
    port map (
            O => \N__42046\,
            I => \N__42035\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__42043\,
            I => \N__42035\
        );

    \I__9433\ : LocalMux
    port map (
            O => \N__42040\,
            I => \nx.n2199\
        );

    \I__9432\ : Odrv4
    port map (
            O => \N__42035\,
            I => \nx.n2199\
        );

    \I__9431\ : InMux
    port map (
            O => \N__42030\,
            I => \N__42027\
        );

    \I__9430\ : LocalMux
    port map (
            O => \N__42027\,
            I => \nx.n2260\
        );

    \I__9429\ : CascadeMux
    port map (
            O => \N__42024\,
            I => \N__42021\
        );

    \I__9428\ : InMux
    port map (
            O => \N__42021\,
            I => \N__42017\
        );

    \I__9427\ : CascadeMux
    port map (
            O => \N__42020\,
            I => \N__42014\
        );

    \I__9426\ : LocalMux
    port map (
            O => \N__42017\,
            I => \N__42010\
        );

    \I__9425\ : InMux
    port map (
            O => \N__42014\,
            I => \N__42007\
        );

    \I__9424\ : CascadeMux
    port map (
            O => \N__42013\,
            I => \N__42004\
        );

    \I__9423\ : Span4Mux_v
    port map (
            O => \N__42010\,
            I => \N__41999\
        );

    \I__9422\ : LocalMux
    port map (
            O => \N__42007\,
            I => \N__41999\
        );

    \I__9421\ : InMux
    port map (
            O => \N__42004\,
            I => \N__41996\
        );

    \I__9420\ : Odrv4
    port map (
            O => \N__41999\,
            I => \nx.n2193\
        );

    \I__9419\ : LocalMux
    port map (
            O => \N__41996\,
            I => \nx.n2193\
        );

    \I__9418\ : CascadeMux
    port map (
            O => \N__41991\,
            I => \N__41985\
        );

    \I__9417\ : CascadeMux
    port map (
            O => \N__41990\,
            I => \N__41982\
        );

    \I__9416\ : CascadeMux
    port map (
            O => \N__41989\,
            I => \N__41978\
        );

    \I__9415\ : CascadeMux
    port map (
            O => \N__41988\,
            I => \N__41969\
        );

    \I__9414\ : InMux
    port map (
            O => \N__41985\,
            I => \N__41958\
        );

    \I__9413\ : InMux
    port map (
            O => \N__41982\,
            I => \N__41958\
        );

    \I__9412\ : InMux
    port map (
            O => \N__41981\,
            I => \N__41958\
        );

    \I__9411\ : InMux
    port map (
            O => \N__41978\,
            I => \N__41958\
        );

    \I__9410\ : InMux
    port map (
            O => \N__41977\,
            I => \N__41958\
        );

    \I__9409\ : CascadeMux
    port map (
            O => \N__41976\,
            I => \N__41954\
        );

    \I__9408\ : InMux
    port map (
            O => \N__41975\,
            I => \N__41950\
        );

    \I__9407\ : CascadeMux
    port map (
            O => \N__41974\,
            I => \N__41945\
        );

    \I__9406\ : InMux
    port map (
            O => \N__41973\,
            I => \N__41940\
        );

    \I__9405\ : InMux
    port map (
            O => \N__41972\,
            I => \N__41940\
        );

    \I__9404\ : InMux
    port map (
            O => \N__41969\,
            I => \N__41937\
        );

    \I__9403\ : LocalMux
    port map (
            O => \N__41958\,
            I => \N__41934\
        );

    \I__9402\ : CascadeMux
    port map (
            O => \N__41957\,
            I => \N__41929\
        );

    \I__9401\ : InMux
    port map (
            O => \N__41954\,
            I => \N__41923\
        );

    \I__9400\ : InMux
    port map (
            O => \N__41953\,
            I => \N__41923\
        );

    \I__9399\ : LocalMux
    port map (
            O => \N__41950\,
            I => \N__41920\
        );

    \I__9398\ : InMux
    port map (
            O => \N__41949\,
            I => \N__41913\
        );

    \I__9397\ : InMux
    port map (
            O => \N__41948\,
            I => \N__41913\
        );

    \I__9396\ : InMux
    port map (
            O => \N__41945\,
            I => \N__41913\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__41940\,
            I => \N__41910\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__41937\,
            I => \N__41905\
        );

    \I__9393\ : Span4Mux_h
    port map (
            O => \N__41934\,
            I => \N__41905\
        );

    \I__9392\ : InMux
    port map (
            O => \N__41933\,
            I => \N__41896\
        );

    \I__9391\ : InMux
    port map (
            O => \N__41932\,
            I => \N__41896\
        );

    \I__9390\ : InMux
    port map (
            O => \N__41929\,
            I => \N__41896\
        );

    \I__9389\ : InMux
    port map (
            O => \N__41928\,
            I => \N__41896\
        );

    \I__9388\ : LocalMux
    port map (
            O => \N__41923\,
            I => \nx.n2225\
        );

    \I__9387\ : Odrv4
    port map (
            O => \N__41920\,
            I => \nx.n2225\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__41913\,
            I => \nx.n2225\
        );

    \I__9385\ : Odrv4
    port map (
            O => \N__41910\,
            I => \nx.n2225\
        );

    \I__9384\ : Odrv4
    port map (
            O => \N__41905\,
            I => \nx.n2225\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__41896\,
            I => \nx.n2225\
        );

    \I__9382\ : InMux
    port map (
            O => \N__41883\,
            I => \N__41878\
        );

    \I__9381\ : CascadeMux
    port map (
            O => \N__41882\,
            I => \N__41875\
        );

    \I__9380\ : InMux
    port map (
            O => \N__41881\,
            I => \N__41872\
        );

    \I__9379\ : LocalMux
    port map (
            O => \N__41878\,
            I => \N__41869\
        );

    \I__9378\ : InMux
    port map (
            O => \N__41875\,
            I => \N__41866\
        );

    \I__9377\ : LocalMux
    port map (
            O => \N__41872\,
            I => \N__41863\
        );

    \I__9376\ : Span4Mux_h
    port map (
            O => \N__41869\,
            I => \N__41860\
        );

    \I__9375\ : LocalMux
    port map (
            O => \N__41866\,
            I => \N__41857\
        );

    \I__9374\ : Span4Mux_v
    port map (
            O => \N__41863\,
            I => \N__41852\
        );

    \I__9373\ : Span4Mux_h
    port map (
            O => \N__41860\,
            I => \N__41852\
        );

    \I__9372\ : Odrv4
    port map (
            O => \N__41857\,
            I => \nx.n2396\
        );

    \I__9371\ : Odrv4
    port map (
            O => \N__41852\,
            I => \nx.n2396\
        );

    \I__9370\ : CascadeMux
    port map (
            O => \N__41847\,
            I => \N__41844\
        );

    \I__9369\ : InMux
    port map (
            O => \N__41844\,
            I => \N__41840\
        );

    \I__9368\ : InMux
    port map (
            O => \N__41843\,
            I => \N__41837\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__41840\,
            I => \N__41834\
        );

    \I__9366\ : LocalMux
    port map (
            O => \N__41837\,
            I => \N__41829\
        );

    \I__9365\ : Span4Mux_h
    port map (
            O => \N__41834\,
            I => \N__41829\
        );

    \I__9364\ : Odrv4
    port map (
            O => \N__41829\,
            I => \nx.n2395\
        );

    \I__9363\ : InMux
    port map (
            O => \N__41826\,
            I => \N__41823\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__41823\,
            I => \N__41820\
        );

    \I__9361\ : Span4Mux_h
    port map (
            O => \N__41820\,
            I => \N__41817\
        );

    \I__9360\ : Odrv4
    port map (
            O => \N__41817\,
            I => \nx.n2462\
        );

    \I__9359\ : InMux
    port map (
            O => \N__41814\,
            I => \nx.n10741\
        );

    \I__9358\ : CascadeMux
    port map (
            O => \N__41811\,
            I => \N__41808\
        );

    \I__9357\ : InMux
    port map (
            O => \N__41808\,
            I => \N__41805\
        );

    \I__9356\ : LocalMux
    port map (
            O => \N__41805\,
            I => \N__41801\
        );

    \I__9355\ : InMux
    port map (
            O => \N__41804\,
            I => \N__41798\
        );

    \I__9354\ : Span4Mux_v
    port map (
            O => \N__41801\,
            I => \N__41795\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__41798\,
            I => \nx.n2394\
        );

    \I__9352\ : Odrv4
    port map (
            O => \N__41795\,
            I => \nx.n2394\
        );

    \I__9351\ : InMux
    port map (
            O => \N__41790\,
            I => \N__41787\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__41787\,
            I => \N__41784\
        );

    \I__9349\ : Span4Mux_v
    port map (
            O => \N__41784\,
            I => \N__41781\
        );

    \I__9348\ : Span4Mux_h
    port map (
            O => \N__41781\,
            I => \N__41778\
        );

    \I__9347\ : Odrv4
    port map (
            O => \N__41778\,
            I => \nx.n2461\
        );

    \I__9346\ : InMux
    port map (
            O => \N__41775\,
            I => \bfn_14_23_0_\
        );

    \I__9345\ : CascadeMux
    port map (
            O => \N__41772\,
            I => \N__41769\
        );

    \I__9344\ : InMux
    port map (
            O => \N__41769\,
            I => \N__41766\
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__41766\,
            I => \N__41761\
        );

    \I__9342\ : InMux
    port map (
            O => \N__41765\,
            I => \N__41756\
        );

    \I__9341\ : InMux
    port map (
            O => \N__41764\,
            I => \N__41756\
        );

    \I__9340\ : Span4Mux_v
    port map (
            O => \N__41761\,
            I => \N__41753\
        );

    \I__9339\ : LocalMux
    port map (
            O => \N__41756\,
            I => \nx.n2393\
        );

    \I__9338\ : Odrv4
    port map (
            O => \N__41753\,
            I => \nx.n2393\
        );

    \I__9337\ : CascadeMux
    port map (
            O => \N__41748\,
            I => \N__41745\
        );

    \I__9336\ : InMux
    port map (
            O => \N__41745\,
            I => \N__41742\
        );

    \I__9335\ : LocalMux
    port map (
            O => \N__41742\,
            I => \N__41739\
        );

    \I__9334\ : Span4Mux_h
    port map (
            O => \N__41739\,
            I => \N__41736\
        );

    \I__9333\ : Odrv4
    port map (
            O => \N__41736\,
            I => \nx.n2460\
        );

    \I__9332\ : InMux
    port map (
            O => \N__41733\,
            I => \nx.n10743\
        );

    \I__9331\ : CascadeMux
    port map (
            O => \N__41730\,
            I => \N__41727\
        );

    \I__9330\ : InMux
    port map (
            O => \N__41727\,
            I => \N__41724\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__41724\,
            I => \N__41719\
        );

    \I__9328\ : InMux
    port map (
            O => \N__41723\,
            I => \N__41714\
        );

    \I__9327\ : InMux
    port map (
            O => \N__41722\,
            I => \N__41714\
        );

    \I__9326\ : Span4Mux_h
    port map (
            O => \N__41719\,
            I => \N__41711\
        );

    \I__9325\ : LocalMux
    port map (
            O => \N__41714\,
            I => \N__41708\
        );

    \I__9324\ : Odrv4
    port map (
            O => \N__41711\,
            I => \nx.n2392\
        );

    \I__9323\ : Odrv4
    port map (
            O => \N__41708\,
            I => \nx.n2392\
        );

    \I__9322\ : CascadeMux
    port map (
            O => \N__41703\,
            I => \N__41700\
        );

    \I__9321\ : InMux
    port map (
            O => \N__41700\,
            I => \N__41697\
        );

    \I__9320\ : LocalMux
    port map (
            O => \N__41697\,
            I => \N__41694\
        );

    \I__9319\ : Span4Mux_v
    port map (
            O => \N__41694\,
            I => \N__41691\
        );

    \I__9318\ : Odrv4
    port map (
            O => \N__41691\,
            I => \nx.n2459\
        );

    \I__9317\ : InMux
    port map (
            O => \N__41688\,
            I => \nx.n10744\
        );

    \I__9316\ : InMux
    port map (
            O => \N__41685\,
            I => \N__41682\
        );

    \I__9315\ : LocalMux
    port map (
            O => \N__41682\,
            I => \N__41679\
        );

    \I__9314\ : Span4Mux_v
    port map (
            O => \N__41679\,
            I => \N__41676\
        );

    \I__9313\ : Odrv4
    port map (
            O => \N__41676\,
            I => \nx.n2458\
        );

    \I__9312\ : InMux
    port map (
            O => \N__41673\,
            I => \nx.n10745\
        );

    \I__9311\ : CascadeMux
    port map (
            O => \N__41670\,
            I => \N__41666\
        );

    \I__9310\ : InMux
    port map (
            O => \N__41669\,
            I => \N__41657\
        );

    \I__9309\ : InMux
    port map (
            O => \N__41666\,
            I => \N__41654\
        );

    \I__9308\ : CascadeMux
    port map (
            O => \N__41665\,
            I => \N__41650\
        );

    \I__9307\ : CascadeMux
    port map (
            O => \N__41664\,
            I => \N__41647\
        );

    \I__9306\ : CascadeMux
    port map (
            O => \N__41663\,
            I => \N__41644\
        );

    \I__9305\ : CascadeMux
    port map (
            O => \N__41662\,
            I => \N__41641\
        );

    \I__9304\ : CascadeMux
    port map (
            O => \N__41661\,
            I => \N__41637\
        );

    \I__9303\ : InMux
    port map (
            O => \N__41660\,
            I => \N__41632\
        );

    \I__9302\ : LocalMux
    port map (
            O => \N__41657\,
            I => \N__41626\
        );

    \I__9301\ : LocalMux
    port map (
            O => \N__41654\,
            I => \N__41626\
        );

    \I__9300\ : InMux
    port map (
            O => \N__41653\,
            I => \N__41613\
        );

    \I__9299\ : InMux
    port map (
            O => \N__41650\,
            I => \N__41613\
        );

    \I__9298\ : InMux
    port map (
            O => \N__41647\,
            I => \N__41613\
        );

    \I__9297\ : InMux
    port map (
            O => \N__41644\,
            I => \N__41613\
        );

    \I__9296\ : InMux
    port map (
            O => \N__41641\,
            I => \N__41613\
        );

    \I__9295\ : InMux
    port map (
            O => \N__41640\,
            I => \N__41613\
        );

    \I__9294\ : InMux
    port map (
            O => \N__41637\,
            I => \N__41604\
        );

    \I__9293\ : InMux
    port map (
            O => \N__41636\,
            I => \N__41604\
        );

    \I__9292\ : InMux
    port map (
            O => \N__41635\,
            I => \N__41604\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__41632\,
            I => \N__41601\
        );

    \I__9290\ : CascadeMux
    port map (
            O => \N__41631\,
            I => \N__41595\
        );

    \I__9289\ : Span4Mux_v
    port map (
            O => \N__41626\,
            I => \N__41588\
        );

    \I__9288\ : LocalMux
    port map (
            O => \N__41613\,
            I => \N__41588\
        );

    \I__9287\ : InMux
    port map (
            O => \N__41612\,
            I => \N__41585\
        );

    \I__9286\ : InMux
    port map (
            O => \N__41611\,
            I => \N__41582\
        );

    \I__9285\ : LocalMux
    port map (
            O => \N__41604\,
            I => \N__41577\
        );

    \I__9284\ : Span4Mux_v
    port map (
            O => \N__41601\,
            I => \N__41577\
        );

    \I__9283\ : InMux
    port map (
            O => \N__41600\,
            I => \N__41574\
        );

    \I__9282\ : InMux
    port map (
            O => \N__41599\,
            I => \N__41567\
        );

    \I__9281\ : InMux
    port map (
            O => \N__41598\,
            I => \N__41567\
        );

    \I__9280\ : InMux
    port map (
            O => \N__41595\,
            I => \N__41567\
        );

    \I__9279\ : InMux
    port map (
            O => \N__41594\,
            I => \N__41564\
        );

    \I__9278\ : InMux
    port map (
            O => \N__41593\,
            I => \N__41561\
        );

    \I__9277\ : Span4Mux_h
    port map (
            O => \N__41588\,
            I => \N__41558\
        );

    \I__9276\ : LocalMux
    port map (
            O => \N__41585\,
            I => \nx.n2423\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__41582\,
            I => \nx.n2423\
        );

    \I__9274\ : Odrv4
    port map (
            O => \N__41577\,
            I => \nx.n2423\
        );

    \I__9273\ : LocalMux
    port map (
            O => \N__41574\,
            I => \nx.n2423\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__41567\,
            I => \nx.n2423\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__41564\,
            I => \nx.n2423\
        );

    \I__9270\ : LocalMux
    port map (
            O => \N__41561\,
            I => \nx.n2423\
        );

    \I__9269\ : Odrv4
    port map (
            O => \N__41558\,
            I => \nx.n2423\
        );

    \I__9268\ : InMux
    port map (
            O => \N__41541\,
            I => \nx.n10746\
        );

    \I__9267\ : InMux
    port map (
            O => \N__41538\,
            I => \N__41534\
        );

    \I__9266\ : CascadeMux
    port map (
            O => \N__41537\,
            I => \N__41531\
        );

    \I__9265\ : LocalMux
    port map (
            O => \N__41534\,
            I => \N__41528\
        );

    \I__9264\ : InMux
    port map (
            O => \N__41531\,
            I => \N__41525\
        );

    \I__9263\ : Span4Mux_h
    port map (
            O => \N__41528\,
            I => \N__41522\
        );

    \I__9262\ : LocalMux
    port map (
            O => \N__41525\,
            I => \N__41519\
        );

    \I__9261\ : Odrv4
    port map (
            O => \N__41522\,
            I => \nx.n2489\
        );

    \I__9260\ : Odrv4
    port map (
            O => \N__41519\,
            I => \nx.n2489\
        );

    \I__9259\ : InMux
    port map (
            O => \N__41514\,
            I => \N__41510\
        );

    \I__9258\ : CascadeMux
    port map (
            O => \N__41513\,
            I => \N__41507\
        );

    \I__9257\ : LocalMux
    port map (
            O => \N__41510\,
            I => \N__41503\
        );

    \I__9256\ : InMux
    port map (
            O => \N__41507\,
            I => \N__41500\
        );

    \I__9255\ : InMux
    port map (
            O => \N__41506\,
            I => \N__41497\
        );

    \I__9254\ : Span4Mux_h
    port map (
            O => \N__41503\,
            I => \N__41492\
        );

    \I__9253\ : LocalMux
    port map (
            O => \N__41500\,
            I => \N__41492\
        );

    \I__9252\ : LocalMux
    port map (
            O => \N__41497\,
            I => \nx.n2207\
        );

    \I__9251\ : Odrv4
    port map (
            O => \N__41492\,
            I => \nx.n2207\
        );

    \I__9250\ : CascadeMux
    port map (
            O => \N__41487\,
            I => \N__41484\
        );

    \I__9249\ : InMux
    port map (
            O => \N__41484\,
            I => \N__41481\
        );

    \I__9248\ : LocalMux
    port map (
            O => \N__41481\,
            I => \nx.n2274\
        );

    \I__9247\ : CascadeMux
    port map (
            O => \N__41478\,
            I => \N__41474\
        );

    \I__9246\ : InMux
    port map (
            O => \N__41477\,
            I => \N__41468\
        );

    \I__9245\ : InMux
    port map (
            O => \N__41474\,
            I => \N__41468\
        );

    \I__9244\ : CascadeMux
    port map (
            O => \N__41473\,
            I => \N__41465\
        );

    \I__9243\ : LocalMux
    port map (
            O => \N__41468\,
            I => \N__41462\
        );

    \I__9242\ : InMux
    port map (
            O => \N__41465\,
            I => \N__41459\
        );

    \I__9241\ : Span4Mux_h
    port map (
            O => \N__41462\,
            I => \N__41456\
        );

    \I__9240\ : LocalMux
    port map (
            O => \N__41459\,
            I => \nx.n2391\
        );

    \I__9239\ : Odrv4
    port map (
            O => \N__41456\,
            I => \nx.n2391\
        );

    \I__9238\ : InMux
    port map (
            O => \N__41451\,
            I => \N__41448\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__41448\,
            I => \nx.n2470\
        );

    \I__9236\ : InMux
    port map (
            O => \N__41445\,
            I => \nx.n10733\
        );

    \I__9235\ : InMux
    port map (
            O => \N__41442\,
            I => \N__41439\
        );

    \I__9234\ : LocalMux
    port map (
            O => \N__41439\,
            I => \N__41436\
        );

    \I__9233\ : Span4Mux_v
    port map (
            O => \N__41436\,
            I => \N__41433\
        );

    \I__9232\ : Odrv4
    port map (
            O => \N__41433\,
            I => \nx.n2469\
        );

    \I__9231\ : InMux
    port map (
            O => \N__41430\,
            I => \bfn_14_22_0_\
        );

    \I__9230\ : CascadeMux
    port map (
            O => \N__41427\,
            I => \N__41424\
        );

    \I__9229\ : InMux
    port map (
            O => \N__41424\,
            I => \N__41419\
        );

    \I__9228\ : CascadeMux
    port map (
            O => \N__41423\,
            I => \N__41416\
        );

    \I__9227\ : CascadeMux
    port map (
            O => \N__41422\,
            I => \N__41413\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__41419\,
            I => \N__41410\
        );

    \I__9225\ : InMux
    port map (
            O => \N__41416\,
            I => \N__41407\
        );

    \I__9224\ : InMux
    port map (
            O => \N__41413\,
            I => \N__41404\
        );

    \I__9223\ : Span4Mux_h
    port map (
            O => \N__41410\,
            I => \N__41401\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__41407\,
            I => \nx.n2401\
        );

    \I__9221\ : LocalMux
    port map (
            O => \N__41404\,
            I => \nx.n2401\
        );

    \I__9220\ : Odrv4
    port map (
            O => \N__41401\,
            I => \nx.n2401\
        );

    \I__9219\ : InMux
    port map (
            O => \N__41394\,
            I => \N__41391\
        );

    \I__9218\ : LocalMux
    port map (
            O => \N__41391\,
            I => \nx.n2468\
        );

    \I__9217\ : InMux
    port map (
            O => \N__41388\,
            I => \nx.n10735\
        );

    \I__9216\ : InMux
    port map (
            O => \N__41385\,
            I => \N__41382\
        );

    \I__9215\ : LocalMux
    port map (
            O => \N__41382\,
            I => \N__41379\
        );

    \I__9214\ : Span4Mux_h
    port map (
            O => \N__41379\,
            I => \N__41376\
        );

    \I__9213\ : Span4Mux_h
    port map (
            O => \N__41376\,
            I => \N__41373\
        );

    \I__9212\ : Odrv4
    port map (
            O => \N__41373\,
            I => \nx.n2467\
        );

    \I__9211\ : InMux
    port map (
            O => \N__41370\,
            I => \nx.n10736\
        );

    \I__9210\ : CascadeMux
    port map (
            O => \N__41367\,
            I => \N__41363\
        );

    \I__9209\ : InMux
    port map (
            O => \N__41366\,
            I => \N__41359\
        );

    \I__9208\ : InMux
    port map (
            O => \N__41363\,
            I => \N__41356\
        );

    \I__9207\ : InMux
    port map (
            O => \N__41362\,
            I => \N__41353\
        );

    \I__9206\ : LocalMux
    port map (
            O => \N__41359\,
            I => \nx.n2399\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__41356\,
            I => \nx.n2399\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__41353\,
            I => \nx.n2399\
        );

    \I__9203\ : InMux
    port map (
            O => \N__41346\,
            I => \N__41343\
        );

    \I__9202\ : LocalMux
    port map (
            O => \N__41343\,
            I => \N__41340\
        );

    \I__9201\ : Odrv4
    port map (
            O => \N__41340\,
            I => \nx.n2466\
        );

    \I__9200\ : InMux
    port map (
            O => \N__41337\,
            I => \nx.n10737\
        );

    \I__9199\ : CascadeMux
    port map (
            O => \N__41334\,
            I => \N__41331\
        );

    \I__9198\ : InMux
    port map (
            O => \N__41331\,
            I => \N__41328\
        );

    \I__9197\ : LocalMux
    port map (
            O => \N__41328\,
            I => \N__41325\
        );

    \I__9196\ : Span4Mux_v
    port map (
            O => \N__41325\,
            I => \N__41322\
        );

    \I__9195\ : Odrv4
    port map (
            O => \N__41322\,
            I => \nx.n2465\
        );

    \I__9194\ : InMux
    port map (
            O => \N__41319\,
            I => \nx.n10738\
        );

    \I__9193\ : InMux
    port map (
            O => \N__41316\,
            I => \N__41313\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__41313\,
            I => \N__41310\
        );

    \I__9191\ : Span4Mux_h
    port map (
            O => \N__41310\,
            I => \N__41307\
        );

    \I__9190\ : Odrv4
    port map (
            O => \N__41307\,
            I => \nx.n2464\
        );

    \I__9189\ : InMux
    port map (
            O => \N__41304\,
            I => \nx.n10739\
        );

    \I__9188\ : CascadeMux
    port map (
            O => \N__41301\,
            I => \N__41298\
        );

    \I__9187\ : InMux
    port map (
            O => \N__41298\,
            I => \N__41295\
        );

    \I__9186\ : LocalMux
    port map (
            O => \N__41295\,
            I => \N__41292\
        );

    \I__9185\ : Span4Mux_v
    port map (
            O => \N__41292\,
            I => \N__41289\
        );

    \I__9184\ : Odrv4
    port map (
            O => \N__41289\,
            I => \nx.n2463\
        );

    \I__9183\ : InMux
    port map (
            O => \N__41286\,
            I => \nx.n10740\
        );

    \I__9182\ : InMux
    port map (
            O => \N__41283\,
            I => \N__41280\
        );

    \I__9181\ : LocalMux
    port map (
            O => \N__41280\,
            I => \N__41276\
        );

    \I__9180\ : InMux
    port map (
            O => \N__41279\,
            I => \N__41272\
        );

    \I__9179\ : Span4Mux_h
    port map (
            O => \N__41276\,
            I => \N__41269\
        );

    \I__9178\ : InMux
    port map (
            O => \N__41275\,
            I => \N__41265\
        );

    \I__9177\ : LocalMux
    port map (
            O => \N__41272\,
            I => \N__41262\
        );

    \I__9176\ : Span4Mux_v
    port map (
            O => \N__41269\,
            I => \N__41259\
        );

    \I__9175\ : CascadeMux
    port map (
            O => \N__41268\,
            I => \N__41255\
        );

    \I__9174\ : LocalMux
    port map (
            O => \N__41265\,
            I => \N__41252\
        );

    \I__9173\ : Span4Mux_v
    port map (
            O => \N__41262\,
            I => \N__41247\
        );

    \I__9172\ : Span4Mux_h
    port map (
            O => \N__41259\,
            I => \N__41247\
        );

    \I__9171\ : InMux
    port map (
            O => \N__41258\,
            I => \N__41244\
        );

    \I__9170\ : InMux
    port map (
            O => \N__41255\,
            I => \N__41241\
        );

    \I__9169\ : Span12Mux_v
    port map (
            O => \N__41252\,
            I => \N__41238\
        );

    \I__9168\ : Span4Mux_h
    port map (
            O => \N__41247\,
            I => \N__41235\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__41244\,
            I => \nx.bit_ctr_11\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__41241\,
            I => \nx.bit_ctr_11\
        );

    \I__9165\ : Odrv12
    port map (
            O => \N__41238\,
            I => \nx.bit_ctr_11\
        );

    \I__9164\ : Odrv4
    port map (
            O => \N__41235\,
            I => \nx.bit_ctr_11\
        );

    \I__9163\ : InMux
    port map (
            O => \N__41226\,
            I => \N__41223\
        );

    \I__9162\ : LocalMux
    port map (
            O => \N__41223\,
            I => \N__41220\
        );

    \I__9161\ : Sp12to4
    port map (
            O => \N__41220\,
            I => \N__41217\
        );

    \I__9160\ : Span12Mux_s11_v
    port map (
            O => \N__41217\,
            I => \N__41214\
        );

    \I__9159\ : Odrv12
    port map (
            O => \N__41214\,
            I => \nx.n2477\
        );

    \I__9158\ : InMux
    port map (
            O => \N__41211\,
            I => \bfn_14_21_0_\
        );

    \I__9157\ : CascadeMux
    port map (
            O => \N__41208\,
            I => \N__41205\
        );

    \I__9156\ : InMux
    port map (
            O => \N__41205\,
            I => \N__41200\
        );

    \I__9155\ : CascadeMux
    port map (
            O => \N__41204\,
            I => \N__41197\
        );

    \I__9154\ : CascadeMux
    port map (
            O => \N__41203\,
            I => \N__41194\
        );

    \I__9153\ : LocalMux
    port map (
            O => \N__41200\,
            I => \N__41191\
        );

    \I__9152\ : InMux
    port map (
            O => \N__41197\,
            I => \N__41188\
        );

    \I__9151\ : InMux
    port map (
            O => \N__41194\,
            I => \N__41185\
        );

    \I__9150\ : Span4Mux_h
    port map (
            O => \N__41191\,
            I => \N__41182\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__41188\,
            I => \N__41179\
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__41185\,
            I => \N__41176\
        );

    \I__9147\ : Span4Mux_h
    port map (
            O => \N__41182\,
            I => \N__41173\
        );

    \I__9146\ : Span4Mux_h
    port map (
            O => \N__41179\,
            I => \N__41170\
        );

    \I__9145\ : Odrv12
    port map (
            O => \N__41176\,
            I => \nx.n2409\
        );

    \I__9144\ : Odrv4
    port map (
            O => \N__41173\,
            I => \nx.n2409\
        );

    \I__9143\ : Odrv4
    port map (
            O => \N__41170\,
            I => \nx.n2409\
        );

    \I__9142\ : InMux
    port map (
            O => \N__41163\,
            I => \N__41160\
        );

    \I__9141\ : LocalMux
    port map (
            O => \N__41160\,
            I => \nx.n2476\
        );

    \I__9140\ : InMux
    port map (
            O => \N__41157\,
            I => \nx.n10727\
        );

    \I__9139\ : CascadeMux
    port map (
            O => \N__41154\,
            I => \N__41150\
        );

    \I__9138\ : InMux
    port map (
            O => \N__41153\,
            I => \N__41147\
        );

    \I__9137\ : InMux
    port map (
            O => \N__41150\,
            I => \N__41143\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__41147\,
            I => \N__41140\
        );

    \I__9135\ : CascadeMux
    port map (
            O => \N__41146\,
            I => \N__41137\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__41143\,
            I => \N__41132\
        );

    \I__9133\ : Span4Mux_h
    port map (
            O => \N__41140\,
            I => \N__41132\
        );

    \I__9132\ : InMux
    port map (
            O => \N__41137\,
            I => \N__41129\
        );

    \I__9131\ : Odrv4
    port map (
            O => \N__41132\,
            I => \nx.n2408\
        );

    \I__9130\ : LocalMux
    port map (
            O => \N__41129\,
            I => \nx.n2408\
        );

    \I__9129\ : InMux
    port map (
            O => \N__41124\,
            I => \N__41121\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__41121\,
            I => \N__41118\
        );

    \I__9127\ : Span4Mux_h
    port map (
            O => \N__41118\,
            I => \N__41115\
        );

    \I__9126\ : Odrv4
    port map (
            O => \N__41115\,
            I => \nx.n2475\
        );

    \I__9125\ : InMux
    port map (
            O => \N__41112\,
            I => \nx.n10728\
        );

    \I__9124\ : InMux
    port map (
            O => \N__41109\,
            I => \N__41105\
        );

    \I__9123\ : CascadeMux
    port map (
            O => \N__41108\,
            I => \N__41101\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__41105\,
            I => \N__41098\
        );

    \I__9121\ : InMux
    port map (
            O => \N__41104\,
            I => \N__41095\
        );

    \I__9120\ : InMux
    port map (
            O => \N__41101\,
            I => \N__41092\
        );

    \I__9119\ : Odrv4
    port map (
            O => \N__41098\,
            I => \nx.n2407\
        );

    \I__9118\ : LocalMux
    port map (
            O => \N__41095\,
            I => \nx.n2407\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__41092\,
            I => \nx.n2407\
        );

    \I__9116\ : InMux
    port map (
            O => \N__41085\,
            I => \N__41082\
        );

    \I__9115\ : LocalMux
    port map (
            O => \N__41082\,
            I => \nx.n2474\
        );

    \I__9114\ : InMux
    port map (
            O => \N__41079\,
            I => \nx.n10729\
        );

    \I__9113\ : InMux
    port map (
            O => \N__41076\,
            I => \N__41073\
        );

    \I__9112\ : LocalMux
    port map (
            O => \N__41073\,
            I => \N__41070\
        );

    \I__9111\ : Span4Mux_h
    port map (
            O => \N__41070\,
            I => \N__41067\
        );

    \I__9110\ : Odrv4
    port map (
            O => \N__41067\,
            I => \nx.n2473\
        );

    \I__9109\ : InMux
    port map (
            O => \N__41064\,
            I => \nx.n10730\
        );

    \I__9108\ : InMux
    port map (
            O => \N__41061\,
            I => \N__41056\
        );

    \I__9107\ : InMux
    port map (
            O => \N__41060\,
            I => \N__41053\
        );

    \I__9106\ : CascadeMux
    port map (
            O => \N__41059\,
            I => \N__41050\
        );

    \I__9105\ : LocalMux
    port map (
            O => \N__41056\,
            I => \N__41047\
        );

    \I__9104\ : LocalMux
    port map (
            O => \N__41053\,
            I => \N__41044\
        );

    \I__9103\ : InMux
    port map (
            O => \N__41050\,
            I => \N__41041\
        );

    \I__9102\ : Span4Mux_v
    port map (
            O => \N__41047\,
            I => \N__41036\
        );

    \I__9101\ : Span4Mux_h
    port map (
            O => \N__41044\,
            I => \N__41036\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__41041\,
            I => \nx.n2405\
        );

    \I__9099\ : Odrv4
    port map (
            O => \N__41036\,
            I => \nx.n2405\
        );

    \I__9098\ : CascadeMux
    port map (
            O => \N__41031\,
            I => \N__41028\
        );

    \I__9097\ : InMux
    port map (
            O => \N__41028\,
            I => \N__41025\
        );

    \I__9096\ : LocalMux
    port map (
            O => \N__41025\,
            I => \N__41022\
        );

    \I__9095\ : Span4Mux_h
    port map (
            O => \N__41022\,
            I => \N__41019\
        );

    \I__9094\ : Odrv4
    port map (
            O => \N__41019\,
            I => \nx.n2472\
        );

    \I__9093\ : InMux
    port map (
            O => \N__41016\,
            I => \nx.n10731\
        );

    \I__9092\ : CascadeMux
    port map (
            O => \N__41013\,
            I => \N__41009\
        );

    \I__9091\ : InMux
    port map (
            O => \N__41012\,
            I => \N__41006\
        );

    \I__9090\ : InMux
    port map (
            O => \N__41009\,
            I => \N__41003\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__41006\,
            I => \nx.n2404\
        );

    \I__9088\ : LocalMux
    port map (
            O => \N__41003\,
            I => \nx.n2404\
        );

    \I__9087\ : InMux
    port map (
            O => \N__40998\,
            I => \N__40995\
        );

    \I__9086\ : LocalMux
    port map (
            O => \N__40995\,
            I => \nx.n2471\
        );

    \I__9085\ : InMux
    port map (
            O => \N__40992\,
            I => \nx.n10732\
        );

    \I__9084\ : CascadeMux
    port map (
            O => \N__40989\,
            I => \n13474_cascade_\
        );

    \I__9083\ : CascadeMux
    port map (
            O => \N__40986\,
            I => \N__40982\
        );

    \I__9082\ : InMux
    port map (
            O => \N__40985\,
            I => \N__40979\
        );

    \I__9081\ : InMux
    port map (
            O => \N__40982\,
            I => \N__40976\
        );

    \I__9080\ : LocalMux
    port map (
            O => \N__40979\,
            I => \N__40971\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__40976\,
            I => \N__40971\
        );

    \I__9078\ : Span12Mux_v
    port map (
            O => \N__40971\,
            I => \N__40968\
        );

    \I__9077\ : Span12Mux_v
    port map (
            O => \N__40968\,
            I => \N__40965\
        );

    \I__9076\ : Span12Mux_h
    port map (
            O => \N__40965\,
            I => \N__40962\
        );

    \I__9075\ : Odrv12
    port map (
            O => \N__40962\,
            I => pin_in_12
        );

    \I__9074\ : InMux
    port map (
            O => \N__40959\,
            I => \N__40956\
        );

    \I__9073\ : LocalMux
    port map (
            O => \N__40956\,
            I => n13477
        );

    \I__9072\ : InMux
    port map (
            O => \N__40953\,
            I => \N__40947\
        );

    \I__9071\ : InMux
    port map (
            O => \N__40952\,
            I => \N__40947\
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__40947\,
            I => \N__40944\
        );

    \I__9069\ : Span4Mux_v
    port map (
            O => \N__40944\,
            I => \N__40941\
        );

    \I__9068\ : Sp12to4
    port map (
            O => \N__40941\,
            I => \N__40938\
        );

    \I__9067\ : Span12Mux_h
    port map (
            O => \N__40938\,
            I => \N__40935\
        );

    \I__9066\ : Odrv12
    port map (
            O => \N__40935\,
            I => pin_in_13
        );

    \I__9065\ : CascadeMux
    port map (
            O => \N__40932\,
            I => \N__40929\
        );

    \I__9064\ : InMux
    port map (
            O => \N__40929\,
            I => \N__40923\
        );

    \I__9063\ : InMux
    port map (
            O => \N__40928\,
            I => \N__40923\
        );

    \I__9062\ : LocalMux
    port map (
            O => \N__40923\,
            I => \N__40920\
        );

    \I__9061\ : Span12Mux_v
    port map (
            O => \N__40920\,
            I => \N__40917\
        );

    \I__9060\ : Span12Mux_h
    port map (
            O => \N__40917\,
            I => \N__40914\
        );

    \I__9059\ : Odrv12
    port map (
            O => \N__40914\,
            I => pin_in_15
        );

    \I__9058\ : InMux
    port map (
            O => \N__40911\,
            I => \N__40908\
        );

    \I__9057\ : LocalMux
    port map (
            O => \N__40908\,
            I => n2367
        );

    \I__9056\ : InMux
    port map (
            O => \N__40905\,
            I => \N__40902\
        );

    \I__9055\ : LocalMux
    port map (
            O => \N__40902\,
            I => n33
        );

    \I__9054\ : CascadeMux
    port map (
            O => \N__40899\,
            I => \n2379_cascade_\
        );

    \I__9053\ : InMux
    port map (
            O => \N__40896\,
            I => \N__40893\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__40893\,
            I => n45_adj_772
        );

    \I__9051\ : InMux
    port map (
            O => \N__40890\,
            I => \N__40880\
        );

    \I__9050\ : InMux
    port map (
            O => \N__40889\,
            I => \N__40880\
        );

    \I__9049\ : InMux
    port map (
            O => \N__40888\,
            I => \N__40880\
        );

    \I__9048\ : InMux
    port map (
            O => \N__40887\,
            I => \N__40877\
        );

    \I__9047\ : LocalMux
    port map (
            O => \N__40880\,
            I => \N__40874\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__40877\,
            I => \N__40871\
        );

    \I__9045\ : Span4Mux_h
    port map (
            O => \N__40874\,
            I => \N__40868\
        );

    \I__9044\ : Span4Mux_v
    port map (
            O => \N__40871\,
            I => \N__40865\
        );

    \I__9043\ : Span4Mux_h
    port map (
            O => \N__40868\,
            I => \N__40861\
        );

    \I__9042\ : Span4Mux_v
    port map (
            O => \N__40865\,
            I => \N__40858\
        );

    \I__9041\ : InMux
    port map (
            O => \N__40864\,
            I => \N__40855\
        );

    \I__9040\ : Span4Mux_v
    port map (
            O => \N__40861\,
            I => \N__40852\
        );

    \I__9039\ : Span4Mux_h
    port map (
            O => \N__40858\,
            I => \N__40849\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__40855\,
            I => neopxl_color_4
        );

    \I__9037\ : Odrv4
    port map (
            O => \N__40852\,
            I => neopxl_color_4
        );

    \I__9036\ : Odrv4
    port map (
            O => \N__40849\,
            I => neopxl_color_4
        );

    \I__9035\ : SRMux
    port map (
            O => \N__40842\,
            I => \N__40839\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__40839\,
            I => \N__40836\
        );

    \I__9033\ : Span4Mux_v
    port map (
            O => \N__40836\,
            I => \N__40833\
        );

    \I__9032\ : Span4Mux_h
    port map (
            O => \N__40833\,
            I => \N__40830\
        );

    \I__9031\ : Span4Mux_v
    port map (
            O => \N__40830\,
            I => \N__40827\
        );

    \I__9030\ : Odrv4
    port map (
            O => \N__40827\,
            I => n22_adj_732
        );

    \I__9029\ : CEMux
    port map (
            O => \N__40824\,
            I => \N__40821\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__40821\,
            I => \N__40817\
        );

    \I__9027\ : CEMux
    port map (
            O => \N__40820\,
            I => \N__40814\
        );

    \I__9026\ : Span4Mux_v
    port map (
            O => \N__40817\,
            I => \N__40807\
        );

    \I__9025\ : LocalMux
    port map (
            O => \N__40814\,
            I => \N__40807\
        );

    \I__9024\ : CEMux
    port map (
            O => \N__40813\,
            I => \N__40803\
        );

    \I__9023\ : CEMux
    port map (
            O => \N__40812\,
            I => \N__40800\
        );

    \I__9022\ : Span4Mux_v
    port map (
            O => \N__40807\,
            I => \N__40797\
        );

    \I__9021\ : InMux
    port map (
            O => \N__40806\,
            I => \N__40794\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__40803\,
            I => \N__40789\
        );

    \I__9019\ : LocalMux
    port map (
            O => \N__40800\,
            I => \N__40789\
        );

    \I__9018\ : Span4Mux_h
    port map (
            O => \N__40797\,
            I => \N__40784\
        );

    \I__9017\ : LocalMux
    port map (
            O => \N__40794\,
            I => \N__40784\
        );

    \I__9016\ : Span4Mux_v
    port map (
            O => \N__40789\,
            I => \N__40779\
        );

    \I__9015\ : Span4Mux_v
    port map (
            O => \N__40784\,
            I => \N__40779\
        );

    \I__9014\ : Span4Mux_v
    port map (
            O => \N__40779\,
            I => \N__40776\
        );

    \I__9013\ : Odrv4
    port map (
            O => \N__40776\,
            I => n7232
        );

    \I__9012\ : InMux
    port map (
            O => \N__40773\,
            I => \N__40770\
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__40770\,
            I => \N__40767\
        );

    \I__9010\ : Odrv4
    port map (
            O => \N__40767\,
            I => n43
        );

    \I__9009\ : InMux
    port map (
            O => \N__40764\,
            I => \N__40761\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__40761\,
            I => n52_adj_770
        );

    \I__9007\ : InMux
    port map (
            O => \N__40758\,
            I => \N__40750\
        );

    \I__9006\ : InMux
    port map (
            O => \N__40757\,
            I => \N__40750\
        );

    \I__9005\ : InMux
    port map (
            O => \N__40756\,
            I => \N__40747\
        );

    \I__9004\ : InMux
    port map (
            O => \N__40755\,
            I => \N__40743\
        );

    \I__9003\ : LocalMux
    port map (
            O => \N__40750\,
            I => \N__40740\
        );

    \I__9002\ : LocalMux
    port map (
            O => \N__40747\,
            I => \N__40737\
        );

    \I__9001\ : InMux
    port map (
            O => \N__40746\,
            I => \N__40734\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__40743\,
            I => \N__40729\
        );

    \I__8999\ : Span12Mux_v
    port map (
            O => \N__40740\,
            I => \N__40729\
        );

    \I__8998\ : Span12Mux_s10_h
    port map (
            O => \N__40737\,
            I => \N__40726\
        );

    \I__8997\ : LocalMux
    port map (
            O => \N__40734\,
            I => neopxl_color_6
        );

    \I__8996\ : Odrv12
    port map (
            O => \N__40729\,
            I => neopxl_color_6
        );

    \I__8995\ : Odrv12
    port map (
            O => \N__40726\,
            I => neopxl_color_6
        );

    \I__8994\ : SRMux
    port map (
            O => \N__40719\,
            I => \N__40716\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__40716\,
            I => \N__40713\
        );

    \I__8992\ : Odrv12
    port map (
            O => \N__40713\,
            I => n22_adj_728
        );

    \I__8991\ : CascadeMux
    port map (
            O => \N__40710\,
            I => \n7150_cascade_\
        );

    \I__8990\ : InMux
    port map (
            O => \N__40707\,
            I => \N__40704\
        );

    \I__8989\ : LocalMux
    port map (
            O => \N__40704\,
            I => \N__40700\
        );

    \I__8988\ : InMux
    port map (
            O => \N__40703\,
            I => \N__40697\
        );

    \I__8987\ : Span4Mux_v
    port map (
            O => \N__40700\,
            I => \N__40694\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__40697\,
            I => \N__40691\
        );

    \I__8985\ : Span4Mux_h
    port map (
            O => \N__40694\,
            I => \N__40688\
        );

    \I__8984\ : Span4Mux_v
    port map (
            O => \N__40691\,
            I => \N__40685\
        );

    \I__8983\ : Sp12to4
    port map (
            O => \N__40688\,
            I => \N__40680\
        );

    \I__8982\ : Sp12to4
    port map (
            O => \N__40685\,
            I => \N__40680\
        );

    \I__8981\ : Span12Mux_s11_h
    port map (
            O => \N__40680\,
            I => \N__40677\
        );

    \I__8980\ : Span12Mux_v
    port map (
            O => \N__40677\,
            I => \N__40674\
        );

    \I__8979\ : Odrv12
    port map (
            O => \N__40674\,
            I => pin_in_11
        );

    \I__8978\ : InMux
    port map (
            O => \N__40671\,
            I => \N__40668\
        );

    \I__8977\ : LocalMux
    port map (
            O => \N__40668\,
            I => n2355
        );

    \I__8976\ : CascadeMux
    port map (
            O => \N__40665\,
            I => \N__40661\
        );

    \I__8975\ : InMux
    port map (
            O => \N__40664\,
            I => \N__40658\
        );

    \I__8974\ : InMux
    port map (
            O => \N__40661\,
            I => \N__40652\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__40658\,
            I => \N__40649\
        );

    \I__8972\ : InMux
    port map (
            O => \N__40657\,
            I => \N__40645\
        );

    \I__8971\ : InMux
    port map (
            O => \N__40656\,
            I => \N__40642\
        );

    \I__8970\ : InMux
    port map (
            O => \N__40655\,
            I => \N__40639\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__40652\,
            I => \N__40636\
        );

    \I__8968\ : Span4Mux_h
    port map (
            O => \N__40649\,
            I => \N__40633\
        );

    \I__8967\ : InMux
    port map (
            O => \N__40648\,
            I => \N__40630\
        );

    \I__8966\ : LocalMux
    port map (
            O => \N__40645\,
            I => \N__40627\
        );

    \I__8965\ : LocalMux
    port map (
            O => \N__40642\,
            I => n21_adj_714
        );

    \I__8964\ : LocalMux
    port map (
            O => \N__40639\,
            I => n21_adj_714
        );

    \I__8963\ : Odrv4
    port map (
            O => \N__40636\,
            I => n21_adj_714
        );

    \I__8962\ : Odrv4
    port map (
            O => \N__40633\,
            I => n21_adj_714
        );

    \I__8961\ : LocalMux
    port map (
            O => \N__40630\,
            I => n21_adj_714
        );

    \I__8960\ : Odrv12
    port map (
            O => \N__40627\,
            I => n21_adj_714
        );

    \I__8959\ : CascadeMux
    port map (
            O => \N__40614\,
            I => \n7_adj_719_cascade_\
        );

    \I__8958\ : InMux
    port map (
            O => \N__40611\,
            I => \N__40606\
        );

    \I__8957\ : InMux
    port map (
            O => \N__40610\,
            I => \N__40603\
        );

    \I__8956\ : InMux
    port map (
            O => \N__40609\,
            I => \N__40600\
        );

    \I__8955\ : LocalMux
    port map (
            O => \N__40606\,
            I => n7150
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__40603\,
            I => n7150
        );

    \I__8953\ : LocalMux
    port map (
            O => \N__40600\,
            I => n7150
        );

    \I__8952\ : CascadeMux
    port map (
            O => \N__40593\,
            I => \N__40590\
        );

    \I__8951\ : InMux
    port map (
            O => \N__40590\,
            I => \N__40587\
        );

    \I__8950\ : LocalMux
    port map (
            O => \N__40587\,
            I => \N__40584\
        );

    \I__8949\ : Sp12to4
    port map (
            O => \N__40584\,
            I => \N__40580\
        );

    \I__8948\ : InMux
    port map (
            O => \N__40583\,
            I => \N__40577\
        );

    \I__8947\ : Span12Mux_v
    port map (
            O => \N__40580\,
            I => \N__40572\
        );

    \I__8946\ : LocalMux
    port map (
            O => \N__40577\,
            I => \N__40572\
        );

    \I__8945\ : Span12Mux_h
    port map (
            O => \N__40572\,
            I => \N__40569\
        );

    \I__8944\ : Span12Mux_v
    port map (
            O => \N__40569\,
            I => \N__40566\
        );

    \I__8943\ : Odrv12
    port map (
            O => \N__40566\,
            I => pin_in_9
        );

    \I__8942\ : InMux
    port map (
            O => \N__40563\,
            I => \N__40560\
        );

    \I__8941\ : LocalMux
    port map (
            O => \N__40560\,
            I => n2337
        );

    \I__8940\ : CascadeMux
    port map (
            O => \N__40557\,
            I => \n2343_cascade_\
        );

    \I__8939\ : InMux
    port map (
            O => \N__40554\,
            I => \N__40551\
        );

    \I__8938\ : LocalMux
    port map (
            O => \N__40551\,
            I => n2325
        );

    \I__8937\ : InMux
    port map (
            O => \N__40548\,
            I => \N__40545\
        );

    \I__8936\ : LocalMux
    port map (
            O => \N__40545\,
            I => \N__40541\
        );

    \I__8935\ : InMux
    port map (
            O => \N__40544\,
            I => \N__40538\
        );

    \I__8934\ : Span4Mux_v
    port map (
            O => \N__40541\,
            I => \N__40535\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__40538\,
            I => \N__40532\
        );

    \I__8932\ : Span4Mux_h
    port map (
            O => \N__40535\,
            I => \N__40529\
        );

    \I__8931\ : Span4Mux_v
    port map (
            O => \N__40532\,
            I => \N__40526\
        );

    \I__8930\ : Sp12to4
    port map (
            O => \N__40529\,
            I => \N__40521\
        );

    \I__8929\ : Sp12to4
    port map (
            O => \N__40526\,
            I => \N__40521\
        );

    \I__8928\ : Odrv12
    port map (
            O => \N__40521\,
            I => pin_in_3
        );

    \I__8927\ : CascadeMux
    port map (
            O => \N__40518\,
            I => \N__40514\
        );

    \I__8926\ : InMux
    port map (
            O => \N__40517\,
            I => \N__40511\
        );

    \I__8925\ : InMux
    port map (
            O => \N__40514\,
            I => \N__40508\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__40511\,
            I => \N__40505\
        );

    \I__8923\ : LocalMux
    port map (
            O => \N__40508\,
            I => \N__40502\
        );

    \I__8922\ : Span4Mux_v
    port map (
            O => \N__40505\,
            I => \N__40499\
        );

    \I__8921\ : Span12Mux_h
    port map (
            O => \N__40502\,
            I => \N__40494\
        );

    \I__8920\ : Sp12to4
    port map (
            O => \N__40499\,
            I => \N__40494\
        );

    \I__8919\ : Span12Mux_h
    port map (
            O => \N__40494\,
            I => \N__40491\
        );

    \I__8918\ : Span12Mux_v
    port map (
            O => \N__40491\,
            I => \N__40488\
        );

    \I__8917\ : Odrv12
    port map (
            O => \N__40488\,
            I => pin_in_1
        );

    \I__8916\ : InMux
    port map (
            O => \N__40485\,
            I => \N__40482\
        );

    \I__8915\ : LocalMux
    port map (
            O => \N__40482\,
            I => n2361
        );

    \I__8914\ : InMux
    port map (
            O => \N__40479\,
            I => \N__40475\
        );

    \I__8913\ : InMux
    port map (
            O => \N__40478\,
            I => \N__40472\
        );

    \I__8912\ : LocalMux
    port map (
            O => \N__40475\,
            I => \N__40469\
        );

    \I__8911\ : LocalMux
    port map (
            O => \N__40472\,
            I => \N__40466\
        );

    \I__8910\ : Span12Mux_v
    port map (
            O => \N__40469\,
            I => \N__40463\
        );

    \I__8909\ : Span4Mux_v
    port map (
            O => \N__40466\,
            I => \N__40460\
        );

    \I__8908\ : Span12Mux_h
    port map (
            O => \N__40463\,
            I => \N__40457\
        );

    \I__8907\ : Sp12to4
    port map (
            O => \N__40460\,
            I => \N__40454\
        );

    \I__8906\ : Odrv12
    port map (
            O => \N__40457\,
            I => pin_in_2
        );

    \I__8905\ : Odrv12
    port map (
            O => \N__40454\,
            I => pin_in_2
        );

    \I__8904\ : InMux
    port map (
            O => \N__40449\,
            I => \N__40445\
        );

    \I__8903\ : CascadeMux
    port map (
            O => \N__40448\,
            I => \N__40438\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__40445\,
            I => \N__40435\
        );

    \I__8901\ : InMux
    port map (
            O => \N__40444\,
            I => \N__40432\
        );

    \I__8900\ : InMux
    port map (
            O => \N__40443\,
            I => \N__40429\
        );

    \I__8899\ : InMux
    port map (
            O => \N__40442\,
            I => \N__40426\
        );

    \I__8898\ : InMux
    port map (
            O => \N__40441\,
            I => \N__40423\
        );

    \I__8897\ : InMux
    port map (
            O => \N__40438\,
            I => \N__40420\
        );

    \I__8896\ : Span4Mux_v
    port map (
            O => \N__40435\,
            I => \N__40417\
        );

    \I__8895\ : LocalMux
    port map (
            O => \N__40432\,
            I => n22_adj_740
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__40429\,
            I => n22_adj_740
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__40426\,
            I => n22_adj_740
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__40423\,
            I => n22_adj_740
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__40420\,
            I => n22_adj_740
        );

    \I__8890\ : Odrv4
    port map (
            O => \N__40417\,
            I => n22_adj_740
        );

    \I__8889\ : CascadeMux
    port map (
            O => \N__40404\,
            I => \n21_adj_741_cascade_\
        );

    \I__8888\ : InMux
    port map (
            O => \N__40401\,
            I => \N__40398\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__40398\,
            I => \N__40394\
        );

    \I__8886\ : InMux
    port map (
            O => \N__40397\,
            I => \N__40391\
        );

    \I__8885\ : Span4Mux_v
    port map (
            O => \N__40394\,
            I => \N__40386\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__40391\,
            I => \N__40386\
        );

    \I__8883\ : Odrv4
    port map (
            O => \N__40386\,
            I => n7128
        );

    \I__8882\ : CascadeMux
    port map (
            O => \N__40383\,
            I => \N__40380\
        );

    \I__8881\ : InMux
    port map (
            O => \N__40380\,
            I => \N__40377\
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__40377\,
            I => \N__40373\
        );

    \I__8879\ : InMux
    port map (
            O => \N__40376\,
            I => \N__40370\
        );

    \I__8878\ : Odrv4
    port map (
            O => \N__40373\,
            I => \nx.n2192\
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__40370\,
            I => \nx.n2192\
        );

    \I__8876\ : InMux
    port map (
            O => \N__40365\,
            I => \nx.n10707\
        );

    \I__8875\ : CascadeMux
    port map (
            O => \N__40362\,
            I => \N__40358\
        );

    \I__8874\ : InMux
    port map (
            O => \N__40361\,
            I => \N__40355\
        );

    \I__8873\ : InMux
    port map (
            O => \N__40358\,
            I => \N__40348\
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__40355\,
            I => \N__40343\
        );

    \I__8871\ : InMux
    port map (
            O => \N__40354\,
            I => \N__40338\
        );

    \I__8870\ : InMux
    port map (
            O => \N__40353\,
            I => \N__40338\
        );

    \I__8869\ : InMux
    port map (
            O => \N__40352\,
            I => \N__40335\
        );

    \I__8868\ : InMux
    port map (
            O => \N__40351\,
            I => \N__40331\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__40348\,
            I => \N__40328\
        );

    \I__8866\ : InMux
    port map (
            O => \N__40347\,
            I => \N__40323\
        );

    \I__8865\ : InMux
    port map (
            O => \N__40346\,
            I => \N__40323\
        );

    \I__8864\ : Span4Mux_v
    port map (
            O => \N__40343\,
            I => \N__40320\
        );

    \I__8863\ : LocalMux
    port map (
            O => \N__40338\,
            I => \N__40317\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__40335\,
            I => \N__40314\
        );

    \I__8861\ : InMux
    port map (
            O => \N__40334\,
            I => \N__40311\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__40331\,
            I => n7155
        );

    \I__8859\ : Odrv4
    port map (
            O => \N__40328\,
            I => n7155
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__40323\,
            I => n7155
        );

    \I__8857\ : Odrv4
    port map (
            O => \N__40320\,
            I => n7155
        );

    \I__8856\ : Odrv4
    port map (
            O => \N__40317\,
            I => n7155
        );

    \I__8855\ : Odrv4
    port map (
            O => \N__40314\,
            I => n7155
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__40311\,
            I => n7155
        );

    \I__8853\ : InMux
    port map (
            O => \N__40296\,
            I => \N__40293\
        );

    \I__8852\ : LocalMux
    port map (
            O => \N__40293\,
            I => n6166
        );

    \I__8851\ : CascadeMux
    port map (
            O => \N__40290\,
            I => \n6166_cascade_\
        );

    \I__8850\ : InMux
    port map (
            O => \N__40287\,
            I => \N__40284\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__40284\,
            I => n7286
        );

    \I__8848\ : CascadeMux
    port map (
            O => \N__40281\,
            I => \n7_adj_753_cascade_\
        );

    \I__8847\ : InMux
    port map (
            O => \N__40278\,
            I => \N__40274\
        );

    \I__8846\ : CascadeMux
    port map (
            O => \N__40277\,
            I => \N__40270\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__40274\,
            I => \N__40267\
        );

    \I__8844\ : InMux
    port map (
            O => \N__40273\,
            I => \N__40264\
        );

    \I__8843\ : InMux
    port map (
            O => \N__40270\,
            I => \N__40261\
        );

    \I__8842\ : Span4Mux_v
    port map (
            O => \N__40267\,
            I => \N__40254\
        );

    \I__8841\ : LocalMux
    port map (
            O => \N__40264\,
            I => \N__40254\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__40261\,
            I => \N__40254\
        );

    \I__8839\ : Odrv4
    port map (
            O => \N__40254\,
            I => \nx.n2201\
        );

    \I__8838\ : InMux
    port map (
            O => \N__40251\,
            I => \N__40248\
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__40248\,
            I => \N__40245\
        );

    \I__8836\ : Odrv4
    port map (
            O => \N__40245\,
            I => \nx.n2268\
        );

    \I__8835\ : InMux
    port map (
            O => \N__40242\,
            I => \nx.n10698\
        );

    \I__8834\ : InMux
    port map (
            O => \N__40239\,
            I => \nx.n10699\
        );

    \I__8833\ : InMux
    port map (
            O => \N__40236\,
            I => \nx.n10700\
        );

    \I__8832\ : InMux
    port map (
            O => \N__40233\,
            I => \nx.n10701\
        );

    \I__8831\ : CascadeMux
    port map (
            O => \N__40230\,
            I => \N__40225\
        );

    \I__8830\ : InMux
    port map (
            O => \N__40229\,
            I => \N__40222\
        );

    \I__8829\ : InMux
    port map (
            O => \N__40228\,
            I => \N__40217\
        );

    \I__8828\ : InMux
    port map (
            O => \N__40225\,
            I => \N__40217\
        );

    \I__8827\ : LocalMux
    port map (
            O => \N__40222\,
            I => \N__40214\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__40217\,
            I => \N__40211\
        );

    \I__8825\ : Odrv4
    port map (
            O => \N__40214\,
            I => \nx.n2197\
        );

    \I__8824\ : Odrv4
    port map (
            O => \N__40211\,
            I => \nx.n2197\
        );

    \I__8823\ : InMux
    port map (
            O => \N__40206\,
            I => \N__40203\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__40203\,
            I => \N__40200\
        );

    \I__8821\ : Span4Mux_v
    port map (
            O => \N__40200\,
            I => \N__40197\
        );

    \I__8820\ : Odrv4
    port map (
            O => \N__40197\,
            I => \nx.n2264\
        );

    \I__8819\ : InMux
    port map (
            O => \N__40194\,
            I => \nx.n10702\
        );

    \I__8818\ : InMux
    port map (
            O => \N__40191\,
            I => \N__40186\
        );

    \I__8817\ : InMux
    port map (
            O => \N__40190\,
            I => \N__40183\
        );

    \I__8816\ : InMux
    port map (
            O => \N__40189\,
            I => \N__40180\
        );

    \I__8815\ : LocalMux
    port map (
            O => \N__40186\,
            I => \N__40177\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__40183\,
            I => \N__40172\
        );

    \I__8813\ : LocalMux
    port map (
            O => \N__40180\,
            I => \N__40172\
        );

    \I__8812\ : Odrv4
    port map (
            O => \N__40177\,
            I => \nx.n2196\
        );

    \I__8811\ : Odrv4
    port map (
            O => \N__40172\,
            I => \nx.n2196\
        );

    \I__8810\ : InMux
    port map (
            O => \N__40167\,
            I => \N__40164\
        );

    \I__8809\ : LocalMux
    port map (
            O => \N__40164\,
            I => \N__40161\
        );

    \I__8808\ : Span4Mux_h
    port map (
            O => \N__40161\,
            I => \N__40158\
        );

    \I__8807\ : Odrv4
    port map (
            O => \N__40158\,
            I => \nx.n2263\
        );

    \I__8806\ : InMux
    port map (
            O => \N__40155\,
            I => \nx.n10703\
        );

    \I__8805\ : CascadeMux
    port map (
            O => \N__40152\,
            I => \N__40148\
        );

    \I__8804\ : InMux
    port map (
            O => \N__40151\,
            I => \N__40145\
        );

    \I__8803\ : InMux
    port map (
            O => \N__40148\,
            I => \N__40142\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__40145\,
            I => \N__40138\
        );

    \I__8801\ : LocalMux
    port map (
            O => \N__40142\,
            I => \N__40135\
        );

    \I__8800\ : InMux
    port map (
            O => \N__40141\,
            I => \N__40132\
        );

    \I__8799\ : Odrv4
    port map (
            O => \N__40138\,
            I => \nx.n2195\
        );

    \I__8798\ : Odrv4
    port map (
            O => \N__40135\,
            I => \nx.n2195\
        );

    \I__8797\ : LocalMux
    port map (
            O => \N__40132\,
            I => \nx.n2195\
        );

    \I__8796\ : CascadeMux
    port map (
            O => \N__40125\,
            I => \N__40122\
        );

    \I__8795\ : InMux
    port map (
            O => \N__40122\,
            I => \N__40119\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__40119\,
            I => \N__40116\
        );

    \I__8793\ : Span4Mux_h
    port map (
            O => \N__40116\,
            I => \N__40113\
        );

    \I__8792\ : Odrv4
    port map (
            O => \N__40113\,
            I => \nx.n2262\
        );

    \I__8791\ : InMux
    port map (
            O => \N__40110\,
            I => \nx.n10704\
        );

    \I__8790\ : CascadeMux
    port map (
            O => \N__40107\,
            I => \N__40103\
        );

    \I__8789\ : CascadeMux
    port map (
            O => \N__40106\,
            I => \N__40100\
        );

    \I__8788\ : InMux
    port map (
            O => \N__40103\,
            I => \N__40097\
        );

    \I__8787\ : InMux
    port map (
            O => \N__40100\,
            I => \N__40094\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__40097\,
            I => \N__40091\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__40094\,
            I => \N__40085\
        );

    \I__8784\ : Span4Mux_h
    port map (
            O => \N__40091\,
            I => \N__40085\
        );

    \I__8783\ : InMux
    port map (
            O => \N__40090\,
            I => \N__40082\
        );

    \I__8782\ : Odrv4
    port map (
            O => \N__40085\,
            I => \nx.n2194\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__40082\,
            I => \nx.n2194\
        );

    \I__8780\ : InMux
    port map (
            O => \N__40077\,
            I => \N__40074\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__40074\,
            I => \N__40071\
        );

    \I__8778\ : Span4Mux_h
    port map (
            O => \N__40071\,
            I => \N__40068\
        );

    \I__8777\ : Odrv4
    port map (
            O => \N__40068\,
            I => \nx.n2261\
        );

    \I__8776\ : InMux
    port map (
            O => \N__40065\,
            I => \bfn_13_25_0_\
        );

    \I__8775\ : InMux
    port map (
            O => \N__40062\,
            I => \nx.n10706\
        );

    \I__8774\ : CascadeMux
    port map (
            O => \N__40059\,
            I => \N__40054\
        );

    \I__8773\ : InMux
    port map (
            O => \N__40058\,
            I => \N__40051\
        );

    \I__8772\ : InMux
    port map (
            O => \N__40057\,
            I => \N__40048\
        );

    \I__8771\ : InMux
    port map (
            O => \N__40054\,
            I => \N__40045\
        );

    \I__8770\ : LocalMux
    port map (
            O => \N__40051\,
            I => \N__40042\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__40048\,
            I => \nx.n2209\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__40045\,
            I => \nx.n2209\
        );

    \I__8767\ : Odrv4
    port map (
            O => \N__40042\,
            I => \nx.n2209\
        );

    \I__8766\ : CascadeMux
    port map (
            O => \N__40035\,
            I => \N__40032\
        );

    \I__8765\ : InMux
    port map (
            O => \N__40032\,
            I => \N__40029\
        );

    \I__8764\ : LocalMux
    port map (
            O => \N__40029\,
            I => \nx.n2276\
        );

    \I__8763\ : InMux
    port map (
            O => \N__40026\,
            I => \nx.n10690\
        );

    \I__8762\ : CascadeMux
    port map (
            O => \N__40023\,
            I => \N__40019\
        );

    \I__8761\ : InMux
    port map (
            O => \N__40022\,
            I => \N__40015\
        );

    \I__8760\ : InMux
    port map (
            O => \N__40019\,
            I => \N__40012\
        );

    \I__8759\ : InMux
    port map (
            O => \N__40018\,
            I => \N__40009\
        );

    \I__8758\ : LocalMux
    port map (
            O => \N__40015\,
            I => \N__40004\
        );

    \I__8757\ : LocalMux
    port map (
            O => \N__40012\,
            I => \N__40004\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__40009\,
            I => \nx.n2208\
        );

    \I__8755\ : Odrv4
    port map (
            O => \N__40004\,
            I => \nx.n2208\
        );

    \I__8754\ : InMux
    port map (
            O => \N__39999\,
            I => \N__39996\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__39996\,
            I => \nx.n2275\
        );

    \I__8752\ : InMux
    port map (
            O => \N__39993\,
            I => \nx.n10691\
        );

    \I__8751\ : InMux
    port map (
            O => \N__39990\,
            I => \nx.n10692\
        );

    \I__8750\ : CascadeMux
    port map (
            O => \N__39987\,
            I => \N__39984\
        );

    \I__8749\ : InMux
    port map (
            O => \N__39984\,
            I => \N__39979\
        );

    \I__8748\ : InMux
    port map (
            O => \N__39983\,
            I => \N__39976\
        );

    \I__8747\ : InMux
    port map (
            O => \N__39982\,
            I => \N__39973\
        );

    \I__8746\ : LocalMux
    port map (
            O => \N__39979\,
            I => \N__39970\
        );

    \I__8745\ : LocalMux
    port map (
            O => \N__39976\,
            I => \nx.n2206\
        );

    \I__8744\ : LocalMux
    port map (
            O => \N__39973\,
            I => \nx.n2206\
        );

    \I__8743\ : Odrv4
    port map (
            O => \N__39970\,
            I => \nx.n2206\
        );

    \I__8742\ : InMux
    port map (
            O => \N__39963\,
            I => \N__39960\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__39960\,
            I => \nx.n2273\
        );

    \I__8740\ : InMux
    port map (
            O => \N__39957\,
            I => \nx.n10693\
        );

    \I__8739\ : CascadeMux
    port map (
            O => \N__39954\,
            I => \N__39951\
        );

    \I__8738\ : InMux
    port map (
            O => \N__39951\,
            I => \N__39946\
        );

    \I__8737\ : InMux
    port map (
            O => \N__39950\,
            I => \N__39941\
        );

    \I__8736\ : InMux
    port map (
            O => \N__39949\,
            I => \N__39941\
        );

    \I__8735\ : LocalMux
    port map (
            O => \N__39946\,
            I => \N__39938\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__39941\,
            I => \nx.n2205\
        );

    \I__8733\ : Odrv4
    port map (
            O => \N__39938\,
            I => \nx.n2205\
        );

    \I__8732\ : CascadeMux
    port map (
            O => \N__39933\,
            I => \N__39930\
        );

    \I__8731\ : InMux
    port map (
            O => \N__39930\,
            I => \N__39927\
        );

    \I__8730\ : LocalMux
    port map (
            O => \N__39927\,
            I => \nx.n2272\
        );

    \I__8729\ : InMux
    port map (
            O => \N__39924\,
            I => \nx.n10694\
        );

    \I__8728\ : InMux
    port map (
            O => \N__39921\,
            I => \nx.n10695\
        );

    \I__8727\ : CascadeMux
    port map (
            O => \N__39918\,
            I => \N__39915\
        );

    \I__8726\ : InMux
    port map (
            O => \N__39915\,
            I => \N__39912\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__39912\,
            I => \N__39907\
        );

    \I__8724\ : InMux
    port map (
            O => \N__39911\,
            I => \N__39904\
        );

    \I__8723\ : InMux
    port map (
            O => \N__39910\,
            I => \N__39901\
        );

    \I__8722\ : Span4Mux_v
    port map (
            O => \N__39907\,
            I => \N__39896\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__39904\,
            I => \N__39896\
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__39901\,
            I => \nx.n2203\
        );

    \I__8719\ : Odrv4
    port map (
            O => \N__39896\,
            I => \nx.n2203\
        );

    \I__8718\ : InMux
    port map (
            O => \N__39891\,
            I => \N__39888\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__39888\,
            I => \nx.n2270\
        );

    \I__8716\ : InMux
    port map (
            O => \N__39885\,
            I => \nx.n10696\
        );

    \I__8715\ : InMux
    port map (
            O => \N__39882\,
            I => \bfn_13_24_0_\
        );

    \I__8714\ : CascadeMux
    port map (
            O => \N__39879\,
            I => \nx.n2300_cascade_\
        );

    \I__8713\ : InMux
    port map (
            O => \N__39876\,
            I => \N__39873\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__39873\,
            I => \nx.n33_adj_644\
        );

    \I__8711\ : InMux
    port map (
            O => \N__39870\,
            I => \N__39867\
        );

    \I__8710\ : LocalMux
    port map (
            O => \N__39867\,
            I => \nx.n34_adj_641\
        );

    \I__8709\ : CascadeMux
    port map (
            O => \N__39864\,
            I => \nx.n32_cascade_\
        );

    \I__8708\ : CascadeMux
    port map (
            O => \N__39861\,
            I => \nx.n2324_cascade_\
        );

    \I__8707\ : InMux
    port map (
            O => \N__39858\,
            I => \N__39853\
        );

    \I__8706\ : InMux
    port map (
            O => \N__39857\,
            I => \N__39850\
        );

    \I__8705\ : InMux
    port map (
            O => \N__39856\,
            I => \N__39847\
        );

    \I__8704\ : LocalMux
    port map (
            O => \N__39853\,
            I => \N__39843\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__39850\,
            I => \N__39838\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__39847\,
            I => \N__39838\
        );

    \I__8701\ : CascadeMux
    port map (
            O => \N__39846\,
            I => \N__39835\
        );

    \I__8700\ : Span4Mux_v
    port map (
            O => \N__39843\,
            I => \N__39832\
        );

    \I__8699\ : Span4Mux_v
    port map (
            O => \N__39838\,
            I => \N__39829\
        );

    \I__8698\ : InMux
    port map (
            O => \N__39835\,
            I => \N__39825\
        );

    \I__8697\ : Span4Mux_h
    port map (
            O => \N__39832\,
            I => \N__39820\
        );

    \I__8696\ : Span4Mux_h
    port map (
            O => \N__39829\,
            I => \N__39820\
        );

    \I__8695\ : InMux
    port map (
            O => \N__39828\,
            I => \N__39817\
        );

    \I__8694\ : LocalMux
    port map (
            O => \N__39825\,
            I => \N__39814\
        );

    \I__8693\ : Span4Mux_h
    port map (
            O => \N__39820\,
            I => \N__39811\
        );

    \I__8692\ : LocalMux
    port map (
            O => \N__39817\,
            I => \nx.bit_ctr_13\
        );

    \I__8691\ : Odrv4
    port map (
            O => \N__39814\,
            I => \nx.bit_ctr_13\
        );

    \I__8690\ : Odrv4
    port map (
            O => \N__39811\,
            I => \nx.bit_ctr_13\
        );

    \I__8689\ : InMux
    port map (
            O => \N__39804\,
            I => \N__39801\
        );

    \I__8688\ : LocalMux
    port map (
            O => \N__39801\,
            I => \nx.n2277\
        );

    \I__8687\ : InMux
    port map (
            O => \N__39798\,
            I => \bfn_13_23_0_\
        );

    \I__8686\ : InMux
    port map (
            O => \N__39795\,
            I => \N__39790\
        );

    \I__8685\ : InMux
    port map (
            O => \N__39794\,
            I => \N__39787\
        );

    \I__8684\ : InMux
    port map (
            O => \N__39793\,
            I => \N__39784\
        );

    \I__8683\ : LocalMux
    port map (
            O => \N__39790\,
            I => \N__39779\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__39787\,
            I => \N__39779\
        );

    \I__8681\ : LocalMux
    port map (
            O => \N__39784\,
            I => \N__39774\
        );

    \I__8680\ : Span4Mux_v
    port map (
            O => \N__39779\,
            I => \N__39771\
        );

    \I__8679\ : InMux
    port map (
            O => \N__39778\,
            I => \N__39768\
        );

    \I__8678\ : InMux
    port map (
            O => \N__39777\,
            I => \N__39765\
        );

    \I__8677\ : Span4Mux_h
    port map (
            O => \N__39774\,
            I => \N__39760\
        );

    \I__8676\ : Span4Mux_h
    port map (
            O => \N__39771\,
            I => \N__39760\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__39768\,
            I => \N__39757\
        );

    \I__8674\ : LocalMux
    port map (
            O => \N__39765\,
            I => \N__39752\
        );

    \I__8673\ : Span4Mux_h
    port map (
            O => \N__39760\,
            I => \N__39752\
        );

    \I__8672\ : Span4Mux_v
    port map (
            O => \N__39757\,
            I => \N__39749\
        );

    \I__8671\ : Odrv4
    port map (
            O => \N__39752\,
            I => neopxl_color_5
        );

    \I__8670\ : Odrv4
    port map (
            O => \N__39749\,
            I => neopxl_color_5
        );

    \I__8669\ : SRMux
    port map (
            O => \N__39744\,
            I => \N__39741\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__39741\,
            I => \N__39738\
        );

    \I__8667\ : Span4Mux_h
    port map (
            O => \N__39738\,
            I => \N__39735\
        );

    \I__8666\ : Span4Mux_h
    port map (
            O => \N__39735\,
            I => \N__39732\
        );

    \I__8665\ : Odrv4
    port map (
            O => \N__39732\,
            I => n22_adj_730
        );

    \I__8664\ : InMux
    port map (
            O => \N__39729\,
            I => \N__39725\
        );

    \I__8663\ : CascadeMux
    port map (
            O => \N__39728\,
            I => \N__39721\
        );

    \I__8662\ : LocalMux
    port map (
            O => \N__39725\,
            I => \N__39718\
        );

    \I__8661\ : InMux
    port map (
            O => \N__39724\,
            I => \N__39715\
        );

    \I__8660\ : InMux
    port map (
            O => \N__39721\,
            I => \N__39712\
        );

    \I__8659\ : Odrv4
    port map (
            O => \N__39718\,
            I => \nx.n2498\
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__39715\,
            I => \nx.n2498\
        );

    \I__8657\ : LocalMux
    port map (
            O => \N__39712\,
            I => \nx.n2498\
        );

    \I__8656\ : CascadeMux
    port map (
            O => \N__39705\,
            I => \nx.n2404_cascade_\
        );

    \I__8655\ : InMux
    port map (
            O => \N__39702\,
            I => \N__39699\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__39699\,
            I => \N__39696\
        );

    \I__8653\ : Odrv4
    port map (
            O => \N__39696\,
            I => \nx.n34_adj_657\
        );

    \I__8652\ : CascadeMux
    port map (
            O => \N__39693\,
            I => \N__39690\
        );

    \I__8651\ : InMux
    port map (
            O => \N__39690\,
            I => \N__39687\
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__39687\,
            I => \N__39682\
        );

    \I__8649\ : InMux
    port map (
            O => \N__39686\,
            I => \N__39679\
        );

    \I__8648\ : InMux
    port map (
            O => \N__39685\,
            I => \N__39676\
        );

    \I__8647\ : Span4Mux_v
    port map (
            O => \N__39682\,
            I => \N__39673\
        );

    \I__8646\ : LocalMux
    port map (
            O => \N__39679\,
            I => \N__39670\
        );

    \I__8645\ : LocalMux
    port map (
            O => \N__39676\,
            I => \nx.n2490\
        );

    \I__8644\ : Odrv4
    port map (
            O => \N__39673\,
            I => \nx.n2490\
        );

    \I__8643\ : Odrv4
    port map (
            O => \N__39670\,
            I => \nx.n2490\
        );

    \I__8642\ : InMux
    port map (
            O => \N__39663\,
            I => \N__39660\
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__39660\,
            I => \N__39656\
        );

    \I__8640\ : CascadeMux
    port map (
            O => \N__39659\,
            I => \N__39653\
        );

    \I__8639\ : Span4Mux_h
    port map (
            O => \N__39656\,
            I => \N__39650\
        );

    \I__8638\ : InMux
    port map (
            O => \N__39653\,
            I => \N__39647\
        );

    \I__8637\ : Odrv4
    port map (
            O => \N__39650\,
            I => \nx.n2504\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__39647\,
            I => \nx.n2504\
        );

    \I__8635\ : CascadeMux
    port map (
            O => \N__39642\,
            I => \nx.n22_adj_637_cascade_\
        );

    \I__8634\ : InMux
    port map (
            O => \N__39639\,
            I => \N__39634\
        );

    \I__8633\ : CascadeMux
    port map (
            O => \N__39638\,
            I => \N__39631\
        );

    \I__8632\ : InMux
    port map (
            O => \N__39637\,
            I => \N__39628\
        );

    \I__8631\ : LocalMux
    port map (
            O => \N__39634\,
            I => \N__39625\
        );

    \I__8630\ : InMux
    port map (
            O => \N__39631\,
            I => \N__39622\
        );

    \I__8629\ : LocalMux
    port map (
            O => \N__39628\,
            I => \N__39619\
        );

    \I__8628\ : Span4Mux_v
    port map (
            O => \N__39625\,
            I => \N__39616\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__39622\,
            I => \N__39613\
        );

    \I__8626\ : Odrv4
    port map (
            O => \N__39619\,
            I => \nx.n2507\
        );

    \I__8625\ : Odrv4
    port map (
            O => \N__39616\,
            I => \nx.n2507\
        );

    \I__8624\ : Odrv4
    port map (
            O => \N__39613\,
            I => \nx.n2507\
        );

    \I__8623\ : InMux
    port map (
            O => \N__39606\,
            I => \N__39603\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__39603\,
            I => \N__39600\
        );

    \I__8621\ : Odrv4
    port map (
            O => \N__39600\,
            I => \nx.n37_adj_638\
        );

    \I__8620\ : InMux
    port map (
            O => \N__39597\,
            I => \N__39594\
        );

    \I__8619\ : LocalMux
    port map (
            O => \N__39594\,
            I => \N__39590\
        );

    \I__8618\ : CascadeMux
    port map (
            O => \N__39593\,
            I => \N__39587\
        );

    \I__8617\ : Span4Mux_h
    port map (
            O => \N__39590\,
            I => \N__39583\
        );

    \I__8616\ : InMux
    port map (
            O => \N__39587\,
            I => \N__39580\
        );

    \I__8615\ : InMux
    port map (
            O => \N__39586\,
            I => \N__39577\
        );

    \I__8614\ : Odrv4
    port map (
            O => \N__39583\,
            I => \nx.n2500\
        );

    \I__8613\ : LocalMux
    port map (
            O => \N__39580\,
            I => \nx.n2500\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__39577\,
            I => \nx.n2500\
        );

    \I__8611\ : InMux
    port map (
            O => \N__39570\,
            I => \N__39567\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__39567\,
            I => \N__39564\
        );

    \I__8609\ : Odrv4
    port map (
            O => \N__39564\,
            I => n13483
        );

    \I__8608\ : InMux
    port map (
            O => \N__39561\,
            I => \N__39558\
        );

    \I__8607\ : LocalMux
    port map (
            O => \N__39558\,
            I => n13360
        );

    \I__8606\ : InMux
    port map (
            O => \N__39555\,
            I => \N__39552\
        );

    \I__8605\ : LocalMux
    port map (
            O => \N__39552\,
            I => \nx.n2575\
        );

    \I__8604\ : CascadeMux
    port map (
            O => \N__39549\,
            I => \N__39545\
        );

    \I__8603\ : CascadeMux
    port map (
            O => \N__39548\,
            I => \N__39541\
        );

    \I__8602\ : InMux
    port map (
            O => \N__39545\,
            I => \N__39533\
        );

    \I__8601\ : InMux
    port map (
            O => \N__39544\,
            I => \N__39530\
        );

    \I__8600\ : InMux
    port map (
            O => \N__39541\,
            I => \N__39527\
        );

    \I__8599\ : CascadeMux
    port map (
            O => \N__39540\,
            I => \N__39520\
        );

    \I__8598\ : CascadeMux
    port map (
            O => \N__39539\,
            I => \N__39514\
        );

    \I__8597\ : CascadeMux
    port map (
            O => \N__39538\,
            I => \N__39510\
        );

    \I__8596\ : CascadeMux
    port map (
            O => \N__39537\,
            I => \N__39504\
        );

    \I__8595\ : CascadeMux
    port map (
            O => \N__39536\,
            I => \N__39500\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__39533\,
            I => \N__39496\
        );

    \I__8593\ : LocalMux
    port map (
            O => \N__39530\,
            I => \N__39491\
        );

    \I__8592\ : LocalMux
    port map (
            O => \N__39527\,
            I => \N__39491\
        );

    \I__8591\ : InMux
    port map (
            O => \N__39526\,
            I => \N__39488\
        );

    \I__8590\ : InMux
    port map (
            O => \N__39525\,
            I => \N__39483\
        );

    \I__8589\ : InMux
    port map (
            O => \N__39524\,
            I => \N__39483\
        );

    \I__8588\ : InMux
    port map (
            O => \N__39523\,
            I => \N__39474\
        );

    \I__8587\ : InMux
    port map (
            O => \N__39520\,
            I => \N__39474\
        );

    \I__8586\ : InMux
    port map (
            O => \N__39519\,
            I => \N__39474\
        );

    \I__8585\ : InMux
    port map (
            O => \N__39518\,
            I => \N__39474\
        );

    \I__8584\ : InMux
    port map (
            O => \N__39517\,
            I => \N__39463\
        );

    \I__8583\ : InMux
    port map (
            O => \N__39514\,
            I => \N__39463\
        );

    \I__8582\ : InMux
    port map (
            O => \N__39513\,
            I => \N__39463\
        );

    \I__8581\ : InMux
    port map (
            O => \N__39510\,
            I => \N__39463\
        );

    \I__8580\ : InMux
    port map (
            O => \N__39509\,
            I => \N__39463\
        );

    \I__8579\ : InMux
    port map (
            O => \N__39508\,
            I => \N__39460\
        );

    \I__8578\ : InMux
    port map (
            O => \N__39507\,
            I => \N__39457\
        );

    \I__8577\ : InMux
    port map (
            O => \N__39504\,
            I => \N__39448\
        );

    \I__8576\ : InMux
    port map (
            O => \N__39503\,
            I => \N__39448\
        );

    \I__8575\ : InMux
    port map (
            O => \N__39500\,
            I => \N__39448\
        );

    \I__8574\ : InMux
    port map (
            O => \N__39499\,
            I => \N__39448\
        );

    \I__8573\ : Span4Mux_v
    port map (
            O => \N__39496\,
            I => \N__39443\
        );

    \I__8572\ : Span4Mux_v
    port map (
            O => \N__39491\,
            I => \N__39443\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__39488\,
            I => \N__39440\
        );

    \I__8570\ : LocalMux
    port map (
            O => \N__39483\,
            I => \nx.n2522\
        );

    \I__8569\ : LocalMux
    port map (
            O => \N__39474\,
            I => \nx.n2522\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__39463\,
            I => \nx.n2522\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__39460\,
            I => \nx.n2522\
        );

    \I__8566\ : LocalMux
    port map (
            O => \N__39457\,
            I => \nx.n2522\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__39448\,
            I => \nx.n2522\
        );

    \I__8564\ : Odrv4
    port map (
            O => \N__39443\,
            I => \nx.n2522\
        );

    \I__8563\ : Odrv4
    port map (
            O => \N__39440\,
            I => \nx.n2522\
        );

    \I__8562\ : InMux
    port map (
            O => \N__39423\,
            I => \N__39419\
        );

    \I__8561\ : CascadeMux
    port map (
            O => \N__39422\,
            I => \N__39416\
        );

    \I__8560\ : LocalMux
    port map (
            O => \N__39419\,
            I => \N__39413\
        );

    \I__8559\ : InMux
    port map (
            O => \N__39416\,
            I => \N__39409\
        );

    \I__8558\ : Span4Mux_v
    port map (
            O => \N__39413\,
            I => \N__39406\
        );

    \I__8557\ : InMux
    port map (
            O => \N__39412\,
            I => \N__39403\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__39409\,
            I => \N__39400\
        );

    \I__8555\ : Span4Mux_h
    port map (
            O => \N__39406\,
            I => \N__39395\
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__39403\,
            I => \N__39395\
        );

    \I__8553\ : Span4Mux_h
    port map (
            O => \N__39400\,
            I => \N__39392\
        );

    \I__8552\ : Odrv4
    port map (
            O => \N__39395\,
            I => \nx.n2607\
        );

    \I__8551\ : Odrv4
    port map (
            O => \N__39392\,
            I => \nx.n2607\
        );

    \I__8550\ : CascadeMux
    port map (
            O => \N__39387\,
            I => \N__39384\
        );

    \I__8549\ : InMux
    port map (
            O => \N__39384\,
            I => \N__39381\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__39381\,
            I => \N__39377\
        );

    \I__8547\ : CascadeMux
    port map (
            O => \N__39380\,
            I => \N__39373\
        );

    \I__8546\ : Span4Mux_v
    port map (
            O => \N__39377\,
            I => \N__39370\
        );

    \I__8545\ : InMux
    port map (
            O => \N__39376\,
            I => \N__39367\
        );

    \I__8544\ : InMux
    port map (
            O => \N__39373\,
            I => \N__39364\
        );

    \I__8543\ : Odrv4
    port map (
            O => \N__39370\,
            I => \nx.n2495\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__39367\,
            I => \nx.n2495\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__39364\,
            I => \nx.n2495\
        );

    \I__8540\ : CascadeMux
    port map (
            O => \N__39357\,
            I => \N__39354\
        );

    \I__8539\ : InMux
    port map (
            O => \N__39354\,
            I => \N__39351\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__39351\,
            I => \N__39347\
        );

    \I__8537\ : CascadeMux
    port map (
            O => \N__39350\,
            I => \N__39344\
        );

    \I__8536\ : Span4Mux_v
    port map (
            O => \N__39347\,
            I => \N__39341\
        );

    \I__8535\ : InMux
    port map (
            O => \N__39344\,
            I => \N__39338\
        );

    \I__8534\ : Odrv4
    port map (
            O => \N__39341\,
            I => \nx.n2503\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__39338\,
            I => \nx.n2503\
        );

    \I__8532\ : CascadeMux
    port map (
            O => \N__39333\,
            I => \nx.n2503_cascade_\
        );

    \I__8531\ : InMux
    port map (
            O => \N__39330\,
            I => \N__39327\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__39327\,
            I => \nx.n36_adj_636\
        );

    \I__8529\ : CascadeMux
    port map (
            O => \N__39324\,
            I => \N__39321\
        );

    \I__8528\ : InMux
    port map (
            O => \N__39321\,
            I => \N__39317\
        );

    \I__8527\ : CascadeMux
    port map (
            O => \N__39320\,
            I => \N__39313\
        );

    \I__8526\ : LocalMux
    port map (
            O => \N__39317\,
            I => \N__39310\
        );

    \I__8525\ : InMux
    port map (
            O => \N__39316\,
            I => \N__39307\
        );

    \I__8524\ : InMux
    port map (
            O => \N__39313\,
            I => \N__39304\
        );

    \I__8523\ : Odrv4
    port map (
            O => \N__39310\,
            I => \nx.n2502\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__39307\,
            I => \nx.n2502\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__39304\,
            I => \nx.n2502\
        );

    \I__8520\ : CascadeMux
    port map (
            O => \N__39297\,
            I => \N__39293\
        );

    \I__8519\ : CascadeMux
    port map (
            O => \N__39296\,
            I => \N__39289\
        );

    \I__8518\ : InMux
    port map (
            O => \N__39293\,
            I => \N__39286\
        );

    \I__8517\ : InMux
    port map (
            O => \N__39292\,
            I => \N__39283\
        );

    \I__8516\ : InMux
    port map (
            O => \N__39289\,
            I => \N__39280\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__39286\,
            I => \nx.n2508\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__39283\,
            I => \nx.n2508\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__39280\,
            I => \nx.n2508\
        );

    \I__8512\ : CascadeMux
    port map (
            O => \N__39273\,
            I => \N__39269\
        );

    \I__8511\ : CascadeMux
    port map (
            O => \N__39272\,
            I => \N__39265\
        );

    \I__8510\ : InMux
    port map (
            O => \N__39269\,
            I => \N__39262\
        );

    \I__8509\ : InMux
    port map (
            O => \N__39268\,
            I => \N__39259\
        );

    \I__8508\ : InMux
    port map (
            O => \N__39265\,
            I => \N__39256\
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__39262\,
            I => \nx.n2506\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__39259\,
            I => \nx.n2506\
        );

    \I__8505\ : LocalMux
    port map (
            O => \N__39256\,
            I => \nx.n2506\
        );

    \I__8504\ : InMux
    port map (
            O => \N__39249\,
            I => \N__39243\
        );

    \I__8503\ : InMux
    port map (
            O => \N__39248\,
            I => \N__39243\
        );

    \I__8502\ : LocalMux
    port map (
            O => \N__39243\,
            I => \N__39240\
        );

    \I__8501\ : Span12Mux_h
    port map (
            O => \N__39240\,
            I => \N__39237\
        );

    \I__8500\ : Span12Mux_v
    port map (
            O => \N__39237\,
            I => \N__39234\
        );

    \I__8499\ : Odrv12
    port map (
            O => \N__39234\,
            I => pin_in_8
        );

    \I__8498\ : CascadeMux
    port map (
            O => \N__39231\,
            I => \n13480_cascade_\
        );

    \I__8497\ : CascadeMux
    port map (
            O => \N__39228\,
            I => \current_pin_7__N_157_cascade_\
        );

    \I__8496\ : InMux
    port map (
            O => \N__39225\,
            I => \N__39222\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__39222\,
            I => \N__39218\
        );

    \I__8494\ : InMux
    port map (
            O => \N__39221\,
            I => \N__39215\
        );

    \I__8493\ : Span4Mux_v
    port map (
            O => \N__39218\,
            I => \N__39212\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__39215\,
            I => \N__39209\
        );

    \I__8491\ : Span4Mux_h
    port map (
            O => \N__39212\,
            I => \N__39204\
        );

    \I__8490\ : Span4Mux_v
    port map (
            O => \N__39209\,
            I => \N__39204\
        );

    \I__8489\ : Span4Mux_h
    port map (
            O => \N__39204\,
            I => \N__39201\
        );

    \I__8488\ : Sp12to4
    port map (
            O => \N__39201\,
            I => \N__39198\
        );

    \I__8487\ : Odrv12
    port map (
            O => \N__39198\,
            I => pin_in_0
        );

    \I__8486\ : InMux
    port map (
            O => \N__39195\,
            I => \N__39191\
        );

    \I__8485\ : CascadeMux
    port map (
            O => \N__39194\,
            I => \N__39188\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__39191\,
            I => \N__39185\
        );

    \I__8483\ : InMux
    port map (
            O => \N__39188\,
            I => \N__39182\
        );

    \I__8482\ : Span4Mux_v
    port map (
            O => \N__39185\,
            I => \N__39179\
        );

    \I__8481\ : LocalMux
    port map (
            O => \N__39182\,
            I => \N__39176\
        );

    \I__8480\ : Span4Mux_v
    port map (
            O => \N__39179\,
            I => \N__39173\
        );

    \I__8479\ : Span4Mux_h
    port map (
            O => \N__39176\,
            I => \N__39170\
        );

    \I__8478\ : Span4Mux_v
    port map (
            O => \N__39173\,
            I => \N__39167\
        );

    \I__8477\ : Sp12to4
    port map (
            O => \N__39170\,
            I => \N__39164\
        );

    \I__8476\ : Sp12to4
    port map (
            O => \N__39167\,
            I => \N__39159\
        );

    \I__8475\ : Span12Mux_v
    port map (
            O => \N__39164\,
            I => \N__39159\
        );

    \I__8474\ : Span12Mux_h
    port map (
            O => \N__39159\,
            I => \N__39156\
        );

    \I__8473\ : Odrv12
    port map (
            O => \N__39156\,
            I => pin_in_10
        );

    \I__8472\ : CascadeMux
    port map (
            O => \N__39153\,
            I => \n2289_cascade_\
        );

    \I__8471\ : CascadeMux
    port map (
            O => \N__39150\,
            I => \N__39146\
        );

    \I__8470\ : InMux
    port map (
            O => \N__39149\,
            I => \N__39143\
        );

    \I__8469\ : InMux
    port map (
            O => \N__39146\,
            I => \N__39140\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__39143\,
            I => \N__39137\
        );

    \I__8467\ : LocalMux
    port map (
            O => \N__39140\,
            I => \N__39134\
        );

    \I__8466\ : Span4Mux_v
    port map (
            O => \N__39137\,
            I => \N__39131\
        );

    \I__8465\ : Span4Mux_h
    port map (
            O => \N__39134\,
            I => \N__39128\
        );

    \I__8464\ : Span4Mux_v
    port map (
            O => \N__39131\,
            I => \N__39125\
        );

    \I__8463\ : Sp12to4
    port map (
            O => \N__39128\,
            I => \N__39122\
        );

    \I__8462\ : Span4Mux_v
    port map (
            O => \N__39125\,
            I => \N__39119\
        );

    \I__8461\ : Span12Mux_v
    port map (
            O => \N__39122\,
            I => \N__39116\
        );

    \I__8460\ : Span4Mux_h
    port map (
            O => \N__39119\,
            I => \N__39113\
        );

    \I__8459\ : Odrv12
    port map (
            O => \N__39116\,
            I => pin_in_6
        );

    \I__8458\ : Odrv4
    port map (
            O => \N__39113\,
            I => pin_in_6
        );

    \I__8457\ : InMux
    port map (
            O => \N__39108\,
            I => \N__39105\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__39105\,
            I => \N__39102\
        );

    \I__8455\ : Span4Mux_h
    port map (
            O => \N__39102\,
            I => \N__39099\
        );

    \I__8454\ : Odrv4
    port map (
            O => \N__39099\,
            I => n13453
        );

    \I__8453\ : CascadeMux
    port map (
            O => \N__39096\,
            I => \n13364_cascade_\
        );

    \I__8452\ : InMux
    port map (
            O => \N__39093\,
            I => \N__39090\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__39090\,
            I => n150
        );

    \I__8450\ : CascadeMux
    port map (
            O => \N__39087\,
            I => \n7155_cascade_\
        );

    \I__8449\ : InMux
    port map (
            O => \N__39084\,
            I => \N__39081\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__39081\,
            I => \N__39078\
        );

    \I__8447\ : Odrv4
    port map (
            O => \N__39078\,
            I => n6190
        );

    \I__8446\ : CascadeMux
    port map (
            O => \N__39075\,
            I => \n6190_cascade_\
        );

    \I__8445\ : InMux
    port map (
            O => \N__39072\,
            I => \N__39069\
        );

    \I__8444\ : LocalMux
    port map (
            O => \N__39069\,
            I => \N__39066\
        );

    \I__8443\ : Odrv4
    port map (
            O => \N__39066\,
            I => n7334
        );

    \I__8442\ : InMux
    port map (
            O => \N__39063\,
            I => \N__39057\
        );

    \I__8441\ : InMux
    port map (
            O => \N__39062\,
            I => \N__39057\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__39057\,
            I => n6170
        );

    \I__8439\ : InMux
    port map (
            O => \N__39054\,
            I => \N__39050\
        );

    \I__8438\ : InMux
    port map (
            O => \N__39053\,
            I => \N__39047\
        );

    \I__8437\ : LocalMux
    port map (
            O => \N__39050\,
            I => n9415
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__39047\,
            I => n9415
        );

    \I__8435\ : InMux
    port map (
            O => \N__39042\,
            I => \N__39038\
        );

    \I__8434\ : InMux
    port map (
            O => \N__39041\,
            I => \N__39035\
        );

    \I__8433\ : LocalMux
    port map (
            O => \N__39038\,
            I => delay_counter_28
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__39035\,
            I => delay_counter_28
        );

    \I__8431\ : InMux
    port map (
            O => \N__39030\,
            I => n10544
        );

    \I__8430\ : InMux
    port map (
            O => \N__39027\,
            I => \N__39023\
        );

    \I__8429\ : InMux
    port map (
            O => \N__39026\,
            I => \N__39020\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__39023\,
            I => delay_counter_29
        );

    \I__8427\ : LocalMux
    port map (
            O => \N__39020\,
            I => delay_counter_29
        );

    \I__8426\ : InMux
    port map (
            O => \N__39015\,
            I => n10545
        );

    \I__8425\ : InMux
    port map (
            O => \N__39012\,
            I => \N__39008\
        );

    \I__8424\ : InMux
    port map (
            O => \N__39011\,
            I => \N__39005\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__39008\,
            I => delay_counter_30
        );

    \I__8422\ : LocalMux
    port map (
            O => \N__39005\,
            I => delay_counter_30
        );

    \I__8421\ : InMux
    port map (
            O => \N__39000\,
            I => n10546
        );

    \I__8420\ : InMux
    port map (
            O => \N__38997\,
            I => n10547
        );

    \I__8419\ : SRMux
    port map (
            O => \N__38994\,
            I => \N__38990\
        );

    \I__8418\ : SRMux
    port map (
            O => \N__38993\,
            I => \N__38986\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__38990\,
            I => \N__38983\
        );

    \I__8416\ : SRMux
    port map (
            O => \N__38989\,
            I => \N__38980\
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__38986\,
            I => \N__38977\
        );

    \I__8414\ : Span4Mux_v
    port map (
            O => \N__38983\,
            I => \N__38973\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__38980\,
            I => \N__38970\
        );

    \I__8412\ : Span4Mux_h
    port map (
            O => \N__38977\,
            I => \N__38967\
        );

    \I__8411\ : SRMux
    port map (
            O => \N__38976\,
            I => \N__38964\
        );

    \I__8410\ : Odrv4
    port map (
            O => \N__38973\,
            I => n7442
        );

    \I__8409\ : Odrv12
    port map (
            O => \N__38970\,
            I => n7442
        );

    \I__8408\ : Odrv4
    port map (
            O => \N__38967\,
            I => n7442
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__38964\,
            I => n7442
        );

    \I__8406\ : CascadeMux
    port map (
            O => \N__38955\,
            I => \n10_adj_779_cascade_\
        );

    \I__8405\ : InMux
    port map (
            O => \N__38952\,
            I => \N__38949\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__38949\,
            I => n10_adj_779
        );

    \I__8403\ : CascadeMux
    port map (
            O => \N__38946\,
            I => \n7290_cascade_\
        );

    \I__8402\ : IoInMux
    port map (
            O => \N__38943\,
            I => \N__38940\
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__38940\,
            I => \N__38937\
        );

    \I__8400\ : Span4Mux_s3_v
    port map (
            O => \N__38937\,
            I => \N__38934\
        );

    \I__8399\ : Span4Mux_h
    port map (
            O => \N__38934\,
            I => \N__38931\
        );

    \I__8398\ : Sp12to4
    port map (
            O => \N__38931\,
            I => \N__38928\
        );

    \I__8397\ : Span12Mux_v
    port map (
            O => \N__38928\,
            I => \N__38923\
        );

    \I__8396\ : InMux
    port map (
            O => \N__38927\,
            I => \N__38920\
        );

    \I__8395\ : InMux
    port map (
            O => \N__38926\,
            I => \N__38917\
        );

    \I__8394\ : Odrv12
    port map (
            O => \N__38923\,
            I => pin_out_10
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__38920\,
            I => pin_out_10
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__38917\,
            I => pin_out_10
        );

    \I__8391\ : InMux
    port map (
            O => \N__38910\,
            I => \N__38907\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__38907\,
            I => \N__38903\
        );

    \I__8389\ : InMux
    port map (
            O => \N__38906\,
            I => \N__38900\
        );

    \I__8388\ : Span4Mux_h
    port map (
            O => \N__38903\,
            I => \N__38897\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__38900\,
            I => \N__38894\
        );

    \I__8386\ : Odrv4
    port map (
            O => \N__38897\,
            I => n7135
        );

    \I__8385\ : Odrv4
    port map (
            O => \N__38894\,
            I => n7135
        );

    \I__8384\ : InMux
    port map (
            O => \N__38889\,
            I => \N__38885\
        );

    \I__8383\ : InMux
    port map (
            O => \N__38888\,
            I => \N__38882\
        );

    \I__8382\ : LocalMux
    port map (
            O => \N__38885\,
            I => \N__38879\
        );

    \I__8381\ : LocalMux
    port map (
            O => \N__38882\,
            I => delay_counter_20
        );

    \I__8380\ : Odrv4
    port map (
            O => \N__38879\,
            I => delay_counter_20
        );

    \I__8379\ : InMux
    port map (
            O => \N__38874\,
            I => n10536
        );

    \I__8378\ : InMux
    port map (
            O => \N__38871\,
            I => \N__38867\
        );

    \I__8377\ : InMux
    port map (
            O => \N__38870\,
            I => \N__38864\
        );

    \I__8376\ : LocalMux
    port map (
            O => \N__38867\,
            I => delay_counter_21
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__38864\,
            I => delay_counter_21
        );

    \I__8374\ : InMux
    port map (
            O => \N__38859\,
            I => n10537
        );

    \I__8373\ : CascadeMux
    port map (
            O => \N__38856\,
            I => \N__38852\
        );

    \I__8372\ : InMux
    port map (
            O => \N__38855\,
            I => \N__38849\
        );

    \I__8371\ : InMux
    port map (
            O => \N__38852\,
            I => \N__38846\
        );

    \I__8370\ : LocalMux
    port map (
            O => \N__38849\,
            I => delay_counter_22
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__38846\,
            I => delay_counter_22
        );

    \I__8368\ : InMux
    port map (
            O => \N__38841\,
            I => n10538
        );

    \I__8367\ : InMux
    port map (
            O => \N__38838\,
            I => \N__38834\
        );

    \I__8366\ : InMux
    port map (
            O => \N__38837\,
            I => \N__38831\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__38834\,
            I => delay_counter_23
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__38831\,
            I => delay_counter_23
        );

    \I__8363\ : InMux
    port map (
            O => \N__38826\,
            I => n10539
        );

    \I__8362\ : InMux
    port map (
            O => \N__38823\,
            I => \N__38819\
        );

    \I__8361\ : InMux
    port map (
            O => \N__38822\,
            I => \N__38816\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__38819\,
            I => delay_counter_24
        );

    \I__8359\ : LocalMux
    port map (
            O => \N__38816\,
            I => delay_counter_24
        );

    \I__8358\ : InMux
    port map (
            O => \N__38811\,
            I => \bfn_12_29_0_\
        );

    \I__8357\ : InMux
    port map (
            O => \N__38808\,
            I => \N__38804\
        );

    \I__8356\ : InMux
    port map (
            O => \N__38807\,
            I => \N__38801\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__38804\,
            I => delay_counter_25
        );

    \I__8354\ : LocalMux
    port map (
            O => \N__38801\,
            I => delay_counter_25
        );

    \I__8353\ : InMux
    port map (
            O => \N__38796\,
            I => n10541
        );

    \I__8352\ : InMux
    port map (
            O => \N__38793\,
            I => \N__38789\
        );

    \I__8351\ : InMux
    port map (
            O => \N__38792\,
            I => \N__38786\
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__38789\,
            I => delay_counter_26
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__38786\,
            I => delay_counter_26
        );

    \I__8348\ : InMux
    port map (
            O => \N__38781\,
            I => n10542
        );

    \I__8347\ : CascadeMux
    port map (
            O => \N__38778\,
            I => \N__38774\
        );

    \I__8346\ : InMux
    port map (
            O => \N__38777\,
            I => \N__38771\
        );

    \I__8345\ : InMux
    port map (
            O => \N__38774\,
            I => \N__38768\
        );

    \I__8344\ : LocalMux
    port map (
            O => \N__38771\,
            I => delay_counter_27
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__38768\,
            I => delay_counter_27
        );

    \I__8342\ : InMux
    port map (
            O => \N__38763\,
            I => n10543
        );

    \I__8341\ : InMux
    port map (
            O => \N__38760\,
            I => \N__38756\
        );

    \I__8340\ : InMux
    port map (
            O => \N__38759\,
            I => \N__38753\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__38756\,
            I => delay_counter_12
        );

    \I__8338\ : LocalMux
    port map (
            O => \N__38753\,
            I => delay_counter_12
        );

    \I__8337\ : InMux
    port map (
            O => \N__38748\,
            I => n10528
        );

    \I__8336\ : InMux
    port map (
            O => \N__38745\,
            I => \N__38741\
        );

    \I__8335\ : InMux
    port map (
            O => \N__38744\,
            I => \N__38738\
        );

    \I__8334\ : LocalMux
    port map (
            O => \N__38741\,
            I => delay_counter_13
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__38738\,
            I => delay_counter_13
        );

    \I__8332\ : InMux
    port map (
            O => \N__38733\,
            I => n10529
        );

    \I__8331\ : InMux
    port map (
            O => \N__38730\,
            I => \N__38726\
        );

    \I__8330\ : InMux
    port map (
            O => \N__38729\,
            I => \N__38723\
        );

    \I__8329\ : LocalMux
    port map (
            O => \N__38726\,
            I => delay_counter_14
        );

    \I__8328\ : LocalMux
    port map (
            O => \N__38723\,
            I => delay_counter_14
        );

    \I__8327\ : InMux
    port map (
            O => \N__38718\,
            I => n10530
        );

    \I__8326\ : CascadeMux
    port map (
            O => \N__38715\,
            I => \N__38712\
        );

    \I__8325\ : InMux
    port map (
            O => \N__38712\,
            I => \N__38709\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__38709\,
            I => \N__38705\
        );

    \I__8323\ : InMux
    port map (
            O => \N__38708\,
            I => \N__38702\
        );

    \I__8322\ : Span4Mux_h
    port map (
            O => \N__38705\,
            I => \N__38699\
        );

    \I__8321\ : LocalMux
    port map (
            O => \N__38702\,
            I => delay_counter_15
        );

    \I__8320\ : Odrv4
    port map (
            O => \N__38699\,
            I => delay_counter_15
        );

    \I__8319\ : InMux
    port map (
            O => \N__38694\,
            I => n10531
        );

    \I__8318\ : InMux
    port map (
            O => \N__38691\,
            I => \N__38687\
        );

    \I__8317\ : InMux
    port map (
            O => \N__38690\,
            I => \N__38684\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__38687\,
            I => \N__38681\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__38684\,
            I => delay_counter_16
        );

    \I__8314\ : Odrv4
    port map (
            O => \N__38681\,
            I => delay_counter_16
        );

    \I__8313\ : InMux
    port map (
            O => \N__38676\,
            I => \bfn_12_28_0_\
        );

    \I__8312\ : InMux
    port map (
            O => \N__38673\,
            I => \N__38670\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__38670\,
            I => \N__38666\
        );

    \I__8310\ : InMux
    port map (
            O => \N__38669\,
            I => \N__38663\
        );

    \I__8309\ : Span4Mux_h
    port map (
            O => \N__38666\,
            I => \N__38660\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__38663\,
            I => delay_counter_17
        );

    \I__8307\ : Odrv4
    port map (
            O => \N__38660\,
            I => delay_counter_17
        );

    \I__8306\ : InMux
    port map (
            O => \N__38655\,
            I => n10533
        );

    \I__8305\ : InMux
    port map (
            O => \N__38652\,
            I => \N__38649\
        );

    \I__8304\ : LocalMux
    port map (
            O => \N__38649\,
            I => \N__38645\
        );

    \I__8303\ : InMux
    port map (
            O => \N__38648\,
            I => \N__38642\
        );

    \I__8302\ : Span4Mux_h
    port map (
            O => \N__38645\,
            I => \N__38639\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__38642\,
            I => delay_counter_18
        );

    \I__8300\ : Odrv4
    port map (
            O => \N__38639\,
            I => delay_counter_18
        );

    \I__8299\ : InMux
    port map (
            O => \N__38634\,
            I => n10534
        );

    \I__8298\ : InMux
    port map (
            O => \N__38631\,
            I => \N__38627\
        );

    \I__8297\ : InMux
    port map (
            O => \N__38630\,
            I => \N__38624\
        );

    \I__8296\ : LocalMux
    port map (
            O => \N__38627\,
            I => \N__38621\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__38624\,
            I => delay_counter_19
        );

    \I__8294\ : Odrv4
    port map (
            O => \N__38621\,
            I => delay_counter_19
        );

    \I__8293\ : InMux
    port map (
            O => \N__38616\,
            I => n10535
        );

    \I__8292\ : InMux
    port map (
            O => \N__38613\,
            I => \N__38609\
        );

    \I__8291\ : InMux
    port map (
            O => \N__38612\,
            I => \N__38606\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__38609\,
            I => delay_counter_3
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__38606\,
            I => delay_counter_3
        );

    \I__8288\ : InMux
    port map (
            O => \N__38601\,
            I => n10519
        );

    \I__8287\ : InMux
    port map (
            O => \N__38598\,
            I => \N__38594\
        );

    \I__8286\ : InMux
    port map (
            O => \N__38597\,
            I => \N__38591\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__38594\,
            I => delay_counter_4
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__38591\,
            I => delay_counter_4
        );

    \I__8283\ : InMux
    port map (
            O => \N__38586\,
            I => n10520
        );

    \I__8282\ : InMux
    port map (
            O => \N__38583\,
            I => \N__38579\
        );

    \I__8281\ : InMux
    port map (
            O => \N__38582\,
            I => \N__38576\
        );

    \I__8280\ : LocalMux
    port map (
            O => \N__38579\,
            I => delay_counter_5
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__38576\,
            I => delay_counter_5
        );

    \I__8278\ : InMux
    port map (
            O => \N__38571\,
            I => n10521
        );

    \I__8277\ : InMux
    port map (
            O => \N__38568\,
            I => \N__38564\
        );

    \I__8276\ : InMux
    port map (
            O => \N__38567\,
            I => \N__38561\
        );

    \I__8275\ : LocalMux
    port map (
            O => \N__38564\,
            I => delay_counter_6
        );

    \I__8274\ : LocalMux
    port map (
            O => \N__38561\,
            I => delay_counter_6
        );

    \I__8273\ : InMux
    port map (
            O => \N__38556\,
            I => n10522
        );

    \I__8272\ : InMux
    port map (
            O => \N__38553\,
            I => \N__38549\
        );

    \I__8271\ : InMux
    port map (
            O => \N__38552\,
            I => \N__38546\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__38549\,
            I => delay_counter_7
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__38546\,
            I => delay_counter_7
        );

    \I__8268\ : InMux
    port map (
            O => \N__38541\,
            I => n10523
        );

    \I__8267\ : InMux
    port map (
            O => \N__38538\,
            I => \N__38534\
        );

    \I__8266\ : InMux
    port map (
            O => \N__38537\,
            I => \N__38531\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__38534\,
            I => delay_counter_8
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__38531\,
            I => delay_counter_8
        );

    \I__8263\ : InMux
    port map (
            O => \N__38526\,
            I => \bfn_12_27_0_\
        );

    \I__8262\ : CascadeMux
    port map (
            O => \N__38523\,
            I => \N__38519\
        );

    \I__8261\ : InMux
    port map (
            O => \N__38522\,
            I => \N__38516\
        );

    \I__8260\ : InMux
    port map (
            O => \N__38519\,
            I => \N__38513\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__38516\,
            I => delay_counter_9
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__38513\,
            I => delay_counter_9
        );

    \I__8257\ : InMux
    port map (
            O => \N__38508\,
            I => n10525
        );

    \I__8256\ : InMux
    port map (
            O => \N__38505\,
            I => \N__38501\
        );

    \I__8255\ : InMux
    port map (
            O => \N__38504\,
            I => \N__38498\
        );

    \I__8254\ : LocalMux
    port map (
            O => \N__38501\,
            I => delay_counter_10
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__38498\,
            I => delay_counter_10
        );

    \I__8252\ : InMux
    port map (
            O => \N__38493\,
            I => n10526
        );

    \I__8251\ : InMux
    port map (
            O => \N__38490\,
            I => \N__38486\
        );

    \I__8250\ : InMux
    port map (
            O => \N__38489\,
            I => \N__38483\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__38486\,
            I => delay_counter_11
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__38483\,
            I => delay_counter_11
        );

    \I__8247\ : InMux
    port map (
            O => \N__38478\,
            I => n10527
        );

    \I__8246\ : CascadeMux
    port map (
            O => \N__38475\,
            I => \N__38472\
        );

    \I__8245\ : InMux
    port map (
            O => \N__38472\,
            I => \N__38469\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__38469\,
            I => \nx.n31\
        );

    \I__8243\ : InMux
    port map (
            O => \N__38466\,
            I => \N__38463\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__38463\,
            I => \nx.n28_adj_601\
        );

    \I__8241\ : InMux
    port map (
            O => \N__38460\,
            I => \N__38457\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__38457\,
            I => \N__38454\
        );

    \I__8239\ : Sp12to4
    port map (
            O => \N__38454\,
            I => \N__38450\
        );

    \I__8238\ : InMux
    port map (
            O => \N__38453\,
            I => \N__38447\
        );

    \I__8237\ : Span12Mux_s10_v
    port map (
            O => \N__38450\,
            I => \N__38442\
        );

    \I__8236\ : LocalMux
    port map (
            O => \N__38447\,
            I => \N__38439\
        );

    \I__8235\ : InMux
    port map (
            O => \N__38446\,
            I => \N__38434\
        );

    \I__8234\ : InMux
    port map (
            O => \N__38445\,
            I => \N__38434\
        );

    \I__8233\ : Odrv12
    port map (
            O => \N__38442\,
            I => neopxl_color_12
        );

    \I__8232\ : Odrv4
    port map (
            O => \N__38439\,
            I => neopxl_color_12
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__38434\,
            I => neopxl_color_12
        );

    \I__8230\ : InMux
    port map (
            O => \N__38427\,
            I => \N__38424\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__38424\,
            I => \N__38421\
        );

    \I__8228\ : Span4Mux_h
    port map (
            O => \N__38421\,
            I => \N__38418\
        );

    \I__8227\ : Span4Mux_h
    port map (
            O => \N__38418\,
            I => \N__38415\
        );

    \I__8226\ : Span4Mux_h
    port map (
            O => \N__38415\,
            I => \N__38412\
        );

    \I__8225\ : Odrv4
    port map (
            O => \N__38412\,
            I => neopxl_color_prev_12
        );

    \I__8224\ : InMux
    port map (
            O => \N__38409\,
            I => \N__38406\
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__38406\,
            I => \nx.n30\
        );

    \I__8222\ : InMux
    port map (
            O => \N__38403\,
            I => \N__38400\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__38400\,
            I => \nx.n22_adj_604\
        );

    \I__8220\ : CascadeMux
    port map (
            O => \N__38397\,
            I => \N__38393\
        );

    \I__8219\ : InMux
    port map (
            O => \N__38396\,
            I => \N__38390\
        );

    \I__8218\ : InMux
    port map (
            O => \N__38393\,
            I => \N__38387\
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__38390\,
            I => delay_counter_0
        );

    \I__8216\ : LocalMux
    port map (
            O => \N__38387\,
            I => delay_counter_0
        );

    \I__8215\ : InMux
    port map (
            O => \N__38382\,
            I => \bfn_12_26_0_\
        );

    \I__8214\ : InMux
    port map (
            O => \N__38379\,
            I => \N__38375\
        );

    \I__8213\ : InMux
    port map (
            O => \N__38378\,
            I => \N__38372\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__38375\,
            I => delay_counter_1
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__38372\,
            I => delay_counter_1
        );

    \I__8210\ : InMux
    port map (
            O => \N__38367\,
            I => n10517
        );

    \I__8209\ : InMux
    port map (
            O => \N__38364\,
            I => \N__38360\
        );

    \I__8208\ : InMux
    port map (
            O => \N__38363\,
            I => \N__38357\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__38360\,
            I => delay_counter_2
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__38357\,
            I => delay_counter_2
        );

    \I__8205\ : InMux
    port map (
            O => \N__38352\,
            I => n10518
        );

    \I__8204\ : InMux
    port map (
            O => \N__38349\,
            I => \N__38346\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__38346\,
            I => \nx.n30_adj_640\
        );

    \I__8202\ : CascadeMux
    port map (
            O => \N__38343\,
            I => \nx.n34_cascade_\
        );

    \I__8201\ : InMux
    port map (
            O => \N__38340\,
            I => \N__38337\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__38337\,
            I => \N__38334\
        );

    \I__8199\ : Odrv4
    port map (
            O => \N__38334\,
            I => \nx.n21\
        );

    \I__8198\ : CascadeMux
    port map (
            O => \N__38331\,
            I => \nx.n2225_cascade_\
        );

    \I__8197\ : InMux
    port map (
            O => \N__38328\,
            I => \N__38325\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__38325\,
            I => \N__38322\
        );

    \I__8195\ : Odrv4
    port map (
            O => \N__38322\,
            I => \nx.n2562\
        );

    \I__8194\ : InMux
    port map (
            O => \N__38319\,
            I => \nx.n10761\
        );

    \I__8193\ : InMux
    port map (
            O => \N__38316\,
            I => \N__38312\
        );

    \I__8192\ : InMux
    port map (
            O => \N__38315\,
            I => \N__38309\
        );

    \I__8191\ : LocalMux
    port map (
            O => \N__38312\,
            I => \nx.n2494\
        );

    \I__8190\ : LocalMux
    port map (
            O => \N__38309\,
            I => \nx.n2494\
        );

    \I__8189\ : InMux
    port map (
            O => \N__38304\,
            I => \N__38301\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__38301\,
            I => \nx.n2561\
        );

    \I__8187\ : InMux
    port map (
            O => \N__38298\,
            I => \bfn_12_22_0_\
        );

    \I__8186\ : InMux
    port map (
            O => \N__38295\,
            I => \N__38292\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__38292\,
            I => \N__38288\
        );

    \I__8184\ : InMux
    port map (
            O => \N__38291\,
            I => \N__38285\
        );

    \I__8183\ : Span4Mux_v
    port map (
            O => \N__38288\,
            I => \N__38279\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__38285\,
            I => \N__38279\
        );

    \I__8181\ : InMux
    port map (
            O => \N__38284\,
            I => \N__38276\
        );

    \I__8180\ : Odrv4
    port map (
            O => \N__38279\,
            I => \nx.n2493\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__38276\,
            I => \nx.n2493\
        );

    \I__8178\ : InMux
    port map (
            O => \N__38271\,
            I => \N__38268\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__38268\,
            I => \N__38265\
        );

    \I__8176\ : Span4Mux_h
    port map (
            O => \N__38265\,
            I => \N__38262\
        );

    \I__8175\ : Odrv4
    port map (
            O => \N__38262\,
            I => \nx.n2560\
        );

    \I__8174\ : InMux
    port map (
            O => \N__38259\,
            I => \nx.n10763\
        );

    \I__8173\ : InMux
    port map (
            O => \N__38256\,
            I => \N__38253\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__38253\,
            I => \N__38249\
        );

    \I__8171\ : InMux
    port map (
            O => \N__38252\,
            I => \N__38245\
        );

    \I__8170\ : Span4Mux_v
    port map (
            O => \N__38249\,
            I => \N__38242\
        );

    \I__8169\ : InMux
    port map (
            O => \N__38248\,
            I => \N__38239\
        );

    \I__8168\ : LocalMux
    port map (
            O => \N__38245\,
            I => \nx.n2492\
        );

    \I__8167\ : Odrv4
    port map (
            O => \N__38242\,
            I => \nx.n2492\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__38239\,
            I => \nx.n2492\
        );

    \I__8165\ : InMux
    port map (
            O => \N__38232\,
            I => \N__38229\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__38229\,
            I => \N__38226\
        );

    \I__8163\ : Odrv4
    port map (
            O => \N__38226\,
            I => \nx.n2559\
        );

    \I__8162\ : InMux
    port map (
            O => \N__38223\,
            I => \nx.n10764\
        );

    \I__8161\ : CascadeMux
    port map (
            O => \N__38220\,
            I => \N__38217\
        );

    \I__8160\ : InMux
    port map (
            O => \N__38217\,
            I => \N__38214\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__38214\,
            I => \N__38210\
        );

    \I__8158\ : InMux
    port map (
            O => \N__38213\,
            I => \N__38207\
        );

    \I__8157\ : Span4Mux_v
    port map (
            O => \N__38210\,
            I => \N__38204\
        );

    \I__8156\ : LocalMux
    port map (
            O => \N__38207\,
            I => \nx.n2491\
        );

    \I__8155\ : Odrv4
    port map (
            O => \N__38204\,
            I => \nx.n2491\
        );

    \I__8154\ : InMux
    port map (
            O => \N__38199\,
            I => \N__38196\
        );

    \I__8153\ : LocalMux
    port map (
            O => \N__38196\,
            I => \N__38193\
        );

    \I__8152\ : Odrv4
    port map (
            O => \N__38193\,
            I => \nx.n2558\
        );

    \I__8151\ : InMux
    port map (
            O => \N__38190\,
            I => \nx.n10765\
        );

    \I__8150\ : CascadeMux
    port map (
            O => \N__38187\,
            I => \N__38184\
        );

    \I__8149\ : InMux
    port map (
            O => \N__38184\,
            I => \N__38181\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__38181\,
            I => \N__38178\
        );

    \I__8147\ : Odrv4
    port map (
            O => \N__38178\,
            I => \nx.n2557\
        );

    \I__8146\ : InMux
    port map (
            O => \N__38175\,
            I => \nx.n10766\
        );

    \I__8145\ : InMux
    port map (
            O => \N__38172\,
            I => \nx.n10767\
        );

    \I__8144\ : InMux
    port map (
            O => \N__38169\,
            I => \N__38165\
        );

    \I__8143\ : InMux
    port map (
            O => \N__38168\,
            I => \N__38162\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__38165\,
            I => \N__38159\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__38162\,
            I => \N__38156\
        );

    \I__8140\ : Span4Mux_v
    port map (
            O => \N__38159\,
            I => \N__38153\
        );

    \I__8139\ : Span4Mux_h
    port map (
            O => \N__38156\,
            I => \N__38150\
        );

    \I__8138\ : Odrv4
    port map (
            O => \N__38153\,
            I => \nx.n2588\
        );

    \I__8137\ : Odrv4
    port map (
            O => \N__38150\,
            I => \nx.n2588\
        );

    \I__8136\ : InMux
    port map (
            O => \N__38145\,
            I => \nx.n10752\
        );

    \I__8135\ : InMux
    port map (
            O => \N__38142\,
            I => \N__38139\
        );

    \I__8134\ : LocalMux
    port map (
            O => \N__38139\,
            I => \nx.n2570\
        );

    \I__8133\ : InMux
    port map (
            O => \N__38136\,
            I => \nx.n10753\
        );

    \I__8132\ : InMux
    port map (
            O => \N__38133\,
            I => \N__38130\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__38130\,
            I => \N__38127\
        );

    \I__8130\ : Odrv4
    port map (
            O => \N__38127\,
            I => \nx.n2569\
        );

    \I__8129\ : InMux
    port map (
            O => \N__38124\,
            I => \bfn_12_21_0_\
        );

    \I__8128\ : InMux
    port map (
            O => \N__38121\,
            I => \N__38115\
        );

    \I__8127\ : InMux
    port map (
            O => \N__38120\,
            I => \N__38115\
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__38115\,
            I => \N__38111\
        );

    \I__8125\ : CascadeMux
    port map (
            O => \N__38114\,
            I => \N__38108\
        );

    \I__8124\ : Span4Mux_h
    port map (
            O => \N__38111\,
            I => \N__38105\
        );

    \I__8123\ : InMux
    port map (
            O => \N__38108\,
            I => \N__38102\
        );

    \I__8122\ : Odrv4
    port map (
            O => \N__38105\,
            I => \nx.n2501\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__38102\,
            I => \nx.n2501\
        );

    \I__8120\ : InMux
    port map (
            O => \N__38097\,
            I => \N__38094\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__38094\,
            I => \N__38091\
        );

    \I__8118\ : Odrv4
    port map (
            O => \N__38091\,
            I => \nx.n2568\
        );

    \I__8117\ : InMux
    port map (
            O => \N__38088\,
            I => \nx.n10755\
        );

    \I__8116\ : InMux
    port map (
            O => \N__38085\,
            I => \N__38082\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__38082\,
            I => \N__38079\
        );

    \I__8114\ : Span4Mux_h
    port map (
            O => \N__38079\,
            I => \N__38076\
        );

    \I__8113\ : Odrv4
    port map (
            O => \N__38076\,
            I => \nx.n2567\
        );

    \I__8112\ : InMux
    port map (
            O => \N__38073\,
            I => \nx.n10756\
        );

    \I__8111\ : CascadeMux
    port map (
            O => \N__38070\,
            I => \N__38067\
        );

    \I__8110\ : InMux
    port map (
            O => \N__38067\,
            I => \N__38062\
        );

    \I__8109\ : CascadeMux
    port map (
            O => \N__38066\,
            I => \N__38059\
        );

    \I__8108\ : InMux
    port map (
            O => \N__38065\,
            I => \N__38056\
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__38062\,
            I => \N__38053\
        );

    \I__8106\ : InMux
    port map (
            O => \N__38059\,
            I => \N__38050\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__38056\,
            I => \N__38047\
        );

    \I__8104\ : Span4Mux_v
    port map (
            O => \N__38053\,
            I => \N__38044\
        );

    \I__8103\ : LocalMux
    port map (
            O => \N__38050\,
            I => \N__38039\
        );

    \I__8102\ : Span4Mux_v
    port map (
            O => \N__38047\,
            I => \N__38039\
        );

    \I__8101\ : Odrv4
    port map (
            O => \N__38044\,
            I => \nx.n2499\
        );

    \I__8100\ : Odrv4
    port map (
            O => \N__38039\,
            I => \nx.n2499\
        );

    \I__8099\ : InMux
    port map (
            O => \N__38034\,
            I => \N__38031\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__38031\,
            I => \N__38028\
        );

    \I__8097\ : Odrv4
    port map (
            O => \N__38028\,
            I => \nx.n2566\
        );

    \I__8096\ : InMux
    port map (
            O => \N__38025\,
            I => \nx.n10757\
        );

    \I__8095\ : CascadeMux
    port map (
            O => \N__38022\,
            I => \N__38019\
        );

    \I__8094\ : InMux
    port map (
            O => \N__38019\,
            I => \N__38016\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__38016\,
            I => \N__38013\
        );

    \I__8092\ : Odrv4
    port map (
            O => \N__38013\,
            I => \nx.n2565\
        );

    \I__8091\ : InMux
    port map (
            O => \N__38010\,
            I => \nx.n10758\
        );

    \I__8090\ : CascadeMux
    port map (
            O => \N__38007\,
            I => \N__38004\
        );

    \I__8089\ : InMux
    port map (
            O => \N__38004\,
            I => \N__38000\
        );

    \I__8088\ : InMux
    port map (
            O => \N__38003\,
            I => \N__37997\
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__38000\,
            I => \N__37994\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__37997\,
            I => \nx.n2497\
        );

    \I__8085\ : Odrv4
    port map (
            O => \N__37994\,
            I => \nx.n2497\
        );

    \I__8084\ : InMux
    port map (
            O => \N__37989\,
            I => \N__37986\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__37986\,
            I => \N__37983\
        );

    \I__8082\ : Span4Mux_h
    port map (
            O => \N__37983\,
            I => \N__37980\
        );

    \I__8081\ : Odrv4
    port map (
            O => \N__37980\,
            I => \nx.n2564\
        );

    \I__8080\ : InMux
    port map (
            O => \N__37977\,
            I => \nx.n10759\
        );

    \I__8079\ : InMux
    port map (
            O => \N__37974\,
            I => \N__37969\
        );

    \I__8078\ : CascadeMux
    port map (
            O => \N__37973\,
            I => \N__37966\
        );

    \I__8077\ : InMux
    port map (
            O => \N__37972\,
            I => \N__37963\
        );

    \I__8076\ : LocalMux
    port map (
            O => \N__37969\,
            I => \N__37960\
        );

    \I__8075\ : InMux
    port map (
            O => \N__37966\,
            I => \N__37957\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__37963\,
            I => \N__37950\
        );

    \I__8073\ : Span4Mux_v
    port map (
            O => \N__37960\,
            I => \N__37950\
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__37957\,
            I => \N__37950\
        );

    \I__8071\ : Odrv4
    port map (
            O => \N__37950\,
            I => \nx.n2496\
        );

    \I__8070\ : CascadeMux
    port map (
            O => \N__37947\,
            I => \N__37944\
        );

    \I__8069\ : InMux
    port map (
            O => \N__37944\,
            I => \N__37941\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__37941\,
            I => \N__37938\
        );

    \I__8067\ : Odrv4
    port map (
            O => \N__37938\,
            I => \nx.n2563\
        );

    \I__8066\ : InMux
    port map (
            O => \N__37935\,
            I => \nx.n10760\
        );

    \I__8065\ : CascadeMux
    port map (
            O => \N__37932\,
            I => \N__37929\
        );

    \I__8064\ : InMux
    port map (
            O => \N__37929\,
            I => \N__37925\
        );

    \I__8063\ : InMux
    port map (
            O => \N__37928\,
            I => \N__37922\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__37925\,
            I => \N__37918\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__37922\,
            I => \N__37915\
        );

    \I__8060\ : InMux
    port map (
            O => \N__37921\,
            I => \N__37912\
        );

    \I__8059\ : Span4Mux_h
    port map (
            O => \N__37918\,
            I => \N__37909\
        );

    \I__8058\ : Odrv4
    port map (
            O => \N__37915\,
            I => \nx.n2605\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__37912\,
            I => \nx.n2605\
        );

    \I__8056\ : Odrv4
    port map (
            O => \N__37909\,
            I => \nx.n2605\
        );

    \I__8055\ : InMux
    port map (
            O => \N__37902\,
            I => \N__37899\
        );

    \I__8054\ : LocalMux
    port map (
            O => \N__37899\,
            I => \nx.n35_adj_639\
        );

    \I__8053\ : InMux
    port map (
            O => \N__37896\,
            I => \N__37893\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__37893\,
            I => \N__37888\
        );

    \I__8051\ : InMux
    port map (
            O => \N__37892\,
            I => \N__37885\
        );

    \I__8050\ : InMux
    port map (
            O => \N__37891\,
            I => \N__37882\
        );

    \I__8049\ : Span4Mux_h
    port map (
            O => \N__37888\,
            I => \N__37878\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__37885\,
            I => \N__37875\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__37882\,
            I => \N__37872\
        );

    \I__8046\ : InMux
    port map (
            O => \N__37881\,
            I => \N__37869\
        );

    \I__8045\ : Span4Mux_v
    port map (
            O => \N__37878\,
            I => \N__37866\
        );

    \I__8044\ : Span4Mux_h
    port map (
            O => \N__37875\,
            I => \N__37863\
        );

    \I__8043\ : Span4Mux_h
    port map (
            O => \N__37872\,
            I => \N__37860\
        );

    \I__8042\ : LocalMux
    port map (
            O => \N__37869\,
            I => \N__37854\
        );

    \I__8041\ : Span4Mux_v
    port map (
            O => \N__37866\,
            I => \N__37854\
        );

    \I__8040\ : Sp12to4
    port map (
            O => \N__37863\,
            I => \N__37849\
        );

    \I__8039\ : Sp12to4
    port map (
            O => \N__37860\,
            I => \N__37849\
        );

    \I__8038\ : InMux
    port map (
            O => \N__37859\,
            I => \N__37846\
        );

    \I__8037\ : Span4Mux_h
    port map (
            O => \N__37854\,
            I => \N__37843\
        );

    \I__8036\ : Span12Mux_v
    port map (
            O => \N__37849\,
            I => \N__37840\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__37846\,
            I => \nx.bit_ctr_10\
        );

    \I__8034\ : Odrv4
    port map (
            O => \N__37843\,
            I => \nx.bit_ctr_10\
        );

    \I__8033\ : Odrv12
    port map (
            O => \N__37840\,
            I => \nx.bit_ctr_10\
        );

    \I__8032\ : InMux
    port map (
            O => \N__37833\,
            I => \N__37830\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__37830\,
            I => \N__37827\
        );

    \I__8030\ : Odrv4
    port map (
            O => \N__37827\,
            I => \nx.n2577\
        );

    \I__8029\ : InMux
    port map (
            O => \N__37824\,
            I => \bfn_12_20_0_\
        );

    \I__8028\ : InMux
    port map (
            O => \N__37821\,
            I => \N__37816\
        );

    \I__8027\ : InMux
    port map (
            O => \N__37820\,
            I => \N__37813\
        );

    \I__8026\ : CascadeMux
    port map (
            O => \N__37819\,
            I => \N__37810\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__37816\,
            I => \N__37807\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__37813\,
            I => \N__37804\
        );

    \I__8023\ : InMux
    port map (
            O => \N__37810\,
            I => \N__37801\
        );

    \I__8022\ : Span4Mux_h
    port map (
            O => \N__37807\,
            I => \N__37798\
        );

    \I__8021\ : Span4Mux_v
    port map (
            O => \N__37804\,
            I => \N__37793\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__37801\,
            I => \N__37793\
        );

    \I__8019\ : Odrv4
    port map (
            O => \N__37798\,
            I => \nx.n2509\
        );

    \I__8018\ : Odrv4
    port map (
            O => \N__37793\,
            I => \nx.n2509\
        );

    \I__8017\ : InMux
    port map (
            O => \N__37788\,
            I => \N__37785\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__37785\,
            I => \N__37782\
        );

    \I__8015\ : Odrv4
    port map (
            O => \N__37782\,
            I => \nx.n2576\
        );

    \I__8014\ : InMux
    port map (
            O => \N__37779\,
            I => \nx.n10747\
        );

    \I__8013\ : InMux
    port map (
            O => \N__37776\,
            I => \nx.n10748\
        );

    \I__8012\ : InMux
    port map (
            O => \N__37773\,
            I => \N__37770\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__37770\,
            I => \nx.n2574\
        );

    \I__8010\ : InMux
    port map (
            O => \N__37767\,
            I => \nx.n10749\
        );

    \I__8009\ : InMux
    port map (
            O => \N__37764\,
            I => \N__37761\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__37761\,
            I => \nx.n2573\
        );

    \I__8007\ : InMux
    port map (
            O => \N__37758\,
            I => \nx.n10750\
        );

    \I__8006\ : CascadeMux
    port map (
            O => \N__37755\,
            I => \N__37751\
        );

    \I__8005\ : InMux
    port map (
            O => \N__37754\,
            I => \N__37748\
        );

    \I__8004\ : InMux
    port map (
            O => \N__37751\,
            I => \N__37745\
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__37748\,
            I => \N__37739\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__37745\,
            I => \N__37739\
        );

    \I__8001\ : CascadeMux
    port map (
            O => \N__37744\,
            I => \N__37736\
        );

    \I__8000\ : Span4Mux_v
    port map (
            O => \N__37739\,
            I => \N__37733\
        );

    \I__7999\ : InMux
    port map (
            O => \N__37736\,
            I => \N__37730\
        );

    \I__7998\ : Odrv4
    port map (
            O => \N__37733\,
            I => \nx.n2505\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__37730\,
            I => \nx.n2505\
        );

    \I__7996\ : CascadeMux
    port map (
            O => \N__37725\,
            I => \N__37722\
        );

    \I__7995\ : InMux
    port map (
            O => \N__37722\,
            I => \N__37719\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__37719\,
            I => \N__37716\
        );

    \I__7993\ : Odrv4
    port map (
            O => \N__37716\,
            I => \nx.n2572\
        );

    \I__7992\ : InMux
    port map (
            O => \N__37713\,
            I => \nx.n10751\
        );

    \I__7991\ : InMux
    port map (
            O => \N__37710\,
            I => \N__37707\
        );

    \I__7990\ : LocalMux
    port map (
            O => \N__37707\,
            I => \nx.n2571\
        );

    \I__7989\ : CascadeMux
    port map (
            O => \N__37704\,
            I => \N__37701\
        );

    \I__7988\ : InMux
    port map (
            O => \N__37701\,
            I => \N__37698\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__37698\,
            I => \N__37695\
        );

    \I__7986\ : Span4Mux_v
    port map (
            O => \N__37695\,
            I => \N__37691\
        );

    \I__7985\ : CascadeMux
    port map (
            O => \N__37694\,
            I => \N__37688\
        );

    \I__7984\ : Span4Mux_h
    port map (
            O => \N__37691\,
            I => \N__37685\
        );

    \I__7983\ : InMux
    port map (
            O => \N__37688\,
            I => \N__37682\
        );

    \I__7982\ : Span4Mux_v
    port map (
            O => \N__37685\,
            I => \N__37676\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__37682\,
            I => \N__37676\
        );

    \I__7980\ : InMux
    port map (
            O => \N__37681\,
            I => \N__37673\
        );

    \I__7979\ : Odrv4
    port map (
            O => \N__37676\,
            I => \nx.n2597\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__37673\,
            I => \nx.n2597\
        );

    \I__7977\ : InMux
    port map (
            O => \N__37668\,
            I => \N__37664\
        );

    \I__7976\ : CascadeMux
    port map (
            O => \N__37667\,
            I => \N__37661\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__37664\,
            I => \N__37657\
        );

    \I__7974\ : InMux
    port map (
            O => \N__37661\,
            I => \N__37654\
        );

    \I__7973\ : InMux
    port map (
            O => \N__37660\,
            I => \N__37651\
        );

    \I__7972\ : Span4Mux_h
    port map (
            O => \N__37657\,
            I => \N__37646\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__37654\,
            I => \N__37646\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__37651\,
            I => \nx.n2601\
        );

    \I__7969\ : Odrv4
    port map (
            O => \N__37646\,
            I => \nx.n2601\
        );

    \I__7968\ : CascadeMux
    port map (
            O => \N__37641\,
            I => \nx.n2497_cascade_\
        );

    \I__7967\ : CascadeMux
    port map (
            O => \N__37638\,
            I => \nx.n26_adj_611_cascade_\
        );

    \I__7966\ : InMux
    port map (
            O => \N__37635\,
            I => \N__37632\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__37632\,
            I => \N__37629\
        );

    \I__7964\ : Span4Mux_h
    port map (
            O => \N__37629\,
            I => \N__37626\
        );

    \I__7963\ : Odrv4
    port map (
            O => \N__37626\,
            I => \nx.n33\
        );

    \I__7962\ : CascadeMux
    port map (
            O => \N__37623\,
            I => \nx.n38_adj_612_cascade_\
        );

    \I__7961\ : CascadeMux
    port map (
            O => \N__37620\,
            I => \nx.n2522_cascade_\
        );

    \I__7960\ : CascadeMux
    port map (
            O => \N__37617\,
            I => \N__37612\
        );

    \I__7959\ : InMux
    port map (
            O => \N__37616\,
            I => \N__37607\
        );

    \I__7958\ : InMux
    port map (
            O => \N__37615\,
            I => \N__37607\
        );

    \I__7957\ : InMux
    port map (
            O => \N__37612\,
            I => \N__37604\
        );

    \I__7956\ : LocalMux
    port map (
            O => \N__37607\,
            I => \N__37601\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__37604\,
            I => \N__37598\
        );

    \I__7954\ : Span4Mux_v
    port map (
            O => \N__37601\,
            I => \N__37595\
        );

    \I__7953\ : Span4Mux_h
    port map (
            O => \N__37598\,
            I => \N__37592\
        );

    \I__7952\ : Odrv4
    port map (
            O => \N__37595\,
            I => \nx.n2600\
        );

    \I__7951\ : Odrv4
    port map (
            O => \N__37592\,
            I => \nx.n2600\
        );

    \I__7950\ : CascadeMux
    port map (
            O => \N__37587\,
            I => \n7166_cascade_\
        );

    \I__7949\ : CascadeMux
    port map (
            O => \N__37584\,
            I => \N__37580\
        );

    \I__7948\ : InMux
    port map (
            O => \N__37583\,
            I => \N__37577\
        );

    \I__7947\ : InMux
    port map (
            O => \N__37580\,
            I => \N__37574\
        );

    \I__7946\ : LocalMux
    port map (
            O => \N__37577\,
            I => \N__37569\
        );

    \I__7945\ : LocalMux
    port map (
            O => \N__37574\,
            I => \N__37569\
        );

    \I__7944\ : Odrv4
    port map (
            O => \N__37569\,
            I => n6152
        );

    \I__7943\ : CascadeMux
    port map (
            O => \N__37566\,
            I => \n8_adj_751_cascade_\
        );

    \I__7942\ : CascadeMux
    port map (
            O => \N__37563\,
            I => \n7294_cascade_\
        );

    \I__7941\ : IoInMux
    port map (
            O => \N__37560\,
            I => \N__37557\
        );

    \I__7940\ : LocalMux
    port map (
            O => \N__37557\,
            I => \N__37554\
        );

    \I__7939\ : IoSpan4Mux
    port map (
            O => \N__37554\,
            I => \N__37551\
        );

    \I__7938\ : Span4Mux_s0_h
    port map (
            O => \N__37551\,
            I => \N__37548\
        );

    \I__7937\ : Sp12to4
    port map (
            O => \N__37548\,
            I => \N__37545\
        );

    \I__7936\ : Span12Mux_s11_h
    port map (
            O => \N__37545\,
            I => \N__37541\
        );

    \I__7935\ : InMux
    port map (
            O => \N__37544\,
            I => \N__37537\
        );

    \I__7934\ : Span12Mux_v
    port map (
            O => \N__37541\,
            I => \N__37534\
        );

    \I__7933\ : InMux
    port map (
            O => \N__37540\,
            I => \N__37531\
        );

    \I__7932\ : LocalMux
    port map (
            O => \N__37537\,
            I => \N__37528\
        );

    \I__7931\ : Odrv12
    port map (
            O => \N__37534\,
            I => pin_out_11
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__37531\,
            I => pin_out_11
        );

    \I__7929\ : Odrv4
    port map (
            O => \N__37528\,
            I => pin_out_11
        );

    \I__7928\ : CascadeMux
    port map (
            O => \N__37521\,
            I => \N__37518\
        );

    \I__7927\ : InMux
    port map (
            O => \N__37518\,
            I => \N__37514\
        );

    \I__7926\ : InMux
    port map (
            O => \N__37517\,
            I => \N__37511\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__37514\,
            I => \N__37508\
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__37511\,
            I => \N__37505\
        );

    \I__7923\ : Span4Mux_h
    port map (
            O => \N__37508\,
            I => \N__37502\
        );

    \I__7922\ : Span4Mux_h
    port map (
            O => \N__37505\,
            I => \N__37499\
        );

    \I__7921\ : Odrv4
    port map (
            O => \N__37502\,
            I => n6154
        );

    \I__7920\ : Odrv4
    port map (
            O => \N__37499\,
            I => n6154
        );

    \I__7919\ : InMux
    port map (
            O => \N__37494\,
            I => \N__37490\
        );

    \I__7918\ : InMux
    port map (
            O => \N__37493\,
            I => \N__37487\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__37490\,
            I => \N__37482\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__37487\,
            I => \N__37482\
        );

    \I__7915\ : Span4Mux_v
    port map (
            O => \N__37482\,
            I => \N__37477\
        );

    \I__7914\ : InMux
    port map (
            O => \N__37481\,
            I => \N__37474\
        );

    \I__7913\ : InMux
    port map (
            O => \N__37480\,
            I => \N__37471\
        );

    \I__7912\ : Odrv4
    port map (
            O => \N__37477\,
            I => n8_adj_744
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__37474\,
            I => n8_adj_744
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__37471\,
            I => n8_adj_744
        );

    \I__7909\ : CascadeMux
    port map (
            O => \N__37464\,
            I => \n13048_cascade_\
        );

    \I__7908\ : InMux
    port map (
            O => \N__37461\,
            I => \N__37458\
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__37458\,
            I => \N__37455\
        );

    \I__7906\ : Odrv4
    port map (
            O => \N__37455\,
            I => n13264
        );

    \I__7905\ : InMux
    port map (
            O => \N__37452\,
            I => \N__37449\
        );

    \I__7904\ : LocalMux
    port map (
            O => \N__37449\,
            I => n12091
        );

    \I__7903\ : CascadeMux
    port map (
            O => \N__37446\,
            I => \n24_adj_720_cascade_\
        );

    \I__7902\ : InMux
    port map (
            O => \N__37443\,
            I => \N__37440\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__37440\,
            I => \N__37437\
        );

    \I__7900\ : Odrv4
    port map (
            O => \N__37437\,
            I => n11898
        );

    \I__7899\ : InMux
    port map (
            O => \N__37434\,
            I => \N__37431\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__37431\,
            I => \N__37427\
        );

    \I__7897\ : CascadeMux
    port map (
            O => \N__37430\,
            I => \N__37424\
        );

    \I__7896\ : Span4Mux_v
    port map (
            O => \N__37427\,
            I => \N__37420\
        );

    \I__7895\ : InMux
    port map (
            O => \N__37424\,
            I => \N__37417\
        );

    \I__7894\ : InMux
    port map (
            O => \N__37423\,
            I => \N__37413\
        );

    \I__7893\ : IoSpan4Mux
    port map (
            O => \N__37420\,
            I => \N__37408\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__37417\,
            I => \N__37408\
        );

    \I__7891\ : InMux
    port map (
            O => \N__37416\,
            I => \N__37405\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__37413\,
            I => \N__37402\
        );

    \I__7889\ : Span4Mux_s2_h
    port map (
            O => \N__37408\,
            I => \N__37399\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__37405\,
            I => \N__37396\
        );

    \I__7887\ : Span4Mux_v
    port map (
            O => \N__37402\,
            I => \N__37390\
        );

    \I__7886\ : Span4Mux_v
    port map (
            O => \N__37399\,
            I => \N__37390\
        );

    \I__7885\ : Span4Mux_v
    port map (
            O => \N__37396\,
            I => \N__37387\
        );

    \I__7884\ : InMux
    port map (
            O => \N__37395\,
            I => \N__37384\
        );

    \I__7883\ : Span4Mux_h
    port map (
            O => \N__37390\,
            I => \N__37381\
        );

    \I__7882\ : Span4Mux_h
    port map (
            O => \N__37387\,
            I => \N__37378\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__37384\,
            I => neopxl_color_7
        );

    \I__7880\ : Odrv4
    port map (
            O => \N__37381\,
            I => neopxl_color_7
        );

    \I__7879\ : Odrv4
    port map (
            O => \N__37378\,
            I => neopxl_color_7
        );

    \I__7878\ : SRMux
    port map (
            O => \N__37371\,
            I => \N__37368\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__37368\,
            I => \N__37365\
        );

    \I__7876\ : Span4Mux_v
    port map (
            O => \N__37365\,
            I => \N__37362\
        );

    \I__7875\ : Span4Mux_h
    port map (
            O => \N__37362\,
            I => \N__37359\
        );

    \I__7874\ : Odrv4
    port map (
            O => \N__37359\,
            I => n22_adj_724
        );

    \I__7873\ : InMux
    port map (
            O => \N__37356\,
            I => \N__37353\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__37353\,
            I => n17_adj_765
        );

    \I__7871\ : CascadeMux
    port map (
            O => \N__37350\,
            I => \n16_adj_764_cascade_\
        );

    \I__7870\ : InMux
    port map (
            O => \N__37347\,
            I => \N__37344\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__37344\,
            I => \N__37341\
        );

    \I__7868\ : Odrv12
    port map (
            O => \N__37341\,
            I => n10978
        );

    \I__7867\ : CEMux
    port map (
            O => \N__37338\,
            I => \N__37335\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__37335\,
            I => \N__37332\
        );

    \I__7865\ : Odrv4
    port map (
            O => \N__37332\,
            I => n36
        );

    \I__7864\ : InMux
    port map (
            O => \N__37329\,
            I => \N__37325\
        );

    \I__7863\ : InMux
    port map (
            O => \N__37328\,
            I => \N__37322\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__37325\,
            I => \N__37317\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__37322\,
            I => \N__37317\
        );

    \I__7860\ : Span4Mux_h
    port map (
            O => \N__37317\,
            I => \N__37313\
        );

    \I__7859\ : InMux
    port map (
            O => \N__37316\,
            I => \N__37310\
        );

    \I__7858\ : Odrv4
    port map (
            O => \N__37313\,
            I => \nx.n2095\
        );

    \I__7857\ : LocalMux
    port map (
            O => \N__37310\,
            I => \nx.n2095\
        );

    \I__7856\ : InMux
    port map (
            O => \N__37305\,
            I => \nx.n10687\
        );

    \I__7855\ : InMux
    port map (
            O => \N__37302\,
            I => \N__37298\
        );

    \I__7854\ : InMux
    port map (
            O => \N__37301\,
            I => \N__37295\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__37298\,
            I => \N__37289\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__37295\,
            I => \N__37289\
        );

    \I__7851\ : InMux
    port map (
            O => \N__37294\,
            I => \N__37286\
        );

    \I__7850\ : Odrv4
    port map (
            O => \N__37289\,
            I => \nx.n2094\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__37286\,
            I => \nx.n2094\
        );

    \I__7848\ : InMux
    port map (
            O => \N__37281\,
            I => \bfn_11_25_0_\
        );

    \I__7847\ : InMux
    port map (
            O => \N__37278\,
            I => \N__37274\
        );

    \I__7846\ : InMux
    port map (
            O => \N__37277\,
            I => \N__37271\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__37274\,
            I => \N__37265\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__37271\,
            I => \N__37265\
        );

    \I__7843\ : InMux
    port map (
            O => \N__37270\,
            I => \N__37262\
        );

    \I__7842\ : Odrv4
    port map (
            O => \N__37265\,
            I => \nx.n2093\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__37262\,
            I => \nx.n2093\
        );

    \I__7840\ : CascadeMux
    port map (
            O => \N__37257\,
            I => \N__37239\
        );

    \I__7839\ : CascadeMux
    port map (
            O => \N__37256\,
            I => \N__37236\
        );

    \I__7838\ : CascadeMux
    port map (
            O => \N__37255\,
            I => \N__37233\
        );

    \I__7837\ : CascadeMux
    port map (
            O => \N__37254\,
            I => \N__37230\
        );

    \I__7836\ : CascadeMux
    port map (
            O => \N__37253\,
            I => \N__37227\
        );

    \I__7835\ : CascadeMux
    port map (
            O => \N__37252\,
            I => \N__37224\
        );

    \I__7834\ : CascadeMux
    port map (
            O => \N__37251\,
            I => \N__37221\
        );

    \I__7833\ : CascadeMux
    port map (
            O => \N__37250\,
            I => \N__37218\
        );

    \I__7832\ : CascadeMux
    port map (
            O => \N__37249\,
            I => \N__37215\
        );

    \I__7831\ : CascadeMux
    port map (
            O => \N__37248\,
            I => \N__37212\
        );

    \I__7830\ : CascadeMux
    port map (
            O => \N__37247\,
            I => \N__37209\
        );

    \I__7829\ : CascadeMux
    port map (
            O => \N__37246\,
            I => \N__37206\
        );

    \I__7828\ : CascadeMux
    port map (
            O => \N__37245\,
            I => \N__37203\
        );

    \I__7827\ : CascadeMux
    port map (
            O => \N__37244\,
            I => \N__37200\
        );

    \I__7826\ : CascadeMux
    port map (
            O => \N__37243\,
            I => \N__37197\
        );

    \I__7825\ : CascadeMux
    port map (
            O => \N__37242\,
            I => \N__37194\
        );

    \I__7824\ : InMux
    port map (
            O => \N__37239\,
            I => \N__37190\
        );

    \I__7823\ : InMux
    port map (
            O => \N__37236\,
            I => \N__37187\
        );

    \I__7822\ : InMux
    port map (
            O => \N__37233\,
            I => \N__37178\
        );

    \I__7821\ : InMux
    port map (
            O => \N__37230\,
            I => \N__37178\
        );

    \I__7820\ : InMux
    port map (
            O => \N__37227\,
            I => \N__37178\
        );

    \I__7819\ : InMux
    port map (
            O => \N__37224\,
            I => \N__37178\
        );

    \I__7818\ : InMux
    port map (
            O => \N__37221\,
            I => \N__37169\
        );

    \I__7817\ : InMux
    port map (
            O => \N__37218\,
            I => \N__37169\
        );

    \I__7816\ : InMux
    port map (
            O => \N__37215\,
            I => \N__37169\
        );

    \I__7815\ : InMux
    port map (
            O => \N__37212\,
            I => \N__37169\
        );

    \I__7814\ : InMux
    port map (
            O => \N__37209\,
            I => \N__37162\
        );

    \I__7813\ : InMux
    port map (
            O => \N__37206\,
            I => \N__37162\
        );

    \I__7812\ : InMux
    port map (
            O => \N__37203\,
            I => \N__37162\
        );

    \I__7811\ : InMux
    port map (
            O => \N__37200\,
            I => \N__37155\
        );

    \I__7810\ : InMux
    port map (
            O => \N__37197\,
            I => \N__37155\
        );

    \I__7809\ : InMux
    port map (
            O => \N__37194\,
            I => \N__37155\
        );

    \I__7808\ : InMux
    port map (
            O => \N__37193\,
            I => \N__37152\
        );

    \I__7807\ : LocalMux
    port map (
            O => \N__37190\,
            I => \nx.n2126\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__37187\,
            I => \nx.n2126\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__37178\,
            I => \nx.n2126\
        );

    \I__7804\ : LocalMux
    port map (
            O => \N__37169\,
            I => \nx.n2126\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__37162\,
            I => \nx.n2126\
        );

    \I__7802\ : LocalMux
    port map (
            O => \N__37155\,
            I => \nx.n2126\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__37152\,
            I => \nx.n2126\
        );

    \I__7800\ : InMux
    port map (
            O => \N__37137\,
            I => \nx.n10689\
        );

    \I__7799\ : CascadeMux
    port map (
            O => \N__37134\,
            I => \N__37131\
        );

    \I__7798\ : InMux
    port map (
            O => \N__37131\,
            I => \N__37128\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__37128\,
            I => n12171
        );

    \I__7796\ : InMux
    port map (
            O => \N__37125\,
            I => \N__37122\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__37122\,
            I => n6_adj_761
        );

    \I__7794\ : CascadeMux
    port map (
            O => \N__37119\,
            I => \n15_cascade_\
        );

    \I__7793\ : InMux
    port map (
            O => \N__37116\,
            I => \N__37113\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__37113\,
            I => n14
        );

    \I__7791\ : InMux
    port map (
            O => \N__37110\,
            I => \N__37106\
        );

    \I__7790\ : InMux
    port map (
            O => \N__37109\,
            I => \N__37103\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__37106\,
            I => \N__37098\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__37103\,
            I => \N__37098\
        );

    \I__7787\ : Span4Mux_h
    port map (
            O => \N__37098\,
            I => \N__37094\
        );

    \I__7786\ : InMux
    port map (
            O => \N__37097\,
            I => \N__37091\
        );

    \I__7785\ : Odrv4
    port map (
            O => \N__37094\,
            I => \nx.n2103\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__37091\,
            I => \nx.n2103\
        );

    \I__7783\ : InMux
    port map (
            O => \N__37086\,
            I => \nx.n10679\
        );

    \I__7782\ : InMux
    port map (
            O => \N__37083\,
            I => \N__37078\
        );

    \I__7781\ : InMux
    port map (
            O => \N__37082\,
            I => \N__37075\
        );

    \I__7780\ : InMux
    port map (
            O => \N__37081\,
            I => \N__37072\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__37078\,
            I => \nx.n2102\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__37075\,
            I => \nx.n2102\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__37072\,
            I => \nx.n2102\
        );

    \I__7776\ : InMux
    port map (
            O => \N__37065\,
            I => \bfn_11_24_0_\
        );

    \I__7775\ : InMux
    port map (
            O => \N__37062\,
            I => \N__37057\
        );

    \I__7774\ : InMux
    port map (
            O => \N__37061\,
            I => \N__37054\
        );

    \I__7773\ : InMux
    port map (
            O => \N__37060\,
            I => \N__37051\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__37057\,
            I => \nx.n2101\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__37054\,
            I => \nx.n2101\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__37051\,
            I => \nx.n2101\
        );

    \I__7769\ : InMux
    port map (
            O => \N__37044\,
            I => \nx.n10681\
        );

    \I__7768\ : InMux
    port map (
            O => \N__37041\,
            I => \N__37037\
        );

    \I__7767\ : InMux
    port map (
            O => \N__37040\,
            I => \N__37034\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__37037\,
            I => \N__37031\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__37034\,
            I => \N__37028\
        );

    \I__7764\ : Span4Mux_v
    port map (
            O => \N__37031\,
            I => \N__37022\
        );

    \I__7763\ : Span4Mux_v
    port map (
            O => \N__37028\,
            I => \N__37022\
        );

    \I__7762\ : InMux
    port map (
            O => \N__37027\,
            I => \N__37019\
        );

    \I__7761\ : Odrv4
    port map (
            O => \N__37022\,
            I => \nx.n2100\
        );

    \I__7760\ : LocalMux
    port map (
            O => \N__37019\,
            I => \nx.n2100\
        );

    \I__7759\ : InMux
    port map (
            O => \N__37014\,
            I => \nx.n10682\
        );

    \I__7758\ : InMux
    port map (
            O => \N__37011\,
            I => \N__37007\
        );

    \I__7757\ : InMux
    port map (
            O => \N__37010\,
            I => \N__37004\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__37007\,
            I => \N__36999\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__37004\,
            I => \N__36999\
        );

    \I__7754\ : Span4Mux_h
    port map (
            O => \N__36999\,
            I => \N__36996\
        );

    \I__7753\ : Odrv4
    port map (
            O => \N__36996\,
            I => \nx.n2099\
        );

    \I__7752\ : InMux
    port map (
            O => \N__36993\,
            I => \nx.n10683\
        );

    \I__7751\ : InMux
    port map (
            O => \N__36990\,
            I => \N__36986\
        );

    \I__7750\ : InMux
    port map (
            O => \N__36989\,
            I => \N__36983\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__36986\,
            I => \N__36980\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__36983\,
            I => \N__36977\
        );

    \I__7747\ : Span4Mux_v
    port map (
            O => \N__36980\,
            I => \N__36971\
        );

    \I__7746\ : Span4Mux_v
    port map (
            O => \N__36977\,
            I => \N__36971\
        );

    \I__7745\ : InMux
    port map (
            O => \N__36976\,
            I => \N__36968\
        );

    \I__7744\ : Odrv4
    port map (
            O => \N__36971\,
            I => \nx.n2098\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__36968\,
            I => \nx.n2098\
        );

    \I__7742\ : InMux
    port map (
            O => \N__36963\,
            I => \nx.n10684\
        );

    \I__7741\ : InMux
    port map (
            O => \N__36960\,
            I => \N__36957\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__36957\,
            I => \N__36953\
        );

    \I__7739\ : InMux
    port map (
            O => \N__36956\,
            I => \N__36950\
        );

    \I__7738\ : Odrv4
    port map (
            O => \N__36953\,
            I => \nx.n2097\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__36950\,
            I => \nx.n2097\
        );

    \I__7736\ : InMux
    port map (
            O => \N__36945\,
            I => \nx.n10685\
        );

    \I__7735\ : InMux
    port map (
            O => \N__36942\,
            I => \N__36937\
        );

    \I__7734\ : InMux
    port map (
            O => \N__36941\,
            I => \N__36934\
        );

    \I__7733\ : InMux
    port map (
            O => \N__36940\,
            I => \N__36931\
        );

    \I__7732\ : LocalMux
    port map (
            O => \N__36937\,
            I => \nx.n2096\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__36934\,
            I => \nx.n2096\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__36931\,
            I => \nx.n2096\
        );

    \I__7729\ : InMux
    port map (
            O => \N__36924\,
            I => \nx.n10686\
        );

    \I__7728\ : CascadeMux
    port map (
            O => \N__36921\,
            I => \nx.n2293_cascade_\
        );

    \I__7727\ : InMux
    port map (
            O => \N__36918\,
            I => \N__36914\
        );

    \I__7726\ : InMux
    port map (
            O => \N__36917\,
            I => \N__36911\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__36914\,
            I => \N__36905\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__36911\,
            I => \N__36905\
        );

    \I__7723\ : InMux
    port map (
            O => \N__36910\,
            I => \N__36902\
        );

    \I__7722\ : Span4Mux_v
    port map (
            O => \N__36905\,
            I => \N__36896\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__36902\,
            I => \N__36896\
        );

    \I__7720\ : InMux
    port map (
            O => \N__36901\,
            I => \N__36892\
        );

    \I__7719\ : Span4Mux_h
    port map (
            O => \N__36896\,
            I => \N__36889\
        );

    \I__7718\ : InMux
    port map (
            O => \N__36895\,
            I => \N__36886\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__36892\,
            I => \N__36881\
        );

    \I__7716\ : Span4Mux_v
    port map (
            O => \N__36889\,
            I => \N__36881\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__36886\,
            I => \nx.bit_ctr_14\
        );

    \I__7714\ : Odrv4
    port map (
            O => \N__36881\,
            I => \nx.bit_ctr_14\
        );

    \I__7713\ : InMux
    port map (
            O => \N__36876\,
            I => \bfn_11_23_0_\
        );

    \I__7712\ : CascadeMux
    port map (
            O => \N__36873\,
            I => \N__36870\
        );

    \I__7711\ : InMux
    port map (
            O => \N__36870\,
            I => \N__36865\
        );

    \I__7710\ : InMux
    port map (
            O => \N__36869\,
            I => \N__36862\
        );

    \I__7709\ : InMux
    port map (
            O => \N__36868\,
            I => \N__36859\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__36865\,
            I => \N__36856\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__36862\,
            I => \nx.n2109\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__36859\,
            I => \nx.n2109\
        );

    \I__7705\ : Odrv4
    port map (
            O => \N__36856\,
            I => \nx.n2109\
        );

    \I__7704\ : CascadeMux
    port map (
            O => \N__36849\,
            I => \N__36845\
        );

    \I__7703\ : CascadeMux
    port map (
            O => \N__36848\,
            I => \N__36842\
        );

    \I__7702\ : InMux
    port map (
            O => \N__36845\,
            I => \N__36839\
        );

    \I__7701\ : InMux
    port map (
            O => \N__36842\,
            I => \N__36836\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__36839\,
            I => \nx.n13436\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__36836\,
            I => \nx.n13436\
        );

    \I__7698\ : InMux
    port map (
            O => \N__36831\,
            I => \nx.n10673\
        );

    \I__7697\ : InMux
    port map (
            O => \N__36828\,
            I => \N__36823\
        );

    \I__7696\ : InMux
    port map (
            O => \N__36827\,
            I => \N__36820\
        );

    \I__7695\ : InMux
    port map (
            O => \N__36826\,
            I => \N__36817\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__36823\,
            I => \nx.n2108\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__36820\,
            I => \nx.n2108\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__36817\,
            I => \nx.n2108\
        );

    \I__7691\ : InMux
    port map (
            O => \N__36810\,
            I => \nx.n10674\
        );

    \I__7690\ : InMux
    port map (
            O => \N__36807\,
            I => \N__36803\
        );

    \I__7689\ : InMux
    port map (
            O => \N__36806\,
            I => \N__36800\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__36803\,
            I => \nx.n2107\
        );

    \I__7687\ : LocalMux
    port map (
            O => \N__36800\,
            I => \nx.n2107\
        );

    \I__7686\ : InMux
    port map (
            O => \N__36795\,
            I => \nx.n10675\
        );

    \I__7685\ : InMux
    port map (
            O => \N__36792\,
            I => \N__36787\
        );

    \I__7684\ : InMux
    port map (
            O => \N__36791\,
            I => \N__36784\
        );

    \I__7683\ : InMux
    port map (
            O => \N__36790\,
            I => \N__36781\
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__36787\,
            I => \nx.n2106\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__36784\,
            I => \nx.n2106\
        );

    \I__7680\ : LocalMux
    port map (
            O => \N__36781\,
            I => \nx.n2106\
        );

    \I__7679\ : InMux
    port map (
            O => \N__36774\,
            I => \nx.n10676\
        );

    \I__7678\ : InMux
    port map (
            O => \N__36771\,
            I => \N__36767\
        );

    \I__7677\ : InMux
    port map (
            O => \N__36770\,
            I => \N__36764\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__36767\,
            I => \N__36759\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__36764\,
            I => \N__36759\
        );

    \I__7674\ : Span4Mux_h
    port map (
            O => \N__36759\,
            I => \N__36756\
        );

    \I__7673\ : Odrv4
    port map (
            O => \N__36756\,
            I => \nx.n2105\
        );

    \I__7672\ : InMux
    port map (
            O => \N__36753\,
            I => \nx.n10677\
        );

    \I__7671\ : InMux
    port map (
            O => \N__36750\,
            I => \N__36746\
        );

    \I__7670\ : InMux
    port map (
            O => \N__36749\,
            I => \N__36743\
        );

    \I__7669\ : LocalMux
    port map (
            O => \N__36746\,
            I => \N__36738\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__36743\,
            I => \N__36738\
        );

    \I__7667\ : Span4Mux_h
    port map (
            O => \N__36738\,
            I => \N__36734\
        );

    \I__7666\ : InMux
    port map (
            O => \N__36737\,
            I => \N__36731\
        );

    \I__7665\ : Odrv4
    port map (
            O => \N__36734\,
            I => \nx.n2104\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__36731\,
            I => \nx.n2104\
        );

    \I__7663\ : InMux
    port map (
            O => \N__36726\,
            I => \nx.n10678\
        );

    \I__7662\ : CascadeMux
    port map (
            O => \N__36723\,
            I => \nx.n2296_cascade_\
        );

    \I__7661\ : CascadeMux
    port map (
            O => \N__36720\,
            I => \nx.n2395_cascade_\
        );

    \I__7660\ : CascadeMux
    port map (
            O => \N__36717\,
            I => \nx.n2494_cascade_\
        );

    \I__7659\ : InMux
    port map (
            O => \N__36714\,
            I => \N__36709\
        );

    \I__7658\ : InMux
    port map (
            O => \N__36713\,
            I => \N__36706\
        );

    \I__7657\ : InMux
    port map (
            O => \N__36712\,
            I => \N__36703\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__36709\,
            I => \N__36700\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__36706\,
            I => \N__36697\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__36703\,
            I => \nx.n2593\
        );

    \I__7653\ : Odrv4
    port map (
            O => \N__36700\,
            I => \nx.n2593\
        );

    \I__7652\ : Odrv4
    port map (
            O => \N__36697\,
            I => \nx.n2593\
        );

    \I__7651\ : CascadeMux
    port map (
            O => \N__36690\,
            I => \nx.n2504_cascade_\
        );

    \I__7650\ : InMux
    port map (
            O => \N__36687\,
            I => \N__36683\
        );

    \I__7649\ : CascadeMux
    port map (
            O => \N__36686\,
            I => \N__36680\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__36683\,
            I => \N__36677\
        );

    \I__7647\ : InMux
    port map (
            O => \N__36680\,
            I => \N__36673\
        );

    \I__7646\ : Span4Mux_h
    port map (
            O => \N__36677\,
            I => \N__36670\
        );

    \I__7645\ : InMux
    port map (
            O => \N__36676\,
            I => \N__36667\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__36673\,
            I => \N__36664\
        );

    \I__7643\ : Odrv4
    port map (
            O => \N__36670\,
            I => \nx.n2603\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__36667\,
            I => \nx.n2603\
        );

    \I__7641\ : Odrv4
    port map (
            O => \N__36664\,
            I => \nx.n2603\
        );

    \I__7640\ : CascadeMux
    port map (
            O => \N__36657\,
            I => \N__36653\
        );

    \I__7639\ : CascadeMux
    port map (
            O => \N__36656\,
            I => \N__36649\
        );

    \I__7638\ : InMux
    port map (
            O => \N__36653\,
            I => \N__36646\
        );

    \I__7637\ : InMux
    port map (
            O => \N__36652\,
            I => \N__36641\
        );

    \I__7636\ : InMux
    port map (
            O => \N__36649\,
            I => \N__36641\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__36646\,
            I => \nx.n2589\
        );

    \I__7634\ : LocalMux
    port map (
            O => \N__36641\,
            I => \nx.n2589\
        );

    \I__7633\ : CascadeMux
    port map (
            O => \N__36636\,
            I => \N__36633\
        );

    \I__7632\ : InMux
    port map (
            O => \N__36633\,
            I => \N__36630\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__36630\,
            I => \N__36626\
        );

    \I__7630\ : InMux
    port map (
            O => \N__36629\,
            I => \N__36622\
        );

    \I__7629\ : Span4Mux_h
    port map (
            O => \N__36626\,
            I => \N__36619\
        );

    \I__7628\ : InMux
    port map (
            O => \N__36625\,
            I => \N__36616\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__36622\,
            I => \nx.n2688\
        );

    \I__7626\ : Odrv4
    port map (
            O => \N__36619\,
            I => \nx.n2688\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__36616\,
            I => \nx.n2688\
        );

    \I__7624\ : CascadeMux
    port map (
            O => \N__36609\,
            I => \N__36606\
        );

    \I__7623\ : InMux
    port map (
            O => \N__36606\,
            I => \N__36602\
        );

    \I__7622\ : CascadeMux
    port map (
            O => \N__36605\,
            I => \N__36597\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__36602\,
            I => \N__36587\
        );

    \I__7620\ : InMux
    port map (
            O => \N__36601\,
            I => \N__36583\
        );

    \I__7619\ : InMux
    port map (
            O => \N__36600\,
            I => \N__36576\
        );

    \I__7618\ : InMux
    port map (
            O => \N__36597\,
            I => \N__36576\
        );

    \I__7617\ : InMux
    port map (
            O => \N__36596\,
            I => \N__36576\
        );

    \I__7616\ : InMux
    port map (
            O => \N__36595\,
            I => \N__36570\
        );

    \I__7615\ : InMux
    port map (
            O => \N__36594\,
            I => \N__36570\
        );

    \I__7614\ : CascadeMux
    port map (
            O => \N__36593\,
            I => \N__36566\
        );

    \I__7613\ : CascadeMux
    port map (
            O => \N__36592\,
            I => \N__36561\
        );

    \I__7612\ : CascadeMux
    port map (
            O => \N__36591\,
            I => \N__36557\
        );

    \I__7611\ : CascadeMux
    port map (
            O => \N__36590\,
            I => \N__36551\
        );

    \I__7610\ : Span4Mux_v
    port map (
            O => \N__36587\,
            I => \N__36545\
        );

    \I__7609\ : InMux
    port map (
            O => \N__36586\,
            I => \N__36542\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__36583\,
            I => \N__36537\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__36576\,
            I => \N__36537\
        );

    \I__7606\ : InMux
    port map (
            O => \N__36575\,
            I => \N__36534\
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__36570\,
            I => \N__36531\
        );

    \I__7604\ : InMux
    port map (
            O => \N__36569\,
            I => \N__36528\
        );

    \I__7603\ : InMux
    port map (
            O => \N__36566\,
            I => \N__36523\
        );

    \I__7602\ : InMux
    port map (
            O => \N__36565\,
            I => \N__36523\
        );

    \I__7601\ : InMux
    port map (
            O => \N__36564\,
            I => \N__36508\
        );

    \I__7600\ : InMux
    port map (
            O => \N__36561\,
            I => \N__36508\
        );

    \I__7599\ : InMux
    port map (
            O => \N__36560\,
            I => \N__36508\
        );

    \I__7598\ : InMux
    port map (
            O => \N__36557\,
            I => \N__36508\
        );

    \I__7597\ : InMux
    port map (
            O => \N__36556\,
            I => \N__36508\
        );

    \I__7596\ : InMux
    port map (
            O => \N__36555\,
            I => \N__36508\
        );

    \I__7595\ : InMux
    port map (
            O => \N__36554\,
            I => \N__36508\
        );

    \I__7594\ : InMux
    port map (
            O => \N__36551\,
            I => \N__36499\
        );

    \I__7593\ : InMux
    port map (
            O => \N__36550\,
            I => \N__36499\
        );

    \I__7592\ : InMux
    port map (
            O => \N__36549\,
            I => \N__36499\
        );

    \I__7591\ : InMux
    port map (
            O => \N__36548\,
            I => \N__36499\
        );

    \I__7590\ : Sp12to4
    port map (
            O => \N__36545\,
            I => \N__36494\
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__36542\,
            I => \N__36494\
        );

    \I__7588\ : Odrv4
    port map (
            O => \N__36537\,
            I => \nx.n2720\
        );

    \I__7587\ : LocalMux
    port map (
            O => \N__36534\,
            I => \nx.n2720\
        );

    \I__7586\ : Odrv12
    port map (
            O => \N__36531\,
            I => \nx.n2720\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__36528\,
            I => \nx.n2720\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__36523\,
            I => \nx.n2720\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__36508\,
            I => \nx.n2720\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__36499\,
            I => \nx.n2720\
        );

    \I__7581\ : Odrv12
    port map (
            O => \N__36494\,
            I => \nx.n2720\
        );

    \I__7580\ : InMux
    port map (
            O => \N__36477\,
            I => \N__36474\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__36474\,
            I => \N__36471\
        );

    \I__7578\ : Span4Mux_h
    port map (
            O => \N__36471\,
            I => \N__36468\
        );

    \I__7577\ : Odrv4
    port map (
            O => \N__36468\,
            I => \nx.n2755\
        );

    \I__7576\ : CascadeMux
    port map (
            O => \N__36465\,
            I => \N__36462\
        );

    \I__7575\ : InMux
    port map (
            O => \N__36462\,
            I => \N__36459\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__36459\,
            I => \N__36454\
        );

    \I__7573\ : InMux
    port map (
            O => \N__36458\,
            I => \N__36449\
        );

    \I__7572\ : InMux
    port map (
            O => \N__36457\,
            I => \N__36449\
        );

    \I__7571\ : Span4Mux_h
    port map (
            O => \N__36454\,
            I => \N__36444\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__36449\,
            I => \N__36444\
        );

    \I__7569\ : Span4Mux_h
    port map (
            O => \N__36444\,
            I => \N__36441\
        );

    \I__7568\ : Odrv4
    port map (
            O => \N__36441\,
            I => \nx.n2787\
        );

    \I__7567\ : CascadeMux
    port map (
            O => \N__36438\,
            I => \N__36435\
        );

    \I__7566\ : InMux
    port map (
            O => \N__36435\,
            I => \N__36431\
        );

    \I__7565\ : CascadeMux
    port map (
            O => \N__36434\,
            I => \N__36428\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__36431\,
            I => \N__36424\
        );

    \I__7563\ : InMux
    port map (
            O => \N__36428\,
            I => \N__36421\
        );

    \I__7562\ : InMux
    port map (
            O => \N__36427\,
            I => \N__36418\
        );

    \I__7561\ : Odrv12
    port map (
            O => \N__36424\,
            I => \nx.n2590\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__36421\,
            I => \nx.n2590\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__36418\,
            I => \nx.n2590\
        );

    \I__7558\ : InMux
    port map (
            O => \N__36411\,
            I => \N__36407\
        );

    \I__7557\ : CascadeMux
    port map (
            O => \N__36410\,
            I => \N__36404\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__36407\,
            I => \N__36400\
        );

    \I__7555\ : InMux
    port map (
            O => \N__36404\,
            I => \N__36397\
        );

    \I__7554\ : InMux
    port map (
            O => \N__36403\,
            I => \N__36394\
        );

    \I__7553\ : Odrv4
    port map (
            O => \N__36400\,
            I => \nx.n2591\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__36397\,
            I => \nx.n2591\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__36394\,
            I => \nx.n2591\
        );

    \I__7550\ : InMux
    port map (
            O => \N__36387\,
            I => \N__36383\
        );

    \I__7549\ : CascadeMux
    port map (
            O => \N__36386\,
            I => \N__36380\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__36383\,
            I => \N__36377\
        );

    \I__7547\ : InMux
    port map (
            O => \N__36380\,
            I => \N__36374\
        );

    \I__7546\ : Odrv4
    port map (
            O => \N__36377\,
            I => \nx.n2596\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__36374\,
            I => \nx.n2596\
        );

    \I__7544\ : InMux
    port map (
            O => \N__36369\,
            I => \N__36366\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__36366\,
            I => \N__36362\
        );

    \I__7542\ : CascadeMux
    port map (
            O => \N__36365\,
            I => \N__36358\
        );

    \I__7541\ : Span4Mux_h
    port map (
            O => \N__36362\,
            I => \N__36355\
        );

    \I__7540\ : InMux
    port map (
            O => \N__36361\,
            I => \N__36352\
        );

    \I__7539\ : InMux
    port map (
            O => \N__36358\,
            I => \N__36349\
        );

    \I__7538\ : Odrv4
    port map (
            O => \N__36355\,
            I => \nx.n2599\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__36352\,
            I => \nx.n2599\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__36349\,
            I => \nx.n2599\
        );

    \I__7535\ : CascadeMux
    port map (
            O => \N__36342\,
            I => \nx.n2596_cascade_\
        );

    \I__7534\ : InMux
    port map (
            O => \N__36339\,
            I => \N__36336\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__36336\,
            I => \N__36332\
        );

    \I__7532\ : CascadeMux
    port map (
            O => \N__36335\,
            I => \N__36328\
        );

    \I__7531\ : Span4Mux_h
    port map (
            O => \N__36332\,
            I => \N__36325\
        );

    \I__7530\ : InMux
    port map (
            O => \N__36331\,
            I => \N__36322\
        );

    \I__7529\ : InMux
    port map (
            O => \N__36328\,
            I => \N__36319\
        );

    \I__7528\ : Odrv4
    port map (
            O => \N__36325\,
            I => \nx.n2604\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__36322\,
            I => \nx.n2604\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__36319\,
            I => \nx.n2604\
        );

    \I__7525\ : InMux
    port map (
            O => \N__36312\,
            I => \N__36309\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__36309\,
            I => \nx.n37\
        );

    \I__7523\ : InMux
    port map (
            O => \N__36306\,
            I => \N__36303\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__36303\,
            I => \N__36298\
        );

    \I__7521\ : CascadeMux
    port map (
            O => \N__36302\,
            I => \N__36295\
        );

    \I__7520\ : CascadeMux
    port map (
            O => \N__36301\,
            I => \N__36292\
        );

    \I__7519\ : Span4Mux_v
    port map (
            O => \N__36298\,
            I => \N__36289\
        );

    \I__7518\ : InMux
    port map (
            O => \N__36295\,
            I => \N__36286\
        );

    \I__7517\ : InMux
    port map (
            O => \N__36292\,
            I => \N__36283\
        );

    \I__7516\ : Odrv4
    port map (
            O => \N__36289\,
            I => \nx.n2598\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__36286\,
            I => \nx.n2598\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__36283\,
            I => \nx.n2598\
        );

    \I__7513\ : InMux
    port map (
            O => \N__36276\,
            I => \N__36273\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__36273\,
            I => \nx.n38\
        );

    \I__7511\ : CascadeMux
    port map (
            O => \N__36270\,
            I => \N__36267\
        );

    \I__7510\ : InMux
    port map (
            O => \N__36267\,
            I => \N__36264\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__36264\,
            I => \N__36260\
        );

    \I__7508\ : CascadeMux
    port map (
            O => \N__36263\,
            I => \N__36256\
        );

    \I__7507\ : Span4Mux_h
    port map (
            O => \N__36260\,
            I => \N__36253\
        );

    \I__7506\ : InMux
    port map (
            O => \N__36259\,
            I => \N__36250\
        );

    \I__7505\ : InMux
    port map (
            O => \N__36256\,
            I => \N__36247\
        );

    \I__7504\ : Odrv4
    port map (
            O => \N__36253\,
            I => \nx.n2602\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__36250\,
            I => \nx.n2602\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__36247\,
            I => \nx.n2602\
        );

    \I__7501\ : CascadeMux
    port map (
            O => \N__36240\,
            I => \N__36237\
        );

    \I__7500\ : InMux
    port map (
            O => \N__36237\,
            I => \N__36233\
        );

    \I__7499\ : InMux
    port map (
            O => \N__36236\,
            I => \N__36230\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__36233\,
            I => \N__36227\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__36230\,
            I => \nx.n2606\
        );

    \I__7496\ : Odrv4
    port map (
            O => \N__36227\,
            I => \nx.n2606\
        );

    \I__7495\ : InMux
    port map (
            O => \N__36222\,
            I => \N__36219\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__36219\,
            I => \N__36216\
        );

    \I__7493\ : Odrv4
    port map (
            O => \N__36216\,
            I => \nx.n2673\
        );

    \I__7492\ : CascadeMux
    port map (
            O => \N__36213\,
            I => \nx.n2606_cascade_\
        );

    \I__7491\ : CascadeMux
    port map (
            O => \N__36210\,
            I => \N__36203\
        );

    \I__7490\ : CascadeMux
    port map (
            O => \N__36209\,
            I => \N__36200\
        );

    \I__7489\ : InMux
    port map (
            O => \N__36208\,
            I => \N__36188\
        );

    \I__7488\ : InMux
    port map (
            O => \N__36207\,
            I => \N__36185\
        );

    \I__7487\ : InMux
    port map (
            O => \N__36206\,
            I => \N__36176\
        );

    \I__7486\ : InMux
    port map (
            O => \N__36203\,
            I => \N__36176\
        );

    \I__7485\ : InMux
    port map (
            O => \N__36200\,
            I => \N__36176\
        );

    \I__7484\ : InMux
    port map (
            O => \N__36199\,
            I => \N__36176\
        );

    \I__7483\ : CascadeMux
    port map (
            O => \N__36198\,
            I => \N__36173\
        );

    \I__7482\ : CascadeMux
    port map (
            O => \N__36197\,
            I => \N__36167\
        );

    \I__7481\ : CascadeMux
    port map (
            O => \N__36196\,
            I => \N__36163\
        );

    \I__7480\ : CascadeMux
    port map (
            O => \N__36195\,
            I => \N__36160\
        );

    \I__7479\ : CascadeMux
    port map (
            O => \N__36194\,
            I => \N__36155\
        );

    \I__7478\ : CascadeMux
    port map (
            O => \N__36193\,
            I => \N__36152\
        );

    \I__7477\ : CascadeMux
    port map (
            O => \N__36192\,
            I => \N__36148\
        );

    \I__7476\ : CascadeMux
    port map (
            O => \N__36191\,
            I => \N__36145\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__36188\,
            I => \N__36141\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__36185\,
            I => \N__36136\
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__36176\,
            I => \N__36136\
        );

    \I__7472\ : InMux
    port map (
            O => \N__36173\,
            I => \N__36133\
        );

    \I__7471\ : InMux
    port map (
            O => \N__36172\,
            I => \N__36130\
        );

    \I__7470\ : InMux
    port map (
            O => \N__36171\,
            I => \N__36121\
        );

    \I__7469\ : InMux
    port map (
            O => \N__36170\,
            I => \N__36121\
        );

    \I__7468\ : InMux
    port map (
            O => \N__36167\,
            I => \N__36121\
        );

    \I__7467\ : InMux
    port map (
            O => \N__36166\,
            I => \N__36121\
        );

    \I__7466\ : InMux
    port map (
            O => \N__36163\,
            I => \N__36114\
        );

    \I__7465\ : InMux
    port map (
            O => \N__36160\,
            I => \N__36114\
        );

    \I__7464\ : InMux
    port map (
            O => \N__36159\,
            I => \N__36114\
        );

    \I__7463\ : InMux
    port map (
            O => \N__36158\,
            I => \N__36099\
        );

    \I__7462\ : InMux
    port map (
            O => \N__36155\,
            I => \N__36099\
        );

    \I__7461\ : InMux
    port map (
            O => \N__36152\,
            I => \N__36099\
        );

    \I__7460\ : InMux
    port map (
            O => \N__36151\,
            I => \N__36099\
        );

    \I__7459\ : InMux
    port map (
            O => \N__36148\,
            I => \N__36099\
        );

    \I__7458\ : InMux
    port map (
            O => \N__36145\,
            I => \N__36099\
        );

    \I__7457\ : InMux
    port map (
            O => \N__36144\,
            I => \N__36099\
        );

    \I__7456\ : Span4Mux_v
    port map (
            O => \N__36141\,
            I => \N__36094\
        );

    \I__7455\ : Span4Mux_v
    port map (
            O => \N__36136\,
            I => \N__36094\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__36133\,
            I => \nx.n2621\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__36130\,
            I => \nx.n2621\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__36121\,
            I => \nx.n2621\
        );

    \I__7451\ : LocalMux
    port map (
            O => \N__36114\,
            I => \nx.n2621\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__36099\,
            I => \nx.n2621\
        );

    \I__7449\ : Odrv4
    port map (
            O => \N__36094\,
            I => \nx.n2621\
        );

    \I__7448\ : CascadeMux
    port map (
            O => \N__36081\,
            I => \N__36077\
        );

    \I__7447\ : InMux
    port map (
            O => \N__36080\,
            I => \N__36074\
        );

    \I__7446\ : InMux
    port map (
            O => \N__36077\,
            I => \N__36071\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__36074\,
            I => \N__36068\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__36071\,
            I => \N__36065\
        );

    \I__7443\ : Odrv4
    port map (
            O => \N__36068\,
            I => \nx.n2705\
        );

    \I__7442\ : Odrv12
    port map (
            O => \N__36065\,
            I => \nx.n2705\
        );

    \I__7441\ : InMux
    port map (
            O => \N__36060\,
            I => \N__36057\
        );

    \I__7440\ : LocalMux
    port map (
            O => \N__36057\,
            I => \N__36054\
        );

    \I__7439\ : Odrv12
    port map (
            O => \N__36054\,
            I => \nx.n2772\
        );

    \I__7438\ : CascadeMux
    port map (
            O => \N__36051\,
            I => \nx.n2705_cascade_\
        );

    \I__7437\ : CascadeMux
    port map (
            O => \N__36048\,
            I => \N__36044\
        );

    \I__7436\ : CascadeMux
    port map (
            O => \N__36047\,
            I => \N__36040\
        );

    \I__7435\ : InMux
    port map (
            O => \N__36044\,
            I => \N__36037\
        );

    \I__7434\ : InMux
    port map (
            O => \N__36043\,
            I => \N__36034\
        );

    \I__7433\ : InMux
    port map (
            O => \N__36040\,
            I => \N__36031\
        );

    \I__7432\ : LocalMux
    port map (
            O => \N__36037\,
            I => \N__36028\
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__36034\,
            I => \N__36025\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__36031\,
            I => \N__36022\
        );

    \I__7429\ : Span4Mux_v
    port map (
            O => \N__36028\,
            I => \N__36015\
        );

    \I__7428\ : Span4Mux_v
    port map (
            O => \N__36025\,
            I => \N__36015\
        );

    \I__7427\ : Span4Mux_h
    port map (
            O => \N__36022\,
            I => \N__36015\
        );

    \I__7426\ : Span4Mux_h
    port map (
            O => \N__36015\,
            I => \N__36012\
        );

    \I__7425\ : Odrv4
    port map (
            O => \N__36012\,
            I => \nx.n2804\
        );

    \I__7424\ : InMux
    port map (
            O => \N__36009\,
            I => \N__36005\
        );

    \I__7423\ : CascadeMux
    port map (
            O => \N__36008\,
            I => \N__36001\
        );

    \I__7422\ : LocalMux
    port map (
            O => \N__36005\,
            I => \N__35998\
        );

    \I__7421\ : InMux
    port map (
            O => \N__36004\,
            I => \N__35995\
        );

    \I__7420\ : InMux
    port map (
            O => \N__36001\,
            I => \N__35992\
        );

    \I__7419\ : Span4Mux_h
    port map (
            O => \N__35998\,
            I => \N__35989\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__35995\,
            I => \nx.n2594\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__35992\,
            I => \nx.n2594\
        );

    \I__7416\ : Odrv4
    port map (
            O => \N__35989\,
            I => \nx.n2594\
        );

    \I__7415\ : CascadeMux
    port map (
            O => \N__35982\,
            I => \N__35978\
        );

    \I__7414\ : InMux
    port map (
            O => \N__35981\,
            I => \N__35975\
        );

    \I__7413\ : InMux
    port map (
            O => \N__35978\,
            I => \N__35972\
        );

    \I__7412\ : LocalMux
    port map (
            O => \N__35975\,
            I => n6156
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__35972\,
            I => n6156
        );

    \I__7410\ : CascadeMux
    port map (
            O => \N__35967\,
            I => \n7266_cascade_\
        );

    \I__7409\ : IoInMux
    port map (
            O => \N__35964\,
            I => \N__35961\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__35961\,
            I => \N__35958\
        );

    \I__7407\ : Span4Mux_s2_h
    port map (
            O => \N__35958\,
            I => \N__35955\
        );

    \I__7406\ : Span4Mux_h
    port map (
            O => \N__35955\,
            I => \N__35952\
        );

    \I__7405\ : Span4Mux_h
    port map (
            O => \N__35952\,
            I => \N__35948\
        );

    \I__7404\ : InMux
    port map (
            O => \N__35951\,
            I => \N__35944\
        );

    \I__7403\ : Sp12to4
    port map (
            O => \N__35948\,
            I => \N__35941\
        );

    \I__7402\ : InMux
    port map (
            O => \N__35947\,
            I => \N__35938\
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__35944\,
            I => \N__35935\
        );

    \I__7400\ : Odrv12
    port map (
            O => \N__35941\,
            I => pin_out_4
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__35938\,
            I => pin_out_4
        );

    \I__7398\ : Odrv4
    port map (
            O => \N__35935\,
            I => pin_out_4
        );

    \I__7397\ : InMux
    port map (
            O => \N__35928\,
            I => \N__35925\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__35925\,
            I => \N__35921\
        );

    \I__7395\ : CascadeMux
    port map (
            O => \N__35924\,
            I => \N__35918\
        );

    \I__7394\ : Span4Mux_h
    port map (
            O => \N__35921\,
            I => \N__35915\
        );

    \I__7393\ : InMux
    port map (
            O => \N__35918\,
            I => \N__35912\
        );

    \I__7392\ : Odrv4
    port map (
            O => \N__35915\,
            I => \nx.n2609\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__35912\,
            I => \nx.n2609\
        );

    \I__7390\ : InMux
    port map (
            O => \N__35907\,
            I => \N__35903\
        );

    \I__7389\ : InMux
    port map (
            O => \N__35906\,
            I => \N__35900\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__35903\,
            I => \N__35896\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__35900\,
            I => \N__35893\
        );

    \I__7386\ : InMux
    port map (
            O => \N__35899\,
            I => \N__35890\
        );

    \I__7385\ : Span4Mux_v
    port map (
            O => \N__35896\,
            I => \N__35887\
        );

    \I__7384\ : Span4Mux_h
    port map (
            O => \N__35893\,
            I => \N__35882\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__35890\,
            I => \N__35882\
        );

    \I__7382\ : Sp12to4
    port map (
            O => \N__35887\,
            I => \N__35877\
        );

    \I__7381\ : Sp12to4
    port map (
            O => \N__35882\,
            I => \N__35874\
        );

    \I__7380\ : InMux
    port map (
            O => \N__35881\,
            I => \N__35871\
        );

    \I__7379\ : InMux
    port map (
            O => \N__35880\,
            I => \N__35868\
        );

    \I__7378\ : Span12Mux_h
    port map (
            O => \N__35877\,
            I => \N__35865\
        );

    \I__7377\ : Span12Mux_v
    port map (
            O => \N__35874\,
            I => \N__35862\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__35871\,
            I => \nx.bit_ctr_9\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__35868\,
            I => \nx.bit_ctr_9\
        );

    \I__7374\ : Odrv12
    port map (
            O => \N__35865\,
            I => \nx.bit_ctr_9\
        );

    \I__7373\ : Odrv12
    port map (
            O => \N__35862\,
            I => \nx.bit_ctr_9\
        );

    \I__7372\ : CascadeMux
    port map (
            O => \N__35853\,
            I => \nx.n2609_cascade_\
        );

    \I__7371\ : CascadeMux
    port map (
            O => \N__35850\,
            I => \nx.n28_adj_599_cascade_\
        );

    \I__7370\ : InMux
    port map (
            O => \N__35847\,
            I => \N__35844\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__35844\,
            I => \N__35841\
        );

    \I__7368\ : Span4Mux_h
    port map (
            O => \N__35841\,
            I => \N__35838\
        );

    \I__7367\ : Odrv4
    port map (
            O => \N__35838\,
            I => \nx.n35\
        );

    \I__7366\ : InMux
    port map (
            O => \N__35835\,
            I => \N__35832\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__35832\,
            I => \N__35829\
        );

    \I__7364\ : Odrv4
    port map (
            O => \N__35829\,
            I => \nx.n40\
        );

    \I__7363\ : InMux
    port map (
            O => \N__35826\,
            I => \N__35822\
        );

    \I__7362\ : CascadeMux
    port map (
            O => \N__35825\,
            I => \N__35818\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__35822\,
            I => \N__35815\
        );

    \I__7360\ : InMux
    port map (
            O => \N__35821\,
            I => \N__35812\
        );

    \I__7359\ : InMux
    port map (
            O => \N__35818\,
            I => \N__35809\
        );

    \I__7358\ : Odrv12
    port map (
            O => \N__35815\,
            I => \nx.n2608\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__35812\,
            I => \nx.n2608\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__35809\,
            I => \nx.n2608\
        );

    \I__7355\ : IoInMux
    port map (
            O => \N__35802\,
            I => \N__35797\
        );

    \I__7354\ : IoInMux
    port map (
            O => \N__35801\,
            I => \N__35790\
        );

    \I__7353\ : IoInMux
    port map (
            O => \N__35800\,
            I => \N__35787\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__35797\,
            I => \N__35784\
        );

    \I__7351\ : IoInMux
    port map (
            O => \N__35796\,
            I => \N__35779\
        );

    \I__7350\ : IoInMux
    port map (
            O => \N__35795\,
            I => \N__35776\
        );

    \I__7349\ : IoInMux
    port map (
            O => \N__35794\,
            I => \N__35773\
        );

    \I__7348\ : IoInMux
    port map (
            O => \N__35793\,
            I => \N__35769\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__35790\,
            I => \N__35761\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__35787\,
            I => \N__35761\
        );

    \I__7345\ : IoSpan4Mux
    port map (
            O => \N__35784\,
            I => \N__35761\
        );

    \I__7344\ : IoInMux
    port map (
            O => \N__35783\,
            I => \N__35758\
        );

    \I__7343\ : IoInMux
    port map (
            O => \N__35782\,
            I => \N__35755\
        );

    \I__7342\ : LocalMux
    port map (
            O => \N__35779\,
            I => \N__35750\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__35776\,
            I => \N__35750\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__35773\,
            I => \N__35747\
        );

    \I__7339\ : IoInMux
    port map (
            O => \N__35772\,
            I => \N__35744\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__35769\,
            I => \N__35741\
        );

    \I__7337\ : IoInMux
    port map (
            O => \N__35768\,
            I => \N__35738\
        );

    \I__7336\ : IoSpan4Mux
    port map (
            O => \N__35761\,
            I => \N__35726\
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__35758\,
            I => \N__35726\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__35755\,
            I => \N__35726\
        );

    \I__7333\ : IoSpan4Mux
    port map (
            O => \N__35750\,
            I => \N__35716\
        );

    \I__7332\ : IoSpan4Mux
    port map (
            O => \N__35747\,
            I => \N__35716\
        );

    \I__7331\ : LocalMux
    port map (
            O => \N__35744\,
            I => \N__35716\
        );

    \I__7330\ : IoSpan4Mux
    port map (
            O => \N__35741\,
            I => \N__35713\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__35738\,
            I => \N__35710\
        );

    \I__7328\ : IoInMux
    port map (
            O => \N__35737\,
            I => \N__35707\
        );

    \I__7327\ : IoInMux
    port map (
            O => \N__35736\,
            I => \N__35704\
        );

    \I__7326\ : IoInMux
    port map (
            O => \N__35735\,
            I => \N__35701\
        );

    \I__7325\ : IoInMux
    port map (
            O => \N__35734\,
            I => \N__35698\
        );

    \I__7324\ : IoInMux
    port map (
            O => \N__35733\,
            I => \N__35695\
        );

    \I__7323\ : IoSpan4Mux
    port map (
            O => \N__35726\,
            I => \N__35692\
        );

    \I__7322\ : IoInMux
    port map (
            O => \N__35725\,
            I => \N__35689\
        );

    \I__7321\ : IoInMux
    port map (
            O => \N__35724\,
            I => \N__35686\
        );

    \I__7320\ : IoInMux
    port map (
            O => \N__35723\,
            I => \N__35683\
        );

    \I__7319\ : IoSpan4Mux
    port map (
            O => \N__35716\,
            I => \N__35680\
        );

    \I__7318\ : IoSpan4Mux
    port map (
            O => \N__35713\,
            I => \N__35676\
        );

    \I__7317\ : IoSpan4Mux
    port map (
            O => \N__35710\,
            I => \N__35671\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__35707\,
            I => \N__35671\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__35704\,
            I => \N__35665\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__35701\,
            I => \N__35662\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__35698\,
            I => \N__35657\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__35695\,
            I => \N__35657\
        );

    \I__7311\ : IoSpan4Mux
    port map (
            O => \N__35692\,
            I => \N__35650\
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__35689\,
            I => \N__35650\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__35686\,
            I => \N__35650\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__35683\,
            I => \N__35647\
        );

    \I__7307\ : Span4Mux_s2_v
    port map (
            O => \N__35680\,
            I => \N__35644\
        );

    \I__7306\ : IoInMux
    port map (
            O => \N__35679\,
            I => \N__35641\
        );

    \I__7305\ : IoSpan4Mux
    port map (
            O => \N__35676\,
            I => \N__35636\
        );

    \I__7304\ : IoSpan4Mux
    port map (
            O => \N__35671\,
            I => \N__35636\
        );

    \I__7303\ : IoInMux
    port map (
            O => \N__35670\,
            I => \N__35633\
        );

    \I__7302\ : IoInMux
    port map (
            O => \N__35669\,
            I => \N__35630\
        );

    \I__7301\ : IoInMux
    port map (
            O => \N__35668\,
            I => \N__35627\
        );

    \I__7300\ : Span4Mux_s2_v
    port map (
            O => \N__35665\,
            I => \N__35624\
        );

    \I__7299\ : Span4Mux_s2_v
    port map (
            O => \N__35662\,
            I => \N__35621\
        );

    \I__7298\ : IoSpan4Mux
    port map (
            O => \N__35657\,
            I => \N__35618\
        );

    \I__7297\ : IoSpan4Mux
    port map (
            O => \N__35650\,
            I => \N__35615\
        );

    \I__7296\ : Span12Mux_s9_h
    port map (
            O => \N__35647\,
            I => \N__35612\
        );

    \I__7295\ : Span4Mux_v
    port map (
            O => \N__35644\,
            I => \N__35609\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__35641\,
            I => \N__35606\
        );

    \I__7293\ : Span4Mux_s2_h
    port map (
            O => \N__35636\,
            I => \N__35603\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__35633\,
            I => \N__35598\
        );

    \I__7291\ : LocalMux
    port map (
            O => \N__35630\,
            I => \N__35598\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__35627\,
            I => \N__35595\
        );

    \I__7289\ : Sp12to4
    port map (
            O => \N__35624\,
            I => \N__35592\
        );

    \I__7288\ : Sp12to4
    port map (
            O => \N__35621\,
            I => \N__35589\
        );

    \I__7287\ : Span4Mux_s3_h
    port map (
            O => \N__35618\,
            I => \N__35586\
        );

    \I__7286\ : Span4Mux_s2_h
    port map (
            O => \N__35615\,
            I => \N__35583\
        );

    \I__7285\ : Span12Mux_h
    port map (
            O => \N__35612\,
            I => \N__35580\
        );

    \I__7284\ : Sp12to4
    port map (
            O => \N__35609\,
            I => \N__35575\
        );

    \I__7283\ : Span12Mux_s6_v
    port map (
            O => \N__35606\,
            I => \N__35575\
        );

    \I__7282\ : Sp12to4
    port map (
            O => \N__35603\,
            I => \N__35572\
        );

    \I__7281\ : Sp12to4
    port map (
            O => \N__35598\,
            I => \N__35569\
        );

    \I__7280\ : Span12Mux_s9_h
    port map (
            O => \N__35595\,
            I => \N__35566\
        );

    \I__7279\ : Span12Mux_h
    port map (
            O => \N__35592\,
            I => \N__35561\
        );

    \I__7278\ : Span12Mux_s10_h
    port map (
            O => \N__35589\,
            I => \N__35561\
        );

    \I__7277\ : Sp12to4
    port map (
            O => \N__35586\,
            I => \N__35558\
        );

    \I__7276\ : Span4Mux_h
    port map (
            O => \N__35583\,
            I => \N__35555\
        );

    \I__7275\ : Span12Mux_v
    port map (
            O => \N__35580\,
            I => \N__35548\
        );

    \I__7274\ : Span12Mux_v
    port map (
            O => \N__35575\,
            I => \N__35548\
        );

    \I__7273\ : Span12Mux_s9_h
    port map (
            O => \N__35572\,
            I => \N__35548\
        );

    \I__7272\ : Span12Mux_v
    port map (
            O => \N__35569\,
            I => \N__35545\
        );

    \I__7271\ : Span12Mux_h
    port map (
            O => \N__35566\,
            I => \N__35538\
        );

    \I__7270\ : Span12Mux_v
    port map (
            O => \N__35561\,
            I => \N__35538\
        );

    \I__7269\ : Span12Mux_s10_h
    port map (
            O => \N__35558\,
            I => \N__35538\
        );

    \I__7268\ : Span4Mux_h
    port map (
            O => \N__35555\,
            I => \N__35535\
        );

    \I__7267\ : Odrv12
    port map (
            O => \N__35548\,
            I => pin_oe_22
        );

    \I__7266\ : Odrv12
    port map (
            O => \N__35545\,
            I => pin_oe_22
        );

    \I__7265\ : Odrv12
    port map (
            O => \N__35538\,
            I => pin_oe_22
        );

    \I__7264\ : Odrv4
    port map (
            O => \N__35535\,
            I => pin_oe_22
        );

    \I__7263\ : InMux
    port map (
            O => \N__35526\,
            I => \N__35522\
        );

    \I__7262\ : InMux
    port map (
            O => \N__35525\,
            I => \N__35519\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__35522\,
            I => \N__35514\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__35519\,
            I => \N__35514\
        );

    \I__7259\ : Span4Mux_h
    port map (
            O => \N__35514\,
            I => \N__35511\
        );

    \I__7258\ : Odrv4
    port map (
            O => \N__35511\,
            I => n6158
        );

    \I__7257\ : CascadeMux
    port map (
            O => \N__35508\,
            I => \N__35505\
        );

    \I__7256\ : InMux
    port map (
            O => \N__35505\,
            I => \N__35499\
        );

    \I__7255\ : InMux
    port map (
            O => \N__35504\,
            I => \N__35494\
        );

    \I__7254\ : InMux
    port map (
            O => \N__35503\,
            I => \N__35494\
        );

    \I__7253\ : InMux
    port map (
            O => \N__35502\,
            I => \N__35491\
        );

    \I__7252\ : LocalMux
    port map (
            O => \N__35499\,
            I => \N__35486\
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__35494\,
            I => \N__35486\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__35491\,
            I => \N__35483\
        );

    \I__7249\ : Span4Mux_h
    port map (
            O => \N__35486\,
            I => \N__35480\
        );

    \I__7248\ : Odrv4
    port map (
            O => \N__35483\,
            I => n8
        );

    \I__7247\ : Odrv4
    port map (
            O => \N__35480\,
            I => n8
        );

    \I__7246\ : CascadeMux
    port map (
            O => \N__35475\,
            I => \n22_adj_740_cascade_\
        );

    \I__7245\ : InMux
    port map (
            O => \N__35472\,
            I => \N__35468\
        );

    \I__7244\ : InMux
    port map (
            O => \N__35471\,
            I => \N__35465\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__35468\,
            I => \N__35460\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__35465\,
            I => \N__35460\
        );

    \I__7241\ : Span4Mux_h
    port map (
            O => \N__35460\,
            I => \N__35457\
        );

    \I__7240\ : Odrv4
    port map (
            O => \N__35457\,
            I => n5907
        );

    \I__7239\ : InMux
    port map (
            O => \N__35454\,
            I => \N__35451\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__35451\,
            I => n6162
        );

    \I__7237\ : CascadeMux
    port map (
            O => \N__35448\,
            I => \n6162_cascade_\
        );

    \I__7236\ : InMux
    port map (
            O => \N__35445\,
            I => \N__35442\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__35442\,
            I => n7278
        );

    \I__7234\ : InMux
    port map (
            O => \N__35439\,
            I => \N__35435\
        );

    \I__7233\ : CascadeMux
    port map (
            O => \N__35438\,
            I => \N__35432\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__35435\,
            I => \N__35429\
        );

    \I__7231\ : InMux
    port map (
            O => \N__35432\,
            I => \N__35426\
        );

    \I__7230\ : Span4Mux_v
    port map (
            O => \N__35429\,
            I => \N__35422\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__35426\,
            I => \N__35419\
        );

    \I__7228\ : CascadeMux
    port map (
            O => \N__35425\,
            I => \N__35416\
        );

    \I__7227\ : Span4Mux_h
    port map (
            O => \N__35422\,
            I => \N__35411\
        );

    \I__7226\ : Span4Mux_h
    port map (
            O => \N__35419\,
            I => \N__35411\
        );

    \I__7225\ : InMux
    port map (
            O => \N__35416\,
            I => \N__35408\
        );

    \I__7224\ : Odrv4
    port map (
            O => \N__35411\,
            I => \nx.n1704\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__35408\,
            I => \nx.n1704\
        );

    \I__7222\ : InMux
    port map (
            O => \N__35403\,
            I => \N__35400\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__35400\,
            I => \nx.n1771\
        );

    \I__7220\ : InMux
    port map (
            O => \N__35397\,
            I => \nx.n10620\
        );

    \I__7219\ : InMux
    port map (
            O => \N__35394\,
            I => \N__35387\
        );

    \I__7218\ : InMux
    port map (
            O => \N__35393\,
            I => \N__35387\
        );

    \I__7217\ : CascadeMux
    port map (
            O => \N__35392\,
            I => \N__35384\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__35387\,
            I => \N__35381\
        );

    \I__7215\ : InMux
    port map (
            O => \N__35384\,
            I => \N__35378\
        );

    \I__7214\ : Odrv4
    port map (
            O => \N__35381\,
            I => \nx.n1703\
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__35378\,
            I => \nx.n1703\
        );

    \I__7212\ : InMux
    port map (
            O => \N__35373\,
            I => \N__35370\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__35370\,
            I => \nx.n1770\
        );

    \I__7210\ : InMux
    port map (
            O => \N__35367\,
            I => \nx.n10621\
        );

    \I__7209\ : CascadeMux
    port map (
            O => \N__35364\,
            I => \N__35361\
        );

    \I__7208\ : InMux
    port map (
            O => \N__35361\,
            I => \N__35358\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__35358\,
            I => \N__35353\
        );

    \I__7206\ : InMux
    port map (
            O => \N__35357\,
            I => \N__35348\
        );

    \I__7205\ : InMux
    port map (
            O => \N__35356\,
            I => \N__35348\
        );

    \I__7204\ : Odrv4
    port map (
            O => \N__35353\,
            I => \nx.n1702\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__35348\,
            I => \nx.n1702\
        );

    \I__7202\ : CascadeMux
    port map (
            O => \N__35343\,
            I => \N__35340\
        );

    \I__7201\ : InMux
    port map (
            O => \N__35340\,
            I => \N__35337\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__35337\,
            I => \N__35334\
        );

    \I__7199\ : Span4Mux_v
    port map (
            O => \N__35334\,
            I => \N__35331\
        );

    \I__7198\ : Span4Mux_h
    port map (
            O => \N__35331\,
            I => \N__35328\
        );

    \I__7197\ : Odrv4
    port map (
            O => \N__35328\,
            I => \nx.n1769\
        );

    \I__7196\ : InMux
    port map (
            O => \N__35325\,
            I => \bfn_10_29_0_\
        );

    \I__7195\ : CascadeMux
    port map (
            O => \N__35322\,
            I => \N__35319\
        );

    \I__7194\ : InMux
    port map (
            O => \N__35319\,
            I => \N__35315\
        );

    \I__7193\ : InMux
    port map (
            O => \N__35318\,
            I => \N__35312\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__35315\,
            I => \N__35309\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__35312\,
            I => \N__35306\
        );

    \I__7190\ : Span4Mux_v
    port map (
            O => \N__35309\,
            I => \N__35301\
        );

    \I__7189\ : Span4Mux_v
    port map (
            O => \N__35306\,
            I => \N__35301\
        );

    \I__7188\ : Odrv4
    port map (
            O => \N__35301\,
            I => \nx.n1701\
        );

    \I__7187\ : InMux
    port map (
            O => \N__35298\,
            I => \N__35295\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__35295\,
            I => \N__35292\
        );

    \I__7185\ : Span4Mux_v
    port map (
            O => \N__35292\,
            I => \N__35289\
        );

    \I__7184\ : Odrv4
    port map (
            O => \N__35289\,
            I => \nx.n1768\
        );

    \I__7183\ : InMux
    port map (
            O => \N__35286\,
            I => \nx.n10623\
        );

    \I__7182\ : InMux
    port map (
            O => \N__35283\,
            I => \N__35280\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__35280\,
            I => \N__35275\
        );

    \I__7180\ : InMux
    port map (
            O => \N__35279\,
            I => \N__35272\
        );

    \I__7179\ : InMux
    port map (
            O => \N__35278\,
            I => \N__35269\
        );

    \I__7178\ : Odrv4
    port map (
            O => \N__35275\,
            I => \nx.n1700\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__35272\,
            I => \nx.n1700\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__35269\,
            I => \nx.n1700\
        );

    \I__7175\ : InMux
    port map (
            O => \N__35262\,
            I => \N__35259\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__35259\,
            I => \N__35256\
        );

    \I__7173\ : Odrv4
    port map (
            O => \N__35256\,
            I => \nx.n1767\
        );

    \I__7172\ : InMux
    port map (
            O => \N__35253\,
            I => \nx.n10624\
        );

    \I__7171\ : CascadeMux
    port map (
            O => \N__35250\,
            I => \N__35246\
        );

    \I__7170\ : CascadeMux
    port map (
            O => \N__35249\,
            I => \N__35243\
        );

    \I__7169\ : InMux
    port map (
            O => \N__35246\,
            I => \N__35239\
        );

    \I__7168\ : InMux
    port map (
            O => \N__35243\,
            I => \N__35234\
        );

    \I__7167\ : InMux
    port map (
            O => \N__35242\,
            I => \N__35234\
        );

    \I__7166\ : LocalMux
    port map (
            O => \N__35239\,
            I => \N__35231\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__35234\,
            I => \N__35228\
        );

    \I__7164\ : Span4Mux_h
    port map (
            O => \N__35231\,
            I => \N__35225\
        );

    \I__7163\ : Span4Mux_h
    port map (
            O => \N__35228\,
            I => \N__35222\
        );

    \I__7162\ : Odrv4
    port map (
            O => \N__35225\,
            I => \nx.n1699\
        );

    \I__7161\ : Odrv4
    port map (
            O => \N__35222\,
            I => \nx.n1699\
        );

    \I__7160\ : InMux
    port map (
            O => \N__35217\,
            I => \N__35214\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__35214\,
            I => \N__35211\
        );

    \I__7158\ : Odrv4
    port map (
            O => \N__35211\,
            I => \nx.n1766\
        );

    \I__7157\ : InMux
    port map (
            O => \N__35208\,
            I => \nx.n10625\
        );

    \I__7156\ : InMux
    port map (
            O => \N__35205\,
            I => \N__35201\
        );

    \I__7155\ : CascadeMux
    port map (
            O => \N__35204\,
            I => \N__35198\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__35201\,
            I => \N__35195\
        );

    \I__7153\ : InMux
    port map (
            O => \N__35198\,
            I => \N__35192\
        );

    \I__7152\ : Span4Mux_h
    port map (
            O => \N__35195\,
            I => \N__35189\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__35192\,
            I => \N__35186\
        );

    \I__7150\ : Span4Mux_v
    port map (
            O => \N__35189\,
            I => \N__35182\
        );

    \I__7149\ : Span4Mux_h
    port map (
            O => \N__35186\,
            I => \N__35179\
        );

    \I__7148\ : InMux
    port map (
            O => \N__35185\,
            I => \N__35176\
        );

    \I__7147\ : Odrv4
    port map (
            O => \N__35182\,
            I => \nx.n1698\
        );

    \I__7146\ : Odrv4
    port map (
            O => \N__35179\,
            I => \nx.n1698\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__35176\,
            I => \nx.n1698\
        );

    \I__7144\ : CascadeMux
    port map (
            O => \N__35169\,
            I => \N__35166\
        );

    \I__7143\ : InMux
    port map (
            O => \N__35166\,
            I => \N__35163\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__35163\,
            I => \N__35160\
        );

    \I__7141\ : Span4Mux_v
    port map (
            O => \N__35160\,
            I => \N__35157\
        );

    \I__7140\ : Odrv4
    port map (
            O => \N__35157\,
            I => \nx.n1765\
        );

    \I__7139\ : InMux
    port map (
            O => \N__35154\,
            I => \nx.n10626\
        );

    \I__7138\ : InMux
    port map (
            O => \N__35151\,
            I => \N__35142\
        );

    \I__7137\ : InMux
    port map (
            O => \N__35150\,
            I => \N__35137\
        );

    \I__7136\ : InMux
    port map (
            O => \N__35149\,
            I => \N__35137\
        );

    \I__7135\ : InMux
    port map (
            O => \N__35148\,
            I => \N__35134\
        );

    \I__7134\ : InMux
    port map (
            O => \N__35147\,
            I => \N__35129\
        );

    \I__7133\ : InMux
    port map (
            O => \N__35146\,
            I => \N__35129\
        );

    \I__7132\ : InMux
    port map (
            O => \N__35145\,
            I => \N__35122\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__35142\,
            I => \N__35115\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__35137\,
            I => \N__35115\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__35134\,
            I => \N__35115\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__35129\,
            I => \N__35112\
        );

    \I__7127\ : CascadeMux
    port map (
            O => \N__35128\,
            I => \N__35109\
        );

    \I__7126\ : InMux
    port map (
            O => \N__35127\,
            I => \N__35100\
        );

    \I__7125\ : InMux
    port map (
            O => \N__35126\,
            I => \N__35100\
        );

    \I__7124\ : InMux
    port map (
            O => \N__35125\,
            I => \N__35100\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__35122\,
            I => \N__35097\
        );

    \I__7122\ : Span4Mux_h
    port map (
            O => \N__35115\,
            I => \N__35094\
        );

    \I__7121\ : Span4Mux_h
    port map (
            O => \N__35112\,
            I => \N__35091\
        );

    \I__7120\ : InMux
    port map (
            O => \N__35109\,
            I => \N__35084\
        );

    \I__7119\ : InMux
    port map (
            O => \N__35108\,
            I => \N__35084\
        );

    \I__7118\ : InMux
    port map (
            O => \N__35107\,
            I => \N__35084\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__35100\,
            I => \nx.n1730\
        );

    \I__7116\ : Odrv4
    port map (
            O => \N__35097\,
            I => \nx.n1730\
        );

    \I__7115\ : Odrv4
    port map (
            O => \N__35094\,
            I => \nx.n1730\
        );

    \I__7114\ : Odrv4
    port map (
            O => \N__35091\,
            I => \nx.n1730\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__35084\,
            I => \nx.n1730\
        );

    \I__7112\ : CascadeMux
    port map (
            O => \N__35073\,
            I => \N__35070\
        );

    \I__7111\ : InMux
    port map (
            O => \N__35070\,
            I => \N__35067\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__35067\,
            I => \N__35064\
        );

    \I__7109\ : Span4Mux_h
    port map (
            O => \N__35064\,
            I => \N__35060\
        );

    \I__7108\ : InMux
    port map (
            O => \N__35063\,
            I => \N__35057\
        );

    \I__7107\ : Odrv4
    port map (
            O => \N__35060\,
            I => \nx.n1697\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__35057\,
            I => \nx.n1697\
        );

    \I__7105\ : InMux
    port map (
            O => \N__35052\,
            I => \nx.n10627\
        );

    \I__7104\ : CascadeMux
    port map (
            O => \N__35049\,
            I => \N__35046\
        );

    \I__7103\ : InMux
    port map (
            O => \N__35046\,
            I => \N__35042\
        );

    \I__7102\ : InMux
    port map (
            O => \N__35045\,
            I => \N__35039\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__35042\,
            I => \N__35036\
        );

    \I__7100\ : LocalMux
    port map (
            O => \N__35039\,
            I => \nx.n1796\
        );

    \I__7099\ : Odrv4
    port map (
            O => \N__35036\,
            I => \nx.n1796\
        );

    \I__7098\ : CascadeMux
    port map (
            O => \N__35031\,
            I => \N__35028\
        );

    \I__7097\ : InMux
    port map (
            O => \N__35028\,
            I => \N__35025\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__35025\,
            I => \N__35022\
        );

    \I__7095\ : Span4Mux_v
    port map (
            O => \N__35022\,
            I => \N__35019\
        );

    \I__7094\ : Odrv4
    port map (
            O => \N__35019\,
            I => \nx.n20_adj_680\
        );

    \I__7093\ : InMux
    port map (
            O => \N__35016\,
            I => \N__35013\
        );

    \I__7092\ : LocalMux
    port map (
            O => \N__35013\,
            I => \nx.n24_adj_685\
        );

    \I__7091\ : CascadeMux
    port map (
            O => \N__35010\,
            I => \nx.n1730_cascade_\
        );

    \I__7090\ : CascadeMux
    port map (
            O => \N__35007\,
            I => \N__35002\
        );

    \I__7089\ : InMux
    port map (
            O => \N__35006\,
            I => \N__34999\
        );

    \I__7088\ : CascadeMux
    port map (
            O => \N__35005\,
            I => \N__34996\
        );

    \I__7087\ : InMux
    port map (
            O => \N__35002\,
            I => \N__34993\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__34999\,
            I => \N__34990\
        );

    \I__7085\ : InMux
    port map (
            O => \N__34996\,
            I => \N__34987\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__34993\,
            I => \N__34982\
        );

    \I__7083\ : Span4Mux_h
    port map (
            O => \N__34990\,
            I => \N__34982\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__34987\,
            I => \nx.n1802\
        );

    \I__7081\ : Odrv4
    port map (
            O => \N__34982\,
            I => \nx.n1802\
        );

    \I__7080\ : InMux
    port map (
            O => \N__34977\,
            I => \N__34972\
        );

    \I__7079\ : InMux
    port map (
            O => \N__34976\,
            I => \N__34969\
        );

    \I__7078\ : InMux
    port map (
            O => \N__34975\,
            I => \N__34966\
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__34972\,
            I => \N__34962\
        );

    \I__7076\ : LocalMux
    port map (
            O => \N__34969\,
            I => \N__34959\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__34966\,
            I => \N__34956\
        );

    \I__7074\ : InMux
    port map (
            O => \N__34965\,
            I => \N__34953\
        );

    \I__7073\ : Span4Mux_s3_h
    port map (
            O => \N__34962\,
            I => \N__34943\
        );

    \I__7072\ : Span4Mux_v
    port map (
            O => \N__34959\,
            I => \N__34943\
        );

    \I__7071\ : Span4Mux_h
    port map (
            O => \N__34956\,
            I => \N__34943\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__34953\,
            I => \N__34943\
        );

    \I__7069\ : InMux
    port map (
            O => \N__34952\,
            I => \N__34940\
        );

    \I__7068\ : Span4Mux_h
    port map (
            O => \N__34943\,
            I => \N__34937\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__34940\,
            I => \nx.bit_ctr_18\
        );

    \I__7066\ : Odrv4
    port map (
            O => \N__34937\,
            I => \nx.bit_ctr_18\
        );

    \I__7065\ : InMux
    port map (
            O => \N__34932\,
            I => \N__34929\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__34929\,
            I => \N__34926\
        );

    \I__7063\ : Span4Mux_v
    port map (
            O => \N__34926\,
            I => \N__34923\
        );

    \I__7062\ : Odrv4
    port map (
            O => \N__34923\,
            I => \nx.n1777\
        );

    \I__7061\ : InMux
    port map (
            O => \N__34920\,
            I => \bfn_10_28_0_\
        );

    \I__7060\ : CascadeMux
    port map (
            O => \N__34917\,
            I => \N__34913\
        );

    \I__7059\ : CascadeMux
    port map (
            O => \N__34916\,
            I => \N__34909\
        );

    \I__7058\ : InMux
    port map (
            O => \N__34913\,
            I => \N__34906\
        );

    \I__7057\ : CascadeMux
    port map (
            O => \N__34912\,
            I => \N__34903\
        );

    \I__7056\ : InMux
    port map (
            O => \N__34909\,
            I => \N__34900\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__34906\,
            I => \N__34897\
        );

    \I__7054\ : InMux
    port map (
            O => \N__34903\,
            I => \N__34894\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__34900\,
            I => \nx.n1709\
        );

    \I__7052\ : Odrv12
    port map (
            O => \N__34897\,
            I => \nx.n1709\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__34894\,
            I => \nx.n1709\
        );

    \I__7050\ : InMux
    port map (
            O => \N__34887\,
            I => \N__34884\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__34884\,
            I => \N__34881\
        );

    \I__7048\ : Span4Mux_v
    port map (
            O => \N__34881\,
            I => \N__34878\
        );

    \I__7047\ : Span4Mux_h
    port map (
            O => \N__34878\,
            I => \N__34875\
        );

    \I__7046\ : Odrv4
    port map (
            O => \N__34875\,
            I => \nx.n1776\
        );

    \I__7045\ : InMux
    port map (
            O => \N__34872\,
            I => \nx.n10615\
        );

    \I__7044\ : CascadeMux
    port map (
            O => \N__34869\,
            I => \N__34864\
        );

    \I__7043\ : InMux
    port map (
            O => \N__34868\,
            I => \N__34861\
        );

    \I__7042\ : CascadeMux
    port map (
            O => \N__34867\,
            I => \N__34858\
        );

    \I__7041\ : InMux
    port map (
            O => \N__34864\,
            I => \N__34855\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__34861\,
            I => \N__34852\
        );

    \I__7039\ : InMux
    port map (
            O => \N__34858\,
            I => \N__34849\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__34855\,
            I => \N__34846\
        );

    \I__7037\ : Span4Mux_v
    port map (
            O => \N__34852\,
            I => \N__34841\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__34849\,
            I => \N__34841\
        );

    \I__7035\ : Span4Mux_v
    port map (
            O => \N__34846\,
            I => \N__34838\
        );

    \I__7034\ : Span4Mux_h
    port map (
            O => \N__34841\,
            I => \N__34835\
        );

    \I__7033\ : Odrv4
    port map (
            O => \N__34838\,
            I => \nx.n1708\
        );

    \I__7032\ : Odrv4
    port map (
            O => \N__34835\,
            I => \nx.n1708\
        );

    \I__7031\ : InMux
    port map (
            O => \N__34830\,
            I => \N__34827\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__34827\,
            I => \N__34824\
        );

    \I__7029\ : Odrv4
    port map (
            O => \N__34824\,
            I => \nx.n1775\
        );

    \I__7028\ : InMux
    port map (
            O => \N__34821\,
            I => \nx.n10616\
        );

    \I__7027\ : CascadeMux
    port map (
            O => \N__34818\,
            I => \N__34815\
        );

    \I__7026\ : InMux
    port map (
            O => \N__34815\,
            I => \N__34811\
        );

    \I__7025\ : InMux
    port map (
            O => \N__34814\,
            I => \N__34808\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__34811\,
            I => \nx.n1707\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__34808\,
            I => \nx.n1707\
        );

    \I__7022\ : InMux
    port map (
            O => \N__34803\,
            I => \N__34800\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__34800\,
            I => \nx.n1774\
        );

    \I__7020\ : InMux
    port map (
            O => \N__34797\,
            I => \nx.n10617\
        );

    \I__7019\ : CascadeMux
    port map (
            O => \N__34794\,
            I => \N__34791\
        );

    \I__7018\ : InMux
    port map (
            O => \N__34791\,
            I => \N__34788\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__34788\,
            I => \N__34784\
        );

    \I__7016\ : InMux
    port map (
            O => \N__34787\,
            I => \N__34781\
        );

    \I__7015\ : Span4Mux_v
    port map (
            O => \N__34784\,
            I => \N__34775\
        );

    \I__7014\ : LocalMux
    port map (
            O => \N__34781\,
            I => \N__34775\
        );

    \I__7013\ : InMux
    port map (
            O => \N__34780\,
            I => \N__34772\
        );

    \I__7012\ : Span4Mux_h
    port map (
            O => \N__34775\,
            I => \N__34769\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__34772\,
            I => \nx.n1706\
        );

    \I__7010\ : Odrv4
    port map (
            O => \N__34769\,
            I => \nx.n1706\
        );

    \I__7009\ : InMux
    port map (
            O => \N__34764\,
            I => \N__34761\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__34761\,
            I => \N__34758\
        );

    \I__7007\ : Span4Mux_h
    port map (
            O => \N__34758\,
            I => \N__34755\
        );

    \I__7006\ : Odrv4
    port map (
            O => \N__34755\,
            I => \nx.n1773\
        );

    \I__7005\ : InMux
    port map (
            O => \N__34752\,
            I => \nx.n10618\
        );

    \I__7004\ : CascadeMux
    port map (
            O => \N__34749\,
            I => \N__34746\
        );

    \I__7003\ : InMux
    port map (
            O => \N__34746\,
            I => \N__34743\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__34743\,
            I => \N__34738\
        );

    \I__7001\ : CascadeMux
    port map (
            O => \N__34742\,
            I => \N__34735\
        );

    \I__7000\ : InMux
    port map (
            O => \N__34741\,
            I => \N__34732\
        );

    \I__6999\ : Span4Mux_h
    port map (
            O => \N__34738\,
            I => \N__34729\
        );

    \I__6998\ : InMux
    port map (
            O => \N__34735\,
            I => \N__34726\
        );

    \I__6997\ : LocalMux
    port map (
            O => \N__34732\,
            I => \N__34723\
        );

    \I__6996\ : Odrv4
    port map (
            O => \N__34729\,
            I => \nx.n1705\
        );

    \I__6995\ : LocalMux
    port map (
            O => \N__34726\,
            I => \nx.n1705\
        );

    \I__6994\ : Odrv4
    port map (
            O => \N__34723\,
            I => \nx.n1705\
        );

    \I__6993\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34713\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__34713\,
            I => \N__34710\
        );

    \I__6991\ : Span4Mux_h
    port map (
            O => \N__34710\,
            I => \N__34707\
        );

    \I__6990\ : Odrv4
    port map (
            O => \N__34707\,
            I => \nx.n1772\
        );

    \I__6989\ : InMux
    port map (
            O => \N__34704\,
            I => \nx.n10619\
        );

    \I__6988\ : CascadeMux
    port map (
            O => \N__34701\,
            I => \nx.n2097_cascade_\
        );

    \I__6987\ : InMux
    port map (
            O => \N__34698\,
            I => \N__34695\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__34695\,
            I => \nx.n27_adj_671\
        );

    \I__6985\ : CascadeMux
    port map (
            O => \N__34692\,
            I => \N__34688\
        );

    \I__6984\ : CascadeMux
    port map (
            O => \N__34691\,
            I => \N__34684\
        );

    \I__6983\ : InMux
    port map (
            O => \N__34688\,
            I => \N__34681\
        );

    \I__6982\ : InMux
    port map (
            O => \N__34687\,
            I => \N__34678\
        );

    \I__6981\ : InMux
    port map (
            O => \N__34684\,
            I => \N__34675\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__34681\,
            I => \N__34672\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__34678\,
            I => \N__34667\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__34675\,
            I => \N__34667\
        );

    \I__6977\ : Span4Mux_h
    port map (
            O => \N__34672\,
            I => \N__34662\
        );

    \I__6976\ : Span4Mux_v
    port map (
            O => \N__34667\,
            I => \N__34662\
        );

    \I__6975\ : Odrv4
    port map (
            O => \N__34662\,
            I => \nx.n2007\
        );

    \I__6974\ : InMux
    port map (
            O => \N__34659\,
            I => \N__34655\
        );

    \I__6973\ : CascadeMux
    port map (
            O => \N__34658\,
            I => \N__34652\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__34655\,
            I => \N__34649\
        );

    \I__6971\ : InMux
    port map (
            O => \N__34652\,
            I => \N__34646\
        );

    \I__6970\ : Span4Mux_v
    port map (
            O => \N__34649\,
            I => \N__34640\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__34646\,
            I => \N__34640\
        );

    \I__6968\ : InMux
    port map (
            O => \N__34645\,
            I => \N__34637\
        );

    \I__6967\ : Span4Mux_h
    port map (
            O => \N__34640\,
            I => \N__34634\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__34637\,
            I => \N__34631\
        );

    \I__6965\ : Odrv4
    port map (
            O => \N__34634\,
            I => \nx.n2002\
        );

    \I__6964\ : Odrv12
    port map (
            O => \N__34631\,
            I => \nx.n2002\
        );

    \I__6963\ : InMux
    port map (
            O => \N__34626\,
            I => \N__34623\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__34623\,
            I => \N__34620\
        );

    \I__6961\ : Odrv4
    port map (
            O => \N__34620\,
            I => \nx.n22_adj_662\
        );

    \I__6960\ : CascadeMux
    port map (
            O => \N__34617\,
            I => \N__34614\
        );

    \I__6959\ : InMux
    port map (
            O => \N__34614\,
            I => \N__34609\
        );

    \I__6958\ : InMux
    port map (
            O => \N__34613\,
            I => \N__34606\
        );

    \I__6957\ : InMux
    port map (
            O => \N__34612\,
            I => \N__34603\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__34609\,
            I => \N__34598\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__34606\,
            I => \N__34598\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__34603\,
            I => \nx.n1803\
        );

    \I__6953\ : Odrv12
    port map (
            O => \N__34598\,
            I => \nx.n1803\
        );

    \I__6952\ : CascadeMux
    port map (
            O => \N__34593\,
            I => \nx.n22_adj_673_cascade_\
        );

    \I__6951\ : InMux
    port map (
            O => \N__34590\,
            I => \N__34587\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__34587\,
            I => \N__34584\
        );

    \I__6949\ : Span4Mux_h
    port map (
            O => \N__34584\,
            I => \N__34581\
        );

    \I__6948\ : Odrv4
    port map (
            O => \N__34581\,
            I => \nx.n16_adj_672\
        );

    \I__6947\ : InMux
    port map (
            O => \N__34578\,
            I => \N__34574\
        );

    \I__6946\ : CascadeMux
    port map (
            O => \N__34577\,
            I => \N__34571\
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__34574\,
            I => \N__34567\
        );

    \I__6944\ : InMux
    port map (
            O => \N__34571\,
            I => \N__34564\
        );

    \I__6943\ : InMux
    port map (
            O => \N__34570\,
            I => \N__34561\
        );

    \I__6942\ : Odrv4
    port map (
            O => \N__34567\,
            I => \nx.n1798\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__34564\,
            I => \nx.n1798\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__34561\,
            I => \nx.n1798\
        );

    \I__6939\ : CascadeMux
    port map (
            O => \N__34554\,
            I => \N__34551\
        );

    \I__6938\ : InMux
    port map (
            O => \N__34551\,
            I => \N__34547\
        );

    \I__6937\ : InMux
    port map (
            O => \N__34550\,
            I => \N__34544\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__34547\,
            I => \N__34541\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__34544\,
            I => \N__34536\
        );

    \I__6934\ : Span4Mux_h
    port map (
            O => \N__34541\,
            I => \N__34536\
        );

    \I__6933\ : Odrv4
    port map (
            O => \N__34536\,
            I => \nx.n1608\
        );

    \I__6932\ : CascadeMux
    port map (
            O => \N__34533\,
            I => \N__34530\
        );

    \I__6931\ : InMux
    port map (
            O => \N__34530\,
            I => \N__34527\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__34527\,
            I => \N__34524\
        );

    \I__6929\ : Span4Mux_h
    port map (
            O => \N__34524\,
            I => \N__34521\
        );

    \I__6928\ : Odrv4
    port map (
            O => \N__34521\,
            I => \nx.n1675\
        );

    \I__6927\ : InMux
    port map (
            O => \N__34518\,
            I => \N__34512\
        );

    \I__6926\ : CascadeMux
    port map (
            O => \N__34517\,
            I => \N__34508\
        );

    \I__6925\ : InMux
    port map (
            O => \N__34516\,
            I => \N__34505\
        );

    \I__6924\ : CascadeMux
    port map (
            O => \N__34515\,
            I => \N__34501\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__34512\,
            I => \N__34496\
        );

    \I__6922\ : InMux
    port map (
            O => \N__34511\,
            I => \N__34491\
        );

    \I__6921\ : InMux
    port map (
            O => \N__34508\,
            I => \N__34491\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__34505\,
            I => \N__34488\
        );

    \I__6919\ : InMux
    port map (
            O => \N__34504\,
            I => \N__34483\
        );

    \I__6918\ : InMux
    port map (
            O => \N__34501\,
            I => \N__34483\
        );

    \I__6917\ : CascadeMux
    port map (
            O => \N__34500\,
            I => \N__34477\
        );

    \I__6916\ : InMux
    port map (
            O => \N__34499\,
            I => \N__34473\
        );

    \I__6915\ : Span4Mux_v
    port map (
            O => \N__34496\,
            I => \N__34468\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__34491\,
            I => \N__34468\
        );

    \I__6913\ : Span4Mux_h
    port map (
            O => \N__34488\,
            I => \N__34463\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__34483\,
            I => \N__34463\
        );

    \I__6911\ : InMux
    port map (
            O => \N__34482\,
            I => \N__34458\
        );

    \I__6910\ : InMux
    port map (
            O => \N__34481\,
            I => \N__34458\
        );

    \I__6909\ : InMux
    port map (
            O => \N__34480\,
            I => \N__34455\
        );

    \I__6908\ : InMux
    port map (
            O => \N__34477\,
            I => \N__34450\
        );

    \I__6907\ : InMux
    port map (
            O => \N__34476\,
            I => \N__34450\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__34473\,
            I => \nx.n1631\
        );

    \I__6905\ : Odrv4
    port map (
            O => \N__34468\,
            I => \nx.n1631\
        );

    \I__6904\ : Odrv4
    port map (
            O => \N__34463\,
            I => \nx.n1631\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__34458\,
            I => \nx.n1631\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__34455\,
            I => \nx.n1631\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__34450\,
            I => \nx.n1631\
        );

    \I__6900\ : CascadeMux
    port map (
            O => \N__34437\,
            I => \nx.n1707_cascade_\
        );

    \I__6899\ : InMux
    port map (
            O => \N__34434\,
            I => \N__34429\
        );

    \I__6898\ : InMux
    port map (
            O => \N__34433\,
            I => \N__34426\
        );

    \I__6897\ : CascadeMux
    port map (
            O => \N__34432\,
            I => \N__34423\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__34429\,
            I => \N__34420\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__34426\,
            I => \N__34417\
        );

    \I__6894\ : InMux
    port map (
            O => \N__34423\,
            I => \N__34414\
        );

    \I__6893\ : Span4Mux_v
    port map (
            O => \N__34420\,
            I => \N__34411\
        );

    \I__6892\ : Odrv4
    port map (
            O => \N__34417\,
            I => \nx.n1806\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__34414\,
            I => \nx.n1806\
        );

    \I__6890\ : Odrv4
    port map (
            O => \N__34411\,
            I => \nx.n1806\
        );

    \I__6889\ : InMux
    port map (
            O => \N__34404\,
            I => \N__34401\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__34401\,
            I => \nx.n2074\
        );

    \I__6887\ : InMux
    port map (
            O => \N__34398\,
            I => \N__34395\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__34395\,
            I => \nx.n2064\
        );

    \I__6885\ : CascadeMux
    port map (
            O => \N__34392\,
            I => \N__34389\
        );

    \I__6884\ : InMux
    port map (
            O => \N__34389\,
            I => \N__34385\
        );

    \I__6883\ : CascadeMux
    port map (
            O => \N__34388\,
            I => \N__34382\
        );

    \I__6882\ : LocalMux
    port map (
            O => \N__34385\,
            I => \N__34379\
        );

    \I__6881\ : InMux
    port map (
            O => \N__34382\,
            I => \N__34376\
        );

    \I__6880\ : Span4Mux_v
    port map (
            O => \N__34379\,
            I => \N__34370\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__34376\,
            I => \N__34370\
        );

    \I__6878\ : InMux
    port map (
            O => \N__34375\,
            I => \N__34367\
        );

    \I__6877\ : Span4Mux_h
    port map (
            O => \N__34370\,
            I => \N__34364\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__34367\,
            I => \N__34361\
        );

    \I__6875\ : Odrv4
    port map (
            O => \N__34364\,
            I => \nx.n1997\
        );

    \I__6874\ : Odrv12
    port map (
            O => \N__34361\,
            I => \nx.n1997\
        );

    \I__6873\ : InMux
    port map (
            O => \N__34356\,
            I => \N__34353\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__34353\,
            I => \nx.n2062\
        );

    \I__6871\ : CascadeMux
    port map (
            O => \N__34350\,
            I => \N__34347\
        );

    \I__6870\ : InMux
    port map (
            O => \N__34347\,
            I => \N__34343\
        );

    \I__6869\ : CascadeMux
    port map (
            O => \N__34346\,
            I => \N__34340\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__34343\,
            I => \N__34336\
        );

    \I__6867\ : InMux
    port map (
            O => \N__34340\,
            I => \N__34333\
        );

    \I__6866\ : CascadeMux
    port map (
            O => \N__34339\,
            I => \N__34330\
        );

    \I__6865\ : Span4Mux_v
    port map (
            O => \N__34336\,
            I => \N__34325\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__34333\,
            I => \N__34325\
        );

    \I__6863\ : InMux
    port map (
            O => \N__34330\,
            I => \N__34322\
        );

    \I__6862\ : Span4Mux_h
    port map (
            O => \N__34325\,
            I => \N__34319\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__34322\,
            I => \N__34316\
        );

    \I__6860\ : Odrv4
    port map (
            O => \N__34319\,
            I => \nx.n1995\
        );

    \I__6859\ : Odrv12
    port map (
            O => \N__34316\,
            I => \nx.n1995\
        );

    \I__6858\ : InMux
    port map (
            O => \N__34311\,
            I => \N__34308\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__34308\,
            I => \N__34305\
        );

    \I__6856\ : Odrv4
    port map (
            O => \N__34305\,
            I => \nx.n26_adj_667\
        );

    \I__6855\ : CascadeMux
    port map (
            O => \N__34302\,
            I => \nx.n30_adj_668_cascade_\
        );

    \I__6854\ : InMux
    port map (
            O => \N__34299\,
            I => \N__34296\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__34296\,
            I => \N__34293\
        );

    \I__6852\ : Odrv4
    port map (
            O => \N__34293\,
            I => \nx.n28_adj_669\
        );

    \I__6851\ : CascadeMux
    port map (
            O => \N__34290\,
            I => \N__34286\
        );

    \I__6850\ : InMux
    port map (
            O => \N__34289\,
            I => \N__34283\
        );

    \I__6849\ : InMux
    port map (
            O => \N__34286\,
            I => \N__34280\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__34283\,
            I => \N__34277\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__34280\,
            I => \N__34273\
        );

    \I__6846\ : Span4Mux_v
    port map (
            O => \N__34277\,
            I => \N__34270\
        );

    \I__6845\ : InMux
    port map (
            O => \N__34276\,
            I => \N__34267\
        );

    \I__6844\ : Span4Mux_h
    port map (
            O => \N__34273\,
            I => \N__34264\
        );

    \I__6843\ : Odrv4
    port map (
            O => \N__34270\,
            I => \nx.n2008\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__34267\,
            I => \nx.n2008\
        );

    \I__6841\ : Odrv4
    port map (
            O => \N__34264\,
            I => \nx.n2008\
        );

    \I__6840\ : CascadeMux
    port map (
            O => \N__34257\,
            I => \N__34254\
        );

    \I__6839\ : InMux
    port map (
            O => \N__34254\,
            I => \N__34251\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__34251\,
            I => \nx.n2075\
        );

    \I__6837\ : CascadeMux
    port map (
            O => \N__34248\,
            I => \nx.n2107_cascade_\
        );

    \I__6836\ : InMux
    port map (
            O => \N__34245\,
            I => \N__34242\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__34242\,
            I => \nx.n29_adj_670\
        );

    \I__6834\ : InMux
    port map (
            O => \N__34239\,
            I => \N__34236\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__34236\,
            I => \nx.n2065\
        );

    \I__6832\ : InMux
    port map (
            O => \N__34233\,
            I => \N__34228\
        );

    \I__6831\ : CascadeMux
    port map (
            O => \N__34232\,
            I => \N__34225\
        );

    \I__6830\ : CascadeMux
    port map (
            O => \N__34231\,
            I => \N__34222\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__34228\,
            I => \N__34219\
        );

    \I__6828\ : InMux
    port map (
            O => \N__34225\,
            I => \N__34216\
        );

    \I__6827\ : InMux
    port map (
            O => \N__34222\,
            I => \N__34213\
        );

    \I__6826\ : Span4Mux_h
    port map (
            O => \N__34219\,
            I => \N__34210\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__34216\,
            I => \N__34205\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__34213\,
            I => \N__34205\
        );

    \I__6823\ : Span4Mux_v
    port map (
            O => \N__34210\,
            I => \N__34200\
        );

    \I__6822\ : Span4Mux_v
    port map (
            O => \N__34205\,
            I => \N__34200\
        );

    \I__6821\ : Odrv4
    port map (
            O => \N__34200\,
            I => \nx.n1998\
        );

    \I__6820\ : CascadeMux
    port map (
            O => \N__34197\,
            I => \N__34186\
        );

    \I__6819\ : CascadeMux
    port map (
            O => \N__34196\,
            I => \N__34180\
        );

    \I__6818\ : CascadeMux
    port map (
            O => \N__34195\,
            I => \N__34177\
        );

    \I__6817\ : InMux
    port map (
            O => \N__34194\,
            I => \N__34172\
        );

    \I__6816\ : InMux
    port map (
            O => \N__34193\,
            I => \N__34172\
        );

    \I__6815\ : InMux
    port map (
            O => \N__34192\,
            I => \N__34169\
        );

    \I__6814\ : CascadeMux
    port map (
            O => \N__34191\,
            I => \N__34165\
        );

    \I__6813\ : CascadeMux
    port map (
            O => \N__34190\,
            I => \N__34161\
        );

    \I__6812\ : InMux
    port map (
            O => \N__34189\,
            I => \N__34156\
        );

    \I__6811\ : InMux
    port map (
            O => \N__34186\,
            I => \N__34143\
        );

    \I__6810\ : InMux
    port map (
            O => \N__34185\,
            I => \N__34143\
        );

    \I__6809\ : InMux
    port map (
            O => \N__34184\,
            I => \N__34143\
        );

    \I__6808\ : InMux
    port map (
            O => \N__34183\,
            I => \N__34143\
        );

    \I__6807\ : InMux
    port map (
            O => \N__34180\,
            I => \N__34143\
        );

    \I__6806\ : InMux
    port map (
            O => \N__34177\,
            I => \N__34143\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__34172\,
            I => \N__34138\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__34169\,
            I => \N__34138\
        );

    \I__6803\ : InMux
    port map (
            O => \N__34168\,
            I => \N__34131\
        );

    \I__6802\ : InMux
    port map (
            O => \N__34165\,
            I => \N__34131\
        );

    \I__6801\ : InMux
    port map (
            O => \N__34164\,
            I => \N__34131\
        );

    \I__6800\ : InMux
    port map (
            O => \N__34161\,
            I => \N__34124\
        );

    \I__6799\ : InMux
    port map (
            O => \N__34160\,
            I => \N__34124\
        );

    \I__6798\ : InMux
    port map (
            O => \N__34159\,
            I => \N__34124\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__34156\,
            I => \nx.n2027\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__34143\,
            I => \nx.n2027\
        );

    \I__6795\ : Odrv4
    port map (
            O => \N__34138\,
            I => \nx.n2027\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__34131\,
            I => \nx.n2027\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__34124\,
            I => \nx.n2027\
        );

    \I__6792\ : CascadeMux
    port map (
            O => \N__34113\,
            I => \nx.n2394_cascade_\
        );

    \I__6791\ : InMux
    port map (
            O => \N__34110\,
            I => \N__34107\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__34107\,
            I => \nx.n2077\
        );

    \I__6789\ : InMux
    port map (
            O => \N__34104\,
            I => \N__34101\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__34101\,
            I => \nx.n2070\
        );

    \I__6787\ : CascadeMux
    port map (
            O => \N__34098\,
            I => \N__34095\
        );

    \I__6786\ : InMux
    port map (
            O => \N__34095\,
            I => \N__34092\
        );

    \I__6785\ : LocalMux
    port map (
            O => \N__34092\,
            I => \nx.n2069\
        );

    \I__6784\ : InMux
    port map (
            O => \N__34089\,
            I => \N__34086\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__34086\,
            I => \nx.n2076\
        );

    \I__6782\ : InMux
    port map (
            O => \N__34083\,
            I => \N__34080\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__34080\,
            I => \N__34077\
        );

    \I__6780\ : Span4Mux_v
    port map (
            O => \N__34077\,
            I => \N__34071\
        );

    \I__6779\ : InMux
    port map (
            O => \N__34076\,
            I => \N__34068\
        );

    \I__6778\ : InMux
    port map (
            O => \N__34075\,
            I => \N__34065\
        );

    \I__6777\ : InMux
    port map (
            O => \N__34074\,
            I => \N__34061\
        );

    \I__6776\ : Sp12to4
    port map (
            O => \N__34071\,
            I => \N__34054\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__34068\,
            I => \N__34054\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__34065\,
            I => \N__34054\
        );

    \I__6773\ : InMux
    port map (
            O => \N__34064\,
            I => \N__34051\
        );

    \I__6772\ : LocalMux
    port map (
            O => \N__34061\,
            I => \N__34046\
        );

    \I__6771\ : Span12Mux_h
    port map (
            O => \N__34054\,
            I => \N__34046\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__34051\,
            I => \nx.bit_ctr_15\
        );

    \I__6769\ : Odrv12
    port map (
            O => \N__34046\,
            I => \nx.bit_ctr_15\
        );

    \I__6768\ : CascadeMux
    port map (
            O => \N__34041\,
            I => \N__34036\
        );

    \I__6767\ : InMux
    port map (
            O => \N__34040\,
            I => \N__34031\
        );

    \I__6766\ : InMux
    port map (
            O => \N__34039\,
            I => \N__34031\
        );

    \I__6765\ : InMux
    port map (
            O => \N__34036\,
            I => \N__34028\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__34031\,
            I => \N__34023\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__34028\,
            I => \N__34023\
        );

    \I__6762\ : Span4Mux_h
    port map (
            O => \N__34023\,
            I => \N__34020\
        );

    \I__6761\ : Odrv4
    port map (
            O => \N__34020\,
            I => \nx.n2003\
        );

    \I__6760\ : CascadeMux
    port map (
            O => \N__34017\,
            I => \N__34012\
        );

    \I__6759\ : CascadeMux
    port map (
            O => \N__34016\,
            I => \N__34009\
        );

    \I__6758\ : InMux
    port map (
            O => \N__34015\,
            I => \N__34004\
        );

    \I__6757\ : InMux
    port map (
            O => \N__34012\,
            I => \N__34004\
        );

    \I__6756\ : InMux
    port map (
            O => \N__34009\,
            I => \N__34001\
        );

    \I__6755\ : LocalMux
    port map (
            O => \N__34004\,
            I => \N__33996\
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__34001\,
            I => \N__33996\
        );

    \I__6753\ : Span4Mux_h
    port map (
            O => \N__33996\,
            I => \N__33993\
        );

    \I__6752\ : Odrv4
    port map (
            O => \N__33993\,
            I => \nx.n2009\
        );

    \I__6751\ : InMux
    port map (
            O => \N__33990\,
            I => \N__33987\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__33987\,
            I => \nx.n27_adj_665\
        );

    \I__6749\ : InMux
    port map (
            O => \N__33984\,
            I => \N__33981\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__33981\,
            I => \nx.n36\
        );

    \I__6747\ : InMux
    port map (
            O => \N__33978\,
            I => \N__33975\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__33975\,
            I => \N__33972\
        );

    \I__6745\ : Span4Mux_h
    port map (
            O => \N__33972\,
            I => \N__33969\
        );

    \I__6744\ : Odrv4
    port map (
            O => \N__33969\,
            I => \nx.n41\
        );

    \I__6743\ : InMux
    port map (
            O => \N__33966\,
            I => \N__33963\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__33963\,
            I => \nx.n2656\
        );

    \I__6741\ : CascadeMux
    port map (
            O => \N__33960\,
            I => \nx.n31_adj_655_cascade_\
        );

    \I__6740\ : InMux
    port map (
            O => \N__33957\,
            I => \N__33954\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__33954\,
            I => \N__33951\
        );

    \I__6738\ : Span4Mux_h
    port map (
            O => \N__33951\,
            I => \N__33948\
        );

    \I__6737\ : Span4Mux_v
    port map (
            O => \N__33948\,
            I => \N__33945\
        );

    \I__6736\ : Odrv4
    port map (
            O => \N__33945\,
            I => \nx.n24_adj_654\
        );

    \I__6735\ : CascadeMux
    port map (
            O => \N__33942\,
            I => \nx.n36_adj_656_cascade_\
        );

    \I__6734\ : InMux
    port map (
            O => \N__33939\,
            I => \N__33936\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__33936\,
            I => \N__33933\
        );

    \I__6732\ : Span4Mux_h
    port map (
            O => \N__33933\,
            I => \N__33930\
        );

    \I__6731\ : Odrv4
    port map (
            O => \N__33930\,
            I => \nx.n33_adj_659\
        );

    \I__6730\ : CascadeMux
    port map (
            O => \N__33927\,
            I => \nx.n2423_cascade_\
        );

    \I__6729\ : CascadeMux
    port map (
            O => \N__33924\,
            I => \nx.n2491_cascade_\
        );

    \I__6728\ : InMux
    port map (
            O => \N__33921\,
            I => \nx.n10788\
        );

    \I__6727\ : InMux
    port map (
            O => \N__33918\,
            I => \nx.n10789\
        );

    \I__6726\ : CascadeMux
    port map (
            O => \N__33915\,
            I => \N__33912\
        );

    \I__6725\ : InMux
    port map (
            O => \N__33912\,
            I => \N__33909\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__33909\,
            I => \nx.n2660\
        );

    \I__6723\ : CascadeMux
    port map (
            O => \N__33906\,
            I => \N__33903\
        );

    \I__6722\ : InMux
    port map (
            O => \N__33903\,
            I => \N__33899\
        );

    \I__6721\ : CascadeMux
    port map (
            O => \N__33902\,
            I => \N__33896\
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__33899\,
            I => \N__33893\
        );

    \I__6719\ : InMux
    port map (
            O => \N__33896\,
            I => \N__33890\
        );

    \I__6718\ : Span4Mux_v
    port map (
            O => \N__33893\,
            I => \N__33885\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__33890\,
            I => \N__33885\
        );

    \I__6716\ : Span4Mux_h
    port map (
            O => \N__33885\,
            I => \N__33881\
        );

    \I__6715\ : InMux
    port map (
            O => \N__33884\,
            I => \N__33878\
        );

    \I__6714\ : Odrv4
    port map (
            O => \N__33881\,
            I => \nx.n2692\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__33878\,
            I => \nx.n2692\
        );

    \I__6712\ : CascadeMux
    port map (
            O => \N__33873\,
            I => \nx.n34_adj_603_cascade_\
        );

    \I__6711\ : CascadeMux
    port map (
            O => \N__33870\,
            I => \nx.n39_cascade_\
        );

    \I__6710\ : CascadeMux
    port map (
            O => \N__33867\,
            I => \nx.n2621_cascade_\
        );

    \I__6709\ : InMux
    port map (
            O => \N__33864\,
            I => \N__33861\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__33861\,
            I => \nx.n2661\
        );

    \I__6707\ : CascadeMux
    port map (
            O => \N__33858\,
            I => \N__33854\
        );

    \I__6706\ : InMux
    port map (
            O => \N__33857\,
            I => \N__33850\
        );

    \I__6705\ : InMux
    port map (
            O => \N__33854\,
            I => \N__33847\
        );

    \I__6704\ : InMux
    port map (
            O => \N__33853\,
            I => \N__33844\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__33850\,
            I => \N__33841\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__33847\,
            I => \N__33838\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__33844\,
            I => \N__33835\
        );

    \I__6700\ : Span4Mux_v
    port map (
            O => \N__33841\,
            I => \N__33830\
        );

    \I__6699\ : Span4Mux_v
    port map (
            O => \N__33838\,
            I => \N__33830\
        );

    \I__6698\ : Span4Mux_h
    port map (
            O => \N__33835\,
            I => \N__33827\
        );

    \I__6697\ : Odrv4
    port map (
            O => \N__33830\,
            I => \nx.n2693\
        );

    \I__6696\ : Odrv4
    port map (
            O => \N__33827\,
            I => \nx.n2693\
        );

    \I__6695\ : InMux
    port map (
            O => \N__33822\,
            I => \N__33819\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__33819\,
            I => \N__33816\
        );

    \I__6693\ : Odrv4
    port map (
            O => \N__33816\,
            I => \nx.n2667\
        );

    \I__6692\ : CascadeMux
    port map (
            O => \N__33813\,
            I => \N__33810\
        );

    \I__6691\ : InMux
    port map (
            O => \N__33810\,
            I => \N__33806\
        );

    \I__6690\ : CascadeMux
    port map (
            O => \N__33809\,
            I => \N__33803\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__33806\,
            I => \N__33800\
        );

    \I__6688\ : InMux
    port map (
            O => \N__33803\,
            I => \N__33797\
        );

    \I__6687\ : Span4Mux_h
    port map (
            O => \N__33800\,
            I => \N__33792\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__33797\,
            I => \N__33792\
        );

    \I__6685\ : Odrv4
    port map (
            O => \N__33792\,
            I => \nx.n2699\
        );

    \I__6684\ : CascadeMux
    port map (
            O => \N__33789\,
            I => \N__33786\
        );

    \I__6683\ : InMux
    port map (
            O => \N__33786\,
            I => \N__33783\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__33783\,
            I => \N__33780\
        );

    \I__6681\ : Span4Mux_h
    port map (
            O => \N__33780\,
            I => \N__33776\
        );

    \I__6680\ : InMux
    port map (
            O => \N__33779\,
            I => \N__33773\
        );

    \I__6679\ : Odrv4
    port map (
            O => \N__33776\,
            I => \nx.n2687\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__33773\,
            I => \nx.n2687\
        );

    \I__6677\ : CascadeMux
    port map (
            O => \N__33768\,
            I => \nx.n2699_cascade_\
        );

    \I__6676\ : CascadeMux
    port map (
            O => \N__33765\,
            I => \N__33762\
        );

    \I__6675\ : InMux
    port map (
            O => \N__33762\,
            I => \N__33759\
        );

    \I__6674\ : LocalMux
    port map (
            O => \N__33759\,
            I => \nx.n2665\
        );

    \I__6673\ : InMux
    port map (
            O => \N__33756\,
            I => \nx.n10779\
        );

    \I__6672\ : InMux
    port map (
            O => \N__33753\,
            I => \N__33750\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__33750\,
            I => \N__33747\
        );

    \I__6670\ : Span4Mux_v
    port map (
            O => \N__33747\,
            I => \N__33744\
        );

    \I__6669\ : Span4Mux_h
    port map (
            O => \N__33744\,
            I => \N__33741\
        );

    \I__6668\ : Odrv4
    port map (
            O => \N__33741\,
            I => \nx.n2664\
        );

    \I__6667\ : InMux
    port map (
            O => \N__33738\,
            I => \nx.n10780\
        );

    \I__6666\ : CascadeMux
    port map (
            O => \N__33735\,
            I => \N__33732\
        );

    \I__6665\ : InMux
    port map (
            O => \N__33732\,
            I => \N__33729\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__33729\,
            I => \nx.n2663\
        );

    \I__6663\ : InMux
    port map (
            O => \N__33726\,
            I => \nx.n10781\
        );

    \I__6662\ : CascadeMux
    port map (
            O => \N__33723\,
            I => \N__33720\
        );

    \I__6661\ : InMux
    port map (
            O => \N__33720\,
            I => \N__33716\
        );

    \I__6660\ : InMux
    port map (
            O => \N__33719\,
            I => \N__33713\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__33716\,
            I => \N__33710\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__33713\,
            I => \N__33707\
        );

    \I__6657\ : Span4Mux_h
    port map (
            O => \N__33710\,
            I => \N__33704\
        );

    \I__6656\ : Odrv4
    port map (
            O => \N__33707\,
            I => \nx.n2595\
        );

    \I__6655\ : Odrv4
    port map (
            O => \N__33704\,
            I => \nx.n2595\
        );

    \I__6654\ : InMux
    port map (
            O => \N__33699\,
            I => \N__33696\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__33696\,
            I => \nx.n2662\
        );

    \I__6652\ : InMux
    port map (
            O => \N__33693\,
            I => \nx.n10782\
        );

    \I__6651\ : InMux
    port map (
            O => \N__33690\,
            I => \bfn_10_19_0_\
        );

    \I__6650\ : InMux
    port map (
            O => \N__33687\,
            I => \nx.n10784\
        );

    \I__6649\ : CascadeMux
    port map (
            O => \N__33684\,
            I => \N__33681\
        );

    \I__6648\ : InMux
    port map (
            O => \N__33681\,
            I => \N__33677\
        );

    \I__6647\ : InMux
    port map (
            O => \N__33680\,
            I => \N__33674\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__33677\,
            I => \nx.n2592\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__33674\,
            I => \nx.n2592\
        );

    \I__6644\ : InMux
    port map (
            O => \N__33669\,
            I => \N__33666\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__33666\,
            I => \nx.n2659\
        );

    \I__6642\ : InMux
    port map (
            O => \N__33663\,
            I => \nx.n10785\
        );

    \I__6641\ : InMux
    port map (
            O => \N__33660\,
            I => \N__33657\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__33657\,
            I => \nx.n2658\
        );

    \I__6639\ : InMux
    port map (
            O => \N__33654\,
            I => \nx.n10786\
        );

    \I__6638\ : InMux
    port map (
            O => \N__33651\,
            I => \N__33648\
        );

    \I__6637\ : LocalMux
    port map (
            O => \N__33648\,
            I => \nx.n2657\
        );

    \I__6636\ : InMux
    port map (
            O => \N__33645\,
            I => \nx.n10787\
        );

    \I__6635\ : InMux
    port map (
            O => \N__33642\,
            I => \nx.n10771\
        );

    \I__6634\ : InMux
    port map (
            O => \N__33639\,
            I => \N__33636\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__33636\,
            I => \N__33633\
        );

    \I__6632\ : Odrv4
    port map (
            O => \N__33633\,
            I => \nx.n2672\
        );

    \I__6631\ : InMux
    port map (
            O => \N__33630\,
            I => \nx.n10772\
        );

    \I__6630\ : InMux
    port map (
            O => \N__33627\,
            I => \N__33624\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__33624\,
            I => \N__33621\
        );

    \I__6628\ : Odrv4
    port map (
            O => \N__33621\,
            I => \nx.n2671\
        );

    \I__6627\ : InMux
    port map (
            O => \N__33618\,
            I => \nx.n10773\
        );

    \I__6626\ : CascadeMux
    port map (
            O => \N__33615\,
            I => \N__33612\
        );

    \I__6625\ : InMux
    port map (
            O => \N__33612\,
            I => \N__33609\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__33609\,
            I => \N__33606\
        );

    \I__6623\ : Odrv4
    port map (
            O => \N__33606\,
            I => \nx.n2670\
        );

    \I__6622\ : InMux
    port map (
            O => \N__33603\,
            I => \nx.n10774\
        );

    \I__6621\ : InMux
    port map (
            O => \N__33600\,
            I => \N__33597\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__33597\,
            I => \N__33594\
        );

    \I__6619\ : Odrv4
    port map (
            O => \N__33594\,
            I => \nx.n2669\
        );

    \I__6618\ : InMux
    port map (
            O => \N__33591\,
            I => \bfn_10_18_0_\
        );

    \I__6617\ : CascadeMux
    port map (
            O => \N__33588\,
            I => \N__33585\
        );

    \I__6616\ : InMux
    port map (
            O => \N__33585\,
            I => \N__33582\
        );

    \I__6615\ : LocalMux
    port map (
            O => \N__33582\,
            I => \N__33579\
        );

    \I__6614\ : Odrv12
    port map (
            O => \N__33579\,
            I => \nx.n2668\
        );

    \I__6613\ : InMux
    port map (
            O => \N__33576\,
            I => \nx.n10776\
        );

    \I__6612\ : InMux
    port map (
            O => \N__33573\,
            I => \nx.n10777\
        );

    \I__6611\ : InMux
    port map (
            O => \N__33570\,
            I => \N__33567\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__33567\,
            I => \nx.n2666\
        );

    \I__6609\ : InMux
    port map (
            O => \N__33564\,
            I => \nx.n10778\
        );

    \I__6608\ : IoInMux
    port map (
            O => \N__33561\,
            I => \N__33558\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__33558\,
            I => \N__33555\
        );

    \I__6606\ : Span4Mux_s2_h
    port map (
            O => \N__33555\,
            I => \N__33552\
        );

    \I__6605\ : Span4Mux_v
    port map (
            O => \N__33552\,
            I => \N__33549\
        );

    \I__6604\ : Sp12to4
    port map (
            O => \N__33549\,
            I => \N__33545\
        );

    \I__6603\ : CascadeMux
    port map (
            O => \N__33548\,
            I => \N__33542\
        );

    \I__6602\ : Span12Mux_s9_h
    port map (
            O => \N__33545\,
            I => \N__33538\
        );

    \I__6601\ : InMux
    port map (
            O => \N__33542\,
            I => \N__33535\
        );

    \I__6600\ : InMux
    port map (
            O => \N__33541\,
            I => \N__33532\
        );

    \I__6599\ : Odrv12
    port map (
            O => \N__33538\,
            I => pin_out_6
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__33535\,
            I => pin_out_6
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__33532\,
            I => pin_out_6
        );

    \I__6596\ : InMux
    port map (
            O => \N__33525\,
            I => \N__33522\
        );

    \I__6595\ : LocalMux
    port map (
            O => \N__33522\,
            I => \N__33519\
        );

    \I__6594\ : Odrv4
    port map (
            O => \N__33519\,
            I => n7262
        );

    \I__6593\ : IoInMux
    port map (
            O => \N__33516\,
            I => \N__33513\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__33513\,
            I => \N__33510\
        );

    \I__6591\ : Span12Mux_s1_h
    port map (
            O => \N__33510\,
            I => \N__33506\
        );

    \I__6590\ : CascadeMux
    port map (
            O => \N__33509\,
            I => \N__33503\
        );

    \I__6589\ : Span12Mux_v
    port map (
            O => \N__33506\,
            I => \N__33499\
        );

    \I__6588\ : InMux
    port map (
            O => \N__33503\,
            I => \N__33496\
        );

    \I__6587\ : InMux
    port map (
            O => \N__33502\,
            I => \N__33493\
        );

    \I__6586\ : Odrv12
    port map (
            O => \N__33499\,
            I => pin_out_7
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__33496\,
            I => pin_out_7
        );

    \I__6584\ : LocalMux
    port map (
            O => \N__33493\,
            I => pin_out_7
        );

    \I__6583\ : InMux
    port map (
            O => \N__33486\,
            I => \N__33483\
        );

    \I__6582\ : LocalMux
    port map (
            O => \N__33483\,
            I => n8_adj_780
        );

    \I__6581\ : CascadeMux
    port map (
            O => \N__33480\,
            I => \n8_adj_780_cascade_\
        );

    \I__6580\ : InMux
    port map (
            O => \N__33477\,
            I => \N__33474\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__33474\,
            I => n7274
        );

    \I__6578\ : InMux
    port map (
            O => \N__33471\,
            I => \N__33468\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__33468\,
            I => \N__33465\
        );

    \I__6576\ : Odrv4
    port map (
            O => \N__33465\,
            I => \nx.n2677\
        );

    \I__6575\ : InMux
    port map (
            O => \N__33462\,
            I => \bfn_10_17_0_\
        );

    \I__6574\ : CascadeMux
    port map (
            O => \N__33459\,
            I => \N__33456\
        );

    \I__6573\ : InMux
    port map (
            O => \N__33456\,
            I => \N__33453\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__33453\,
            I => \N__33450\
        );

    \I__6571\ : Span4Mux_h
    port map (
            O => \N__33450\,
            I => \N__33447\
        );

    \I__6570\ : Odrv4
    port map (
            O => \N__33447\,
            I => \nx.n2676\
        );

    \I__6569\ : InMux
    port map (
            O => \N__33444\,
            I => \nx.n10768\
        );

    \I__6568\ : InMux
    port map (
            O => \N__33441\,
            I => \N__33438\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__33438\,
            I => \N__33435\
        );

    \I__6566\ : Span4Mux_v
    port map (
            O => \N__33435\,
            I => \N__33432\
        );

    \I__6565\ : Odrv4
    port map (
            O => \N__33432\,
            I => \nx.n2675\
        );

    \I__6564\ : InMux
    port map (
            O => \N__33429\,
            I => \nx.n10769\
        );

    \I__6563\ : InMux
    port map (
            O => \N__33426\,
            I => \N__33423\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__33423\,
            I => \N__33420\
        );

    \I__6561\ : Span4Mux_h
    port map (
            O => \N__33420\,
            I => \N__33417\
        );

    \I__6560\ : Odrv4
    port map (
            O => \N__33417\,
            I => \nx.n2674\
        );

    \I__6559\ : InMux
    port map (
            O => \N__33414\,
            I => \nx.n10770\
        );

    \I__6558\ : InMux
    port map (
            O => \N__33411\,
            I => \N__33408\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__33408\,
            I => \N__33405\
        );

    \I__6556\ : Span4Mux_h
    port map (
            O => \N__33405\,
            I => \N__33402\
        );

    \I__6555\ : Odrv4
    port map (
            O => \N__33402\,
            I => \nx.n1668\
        );

    \I__6554\ : CascadeMux
    port map (
            O => \N__33399\,
            I => \N__33396\
        );

    \I__6553\ : InMux
    port map (
            O => \N__33396\,
            I => \N__33393\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__33393\,
            I => \N__33389\
        );

    \I__6551\ : CascadeMux
    port map (
            O => \N__33392\,
            I => \N__33386\
        );

    \I__6550\ : Span4Mux_h
    port map (
            O => \N__33389\,
            I => \N__33382\
        );

    \I__6549\ : InMux
    port map (
            O => \N__33386\,
            I => \N__33379\
        );

    \I__6548\ : InMux
    port map (
            O => \N__33385\,
            I => \N__33376\
        );

    \I__6547\ : Odrv4
    port map (
            O => \N__33382\,
            I => \nx.n1601\
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__33379\,
            I => \nx.n1601\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__33376\,
            I => \nx.n1601\
        );

    \I__6544\ : InMux
    port map (
            O => \N__33369\,
            I => \N__33366\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__33366\,
            I => \N__33363\
        );

    \I__6542\ : Span4Mux_h
    port map (
            O => \N__33363\,
            I => \N__33359\
        );

    \I__6541\ : CascadeMux
    port map (
            O => \N__33362\,
            I => \N__33356\
        );

    \I__6540\ : IoSpan4Mux
    port map (
            O => \N__33359\,
            I => \N__33353\
        );

    \I__6539\ : InMux
    port map (
            O => \N__33356\,
            I => \N__33350\
        );

    \I__6538\ : Span4Mux_s1_v
    port map (
            O => \N__33353\,
            I => \N__33345\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__33350\,
            I => \N__33345\
        );

    \I__6536\ : Span4Mux_h
    port map (
            O => \N__33345\,
            I => \N__33342\
        );

    \I__6535\ : Odrv4
    port map (
            O => \N__33342\,
            I => \nx.n1509\
        );

    \I__6534\ : CascadeMux
    port map (
            O => \N__33339\,
            I => \N__33336\
        );

    \I__6533\ : InMux
    port map (
            O => \N__33336\,
            I => \N__33333\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__33333\,
            I => \N__33330\
        );

    \I__6531\ : Span4Mux_h
    port map (
            O => \N__33330\,
            I => \N__33327\
        );

    \I__6530\ : Odrv4
    port map (
            O => \N__33327\,
            I => \nx.n1576\
        );

    \I__6529\ : CascadeMux
    port map (
            O => \N__33324\,
            I => \nx.n1608_cascade_\
        );

    \I__6528\ : InMux
    port map (
            O => \N__33321\,
            I => \N__33318\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__33318\,
            I => \N__33315\
        );

    \I__6526\ : Odrv4
    port map (
            O => \N__33315\,
            I => \nx.n18\
        );

    \I__6525\ : InMux
    port map (
            O => \N__33312\,
            I => \N__33309\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__33309\,
            I => \N__33305\
        );

    \I__6523\ : CascadeMux
    port map (
            O => \N__33308\,
            I => \N__33302\
        );

    \I__6522\ : Span4Mux_v
    port map (
            O => \N__33305\,
            I => \N__33299\
        );

    \I__6521\ : InMux
    port map (
            O => \N__33302\,
            I => \N__33296\
        );

    \I__6520\ : Odrv4
    port map (
            O => \N__33299\,
            I => \nx.n1506\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__33296\,
            I => \nx.n1506\
        );

    \I__6518\ : CascadeMux
    port map (
            O => \N__33291\,
            I => \N__33288\
        );

    \I__6517\ : InMux
    port map (
            O => \N__33288\,
            I => \N__33285\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__33285\,
            I => \N__33282\
        );

    \I__6515\ : Span4Mux_h
    port map (
            O => \N__33282\,
            I => \N__33279\
        );

    \I__6514\ : Odrv4
    port map (
            O => \N__33279\,
            I => \nx.n1573\
        );

    \I__6513\ : CascadeMux
    port map (
            O => \N__33276\,
            I => \N__33267\
        );

    \I__6512\ : CascadeMux
    port map (
            O => \N__33275\,
            I => \N__33264\
        );

    \I__6511\ : CascadeMux
    port map (
            O => \N__33274\,
            I => \N__33259\
        );

    \I__6510\ : CascadeMux
    port map (
            O => \N__33273\,
            I => \N__33256\
        );

    \I__6509\ : CascadeMux
    port map (
            O => \N__33272\,
            I => \N__33252\
        );

    \I__6508\ : InMux
    port map (
            O => \N__33271\,
            I => \N__33246\
        );

    \I__6507\ : InMux
    port map (
            O => \N__33270\,
            I => \N__33246\
        );

    \I__6506\ : InMux
    port map (
            O => \N__33267\,
            I => \N__33243\
        );

    \I__6505\ : InMux
    port map (
            O => \N__33264\,
            I => \N__33236\
        );

    \I__6504\ : InMux
    port map (
            O => \N__33263\,
            I => \N__33236\
        );

    \I__6503\ : InMux
    port map (
            O => \N__33262\,
            I => \N__33236\
        );

    \I__6502\ : InMux
    port map (
            O => \N__33259\,
            I => \N__33231\
        );

    \I__6501\ : InMux
    port map (
            O => \N__33256\,
            I => \N__33231\
        );

    \I__6500\ : InMux
    port map (
            O => \N__33255\,
            I => \N__33224\
        );

    \I__6499\ : InMux
    port map (
            O => \N__33252\,
            I => \N__33224\
        );

    \I__6498\ : InMux
    port map (
            O => \N__33251\,
            I => \N__33224\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__33246\,
            I => \N__33221\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__33243\,
            I => \N__33218\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__33236\,
            I => \nx.n1532\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__33231\,
            I => \nx.n1532\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__33224\,
            I => \nx.n1532\
        );

    \I__6492\ : Odrv4
    port map (
            O => \N__33221\,
            I => \nx.n1532\
        );

    \I__6491\ : Odrv12
    port map (
            O => \N__33218\,
            I => \nx.n1532\
        );

    \I__6490\ : CascadeMux
    port map (
            O => \N__33207\,
            I => \N__33204\
        );

    \I__6489\ : InMux
    port map (
            O => \N__33204\,
            I => \N__33200\
        );

    \I__6488\ : InMux
    port map (
            O => \N__33203\,
            I => \N__33197\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__33200\,
            I => \N__33193\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__33197\,
            I => \N__33190\
        );

    \I__6485\ : InMux
    port map (
            O => \N__33196\,
            I => \N__33187\
        );

    \I__6484\ : Span4Mux_s3_v
    port map (
            O => \N__33193\,
            I => \N__33184\
        );

    \I__6483\ : Odrv4
    port map (
            O => \N__33190\,
            I => \nx.n1605\
        );

    \I__6482\ : LocalMux
    port map (
            O => \N__33187\,
            I => \nx.n1605\
        );

    \I__6481\ : Odrv4
    port map (
            O => \N__33184\,
            I => \nx.n1605\
        );

    \I__6480\ : InMux
    port map (
            O => \N__33177\,
            I => \N__33173\
        );

    \I__6479\ : CascadeMux
    port map (
            O => \N__33176\,
            I => \N__33169\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__33173\,
            I => \N__33166\
        );

    \I__6477\ : InMux
    port map (
            O => \N__33172\,
            I => \N__33163\
        );

    \I__6476\ : InMux
    port map (
            O => \N__33169\,
            I => \N__33160\
        );

    \I__6475\ : Odrv12
    port map (
            O => \N__33166\,
            I => \nx.n1604\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__33163\,
            I => \nx.n1604\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__33160\,
            I => \nx.n1604\
        );

    \I__6472\ : CascadeMux
    port map (
            O => \N__33153\,
            I => \N__33150\
        );

    \I__6471\ : InMux
    port map (
            O => \N__33150\,
            I => \N__33147\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__33147\,
            I => \N__33144\
        );

    \I__6469\ : Span4Mux_h
    port map (
            O => \N__33144\,
            I => \N__33141\
        );

    \I__6468\ : Odrv4
    port map (
            O => \N__33141\,
            I => \nx.n1671\
        );

    \I__6467\ : InMux
    port map (
            O => \N__33138\,
            I => \N__33134\
        );

    \I__6466\ : CascadeMux
    port map (
            O => \N__33137\,
            I => \N__33131\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__33134\,
            I => \N__33128\
        );

    \I__6464\ : InMux
    port map (
            O => \N__33131\,
            I => \N__33125\
        );

    \I__6463\ : Odrv4
    port map (
            O => \N__33128\,
            I => \nx.n1606\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__33125\,
            I => \nx.n1606\
        );

    \I__6461\ : InMux
    port map (
            O => \N__33120\,
            I => \N__33117\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__33117\,
            I => \N__33114\
        );

    \I__6459\ : Span4Mux_h
    port map (
            O => \N__33114\,
            I => \N__33111\
        );

    \I__6458\ : Odrv4
    port map (
            O => \N__33111\,
            I => \nx.n1673\
        );

    \I__6457\ : CascadeMux
    port map (
            O => \N__33108\,
            I => \n21_cascade_\
        );

    \I__6456\ : InMux
    port map (
            O => \N__33105\,
            I => \N__33102\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__33102\,
            I => \N__33099\
        );

    \I__6454\ : Span4Mux_h
    port map (
            O => \N__33099\,
            I => \N__33095\
        );

    \I__6453\ : InMux
    port map (
            O => \N__33098\,
            I => \N__33092\
        );

    \I__6452\ : Odrv4
    port map (
            O => \N__33095\,
            I => n6150
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__33092\,
            I => n6150
        );

    \I__6450\ : InMux
    port map (
            O => \N__33087\,
            I => \N__33084\
        );

    \I__6449\ : LocalMux
    port map (
            O => \N__33084\,
            I => \N__33081\
        );

    \I__6448\ : Odrv4
    port map (
            O => \N__33081\,
            I => \nx.n1870\
        );

    \I__6447\ : InMux
    port map (
            O => \N__33078\,
            I => \nx.n10634\
        );

    \I__6446\ : InMux
    port map (
            O => \N__33075\,
            I => \N__33072\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__33072\,
            I => \N__33069\
        );

    \I__6444\ : Odrv4
    port map (
            O => \N__33069\,
            I => \nx.n1869\
        );

    \I__6443\ : InMux
    port map (
            O => \N__33066\,
            I => \bfn_9_28_0_\
        );

    \I__6442\ : InMux
    port map (
            O => \N__33063\,
            I => \N__33059\
        );

    \I__6441\ : CascadeMux
    port map (
            O => \N__33062\,
            I => \N__33056\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__33059\,
            I => \N__33053\
        );

    \I__6439\ : InMux
    port map (
            O => \N__33056\,
            I => \N__33050\
        );

    \I__6438\ : Span4Mux_h
    port map (
            O => \N__33053\,
            I => \N__33047\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__33050\,
            I => \N__33044\
        );

    \I__6436\ : Odrv4
    port map (
            O => \N__33047\,
            I => \nx.n1801\
        );

    \I__6435\ : Odrv4
    port map (
            O => \N__33044\,
            I => \nx.n1801\
        );

    \I__6434\ : CascadeMux
    port map (
            O => \N__33039\,
            I => \N__33036\
        );

    \I__6433\ : InMux
    port map (
            O => \N__33036\,
            I => \N__33033\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__33033\,
            I => \N__33030\
        );

    \I__6431\ : Odrv4
    port map (
            O => \N__33030\,
            I => \nx.n1868\
        );

    \I__6430\ : InMux
    port map (
            O => \N__33027\,
            I => \nx.n10636\
        );

    \I__6429\ : CascadeMux
    port map (
            O => \N__33024\,
            I => \N__33021\
        );

    \I__6428\ : InMux
    port map (
            O => \N__33021\,
            I => \N__33017\
        );

    \I__6427\ : InMux
    port map (
            O => \N__33020\,
            I => \N__33013\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__33017\,
            I => \N__33010\
        );

    \I__6425\ : InMux
    port map (
            O => \N__33016\,
            I => \N__33007\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__33013\,
            I => \nx.n1800\
        );

    \I__6423\ : Odrv4
    port map (
            O => \N__33010\,
            I => \nx.n1800\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__33007\,
            I => \nx.n1800\
        );

    \I__6421\ : CascadeMux
    port map (
            O => \N__33000\,
            I => \N__32997\
        );

    \I__6420\ : InMux
    port map (
            O => \N__32997\,
            I => \N__32994\
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__32994\,
            I => \N__32991\
        );

    \I__6418\ : Span4Mux_h
    port map (
            O => \N__32991\,
            I => \N__32988\
        );

    \I__6417\ : Odrv4
    port map (
            O => \N__32988\,
            I => \nx.n1867\
        );

    \I__6416\ : InMux
    port map (
            O => \N__32985\,
            I => \nx.n10637\
        );

    \I__6415\ : InMux
    port map (
            O => \N__32982\,
            I => \N__32979\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__32979\,
            I => \N__32975\
        );

    \I__6413\ : InMux
    port map (
            O => \N__32978\,
            I => \N__32972\
        );

    \I__6412\ : Odrv4
    port map (
            O => \N__32975\,
            I => \nx.n1799\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__32972\,
            I => \nx.n1799\
        );

    \I__6410\ : InMux
    port map (
            O => \N__32967\,
            I => \N__32964\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__32964\,
            I => \N__32961\
        );

    \I__6408\ : Odrv4
    port map (
            O => \N__32961\,
            I => \nx.n1866\
        );

    \I__6407\ : InMux
    port map (
            O => \N__32958\,
            I => \nx.n10638\
        );

    \I__6406\ : InMux
    port map (
            O => \N__32955\,
            I => \N__32952\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__32952\,
            I => \N__32949\
        );

    \I__6404\ : Span4Mux_h
    port map (
            O => \N__32949\,
            I => \N__32946\
        );

    \I__6403\ : Odrv4
    port map (
            O => \N__32946\,
            I => \nx.n1865\
        );

    \I__6402\ : InMux
    port map (
            O => \N__32943\,
            I => \nx.n10639\
        );

    \I__6401\ : CascadeMux
    port map (
            O => \N__32940\,
            I => \N__32937\
        );

    \I__6400\ : InMux
    port map (
            O => \N__32937\,
            I => \N__32934\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__32934\,
            I => \N__32930\
        );

    \I__6398\ : InMux
    port map (
            O => \N__32933\,
            I => \N__32927\
        );

    \I__6397\ : Odrv4
    port map (
            O => \N__32930\,
            I => \nx.n1797\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__32927\,
            I => \nx.n1797\
        );

    \I__6395\ : InMux
    port map (
            O => \N__32922\,
            I => \N__32919\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__32919\,
            I => \N__32916\
        );

    \I__6393\ : Odrv4
    port map (
            O => \N__32916\,
            I => \nx.n1864\
        );

    \I__6392\ : InMux
    port map (
            O => \N__32913\,
            I => \nx.n10640\
        );

    \I__6391\ : CascadeMux
    port map (
            O => \N__32910\,
            I => \N__32907\
        );

    \I__6390\ : InMux
    port map (
            O => \N__32907\,
            I => \N__32904\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__32904\,
            I => \N__32893\
        );

    \I__6388\ : InMux
    port map (
            O => \N__32903\,
            I => \N__32888\
        );

    \I__6387\ : InMux
    port map (
            O => \N__32902\,
            I => \N__32888\
        );

    \I__6386\ : CascadeMux
    port map (
            O => \N__32901\,
            I => \N__32884\
        );

    \I__6385\ : CascadeMux
    port map (
            O => \N__32900\,
            I => \N__32879\
        );

    \I__6384\ : CascadeMux
    port map (
            O => \N__32899\,
            I => \N__32875\
        );

    \I__6383\ : InMux
    port map (
            O => \N__32898\,
            I => \N__32867\
        );

    \I__6382\ : InMux
    port map (
            O => \N__32897\,
            I => \N__32867\
        );

    \I__6381\ : InMux
    port map (
            O => \N__32896\,
            I => \N__32867\
        );

    \I__6380\ : Span4Mux_v
    port map (
            O => \N__32893\,
            I => \N__32862\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__32888\,
            I => \N__32862\
        );

    \I__6378\ : InMux
    port map (
            O => \N__32887\,
            I => \N__32859\
        );

    \I__6377\ : InMux
    port map (
            O => \N__32884\,
            I => \N__32854\
        );

    \I__6376\ : InMux
    port map (
            O => \N__32883\,
            I => \N__32854\
        );

    \I__6375\ : InMux
    port map (
            O => \N__32882\,
            I => \N__32851\
        );

    \I__6374\ : InMux
    port map (
            O => \N__32879\,
            I => \N__32842\
        );

    \I__6373\ : InMux
    port map (
            O => \N__32878\,
            I => \N__32842\
        );

    \I__6372\ : InMux
    port map (
            O => \N__32875\,
            I => \N__32842\
        );

    \I__6371\ : InMux
    port map (
            O => \N__32874\,
            I => \N__32842\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__32867\,
            I => \N__32839\
        );

    \I__6369\ : Span4Mux_h
    port map (
            O => \N__32862\,
            I => \N__32836\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__32859\,
            I => \nx.n1829\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__32854\,
            I => \nx.n1829\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__32851\,
            I => \nx.n1829\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__32842\,
            I => \nx.n1829\
        );

    \I__6364\ : Odrv4
    port map (
            O => \N__32839\,
            I => \nx.n1829\
        );

    \I__6363\ : Odrv4
    port map (
            O => \N__32836\,
            I => \nx.n1829\
        );

    \I__6362\ : InMux
    port map (
            O => \N__32823\,
            I => \nx.n10641\
        );

    \I__6361\ : InMux
    port map (
            O => \N__32820\,
            I => \N__32816\
        );

    \I__6360\ : InMux
    port map (
            O => \N__32819\,
            I => \N__32813\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__32816\,
            I => \N__32807\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__32813\,
            I => \N__32807\
        );

    \I__6357\ : InMux
    port map (
            O => \N__32812\,
            I => \N__32804\
        );

    \I__6356\ : Span4Mux_h
    port map (
            O => \N__32807\,
            I => \N__32801\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__32804\,
            I => \N__32798\
        );

    \I__6354\ : Odrv4
    port map (
            O => \N__32801\,
            I => \nx.n1895\
        );

    \I__6353\ : Odrv12
    port map (
            O => \N__32798\,
            I => \nx.n1895\
        );

    \I__6352\ : InMux
    port map (
            O => \N__32793\,
            I => \N__32788\
        );

    \I__6351\ : InMux
    port map (
            O => \N__32792\,
            I => \N__32785\
        );

    \I__6350\ : CascadeMux
    port map (
            O => \N__32791\,
            I => \N__32782\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__32788\,
            I => \N__32777\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__32785\,
            I => \N__32777\
        );

    \I__6347\ : InMux
    port map (
            O => \N__32782\,
            I => \N__32774\
        );

    \I__6346\ : Odrv4
    port map (
            O => \N__32777\,
            I => \nx.n1896\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__32774\,
            I => \nx.n1896\
        );

    \I__6344\ : InMux
    port map (
            O => \N__32769\,
            I => \N__32766\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__32766\,
            I => \N__32760\
        );

    \I__6342\ : InMux
    port map (
            O => \N__32765\,
            I => \N__32757\
        );

    \I__6341\ : InMux
    port map (
            O => \N__32764\,
            I => \N__32754\
        );

    \I__6340\ : InMux
    port map (
            O => \N__32763\,
            I => \N__32751\
        );

    \I__6339\ : Span4Mux_h
    port map (
            O => \N__32760\,
            I => \N__32746\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__32757\,
            I => \N__32746\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__32754\,
            I => \N__32740\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__32751\,
            I => \N__32740\
        );

    \I__6335\ : Span4Mux_h
    port map (
            O => \N__32746\,
            I => \N__32737\
        );

    \I__6334\ : InMux
    port map (
            O => \N__32745\,
            I => \N__32734\
        );

    \I__6333\ : Span4Mux_h
    port map (
            O => \N__32740\,
            I => \N__32731\
        );

    \I__6332\ : Span4Mux_h
    port map (
            O => \N__32737\,
            I => \N__32728\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__32734\,
            I => \nx.bit_ctr_17\
        );

    \I__6330\ : Odrv4
    port map (
            O => \N__32731\,
            I => \nx.bit_ctr_17\
        );

    \I__6329\ : Odrv4
    port map (
            O => \N__32728\,
            I => \nx.bit_ctr_17\
        );

    \I__6328\ : InMux
    port map (
            O => \N__32721\,
            I => \N__32718\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__32718\,
            I => \N__32714\
        );

    \I__6326\ : InMux
    port map (
            O => \N__32717\,
            I => \N__32711\
        );

    \I__6325\ : Span4Mux_h
    port map (
            O => \N__32714\,
            I => \N__32705\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__32711\,
            I => \N__32702\
        );

    \I__6323\ : InMux
    port map (
            O => \N__32710\,
            I => \N__32699\
        );

    \I__6322\ : InMux
    port map (
            O => \N__32709\,
            I => \N__32694\
        );

    \I__6321\ : InMux
    port map (
            O => \N__32708\,
            I => \N__32694\
        );

    \I__6320\ : Span4Mux_h
    port map (
            O => \N__32705\,
            I => \N__32689\
        );

    \I__6319\ : Span4Mux_s3_h
    port map (
            O => \N__32702\,
            I => \N__32689\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__32699\,
            I => \nx.bit_ctr_22\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__32694\,
            I => \nx.bit_ctr_22\
        );

    \I__6316\ : Odrv4
    port map (
            O => \N__32689\,
            I => \nx.bit_ctr_22\
        );

    \I__6315\ : InMux
    port map (
            O => \N__32682\,
            I => \N__32679\
        );

    \I__6314\ : LocalMux
    port map (
            O => \N__32679\,
            I => \N__32676\
        );

    \I__6313\ : Span4Mux_h
    port map (
            O => \N__32676\,
            I => \N__32673\
        );

    \I__6312\ : Span4Mux_h
    port map (
            O => \N__32673\,
            I => \N__32670\
        );

    \I__6311\ : Odrv4
    port map (
            O => \N__32670\,
            I => \nx.n30_adj_703\
        );

    \I__6310\ : CascadeMux
    port map (
            O => \N__32667\,
            I => \N__32663\
        );

    \I__6309\ : InMux
    port map (
            O => \N__32666\,
            I => \N__32659\
        );

    \I__6308\ : InMux
    port map (
            O => \N__32663\,
            I => \N__32656\
        );

    \I__6307\ : InMux
    port map (
            O => \N__32662\,
            I => \N__32653\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__32659\,
            I => \N__32648\
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__32656\,
            I => \N__32648\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__32653\,
            I => \nx.n1809\
        );

    \I__6303\ : Odrv4
    port map (
            O => \N__32648\,
            I => \nx.n1809\
        );

    \I__6302\ : InMux
    port map (
            O => \N__32643\,
            I => \N__32640\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__32640\,
            I => \N__32637\
        );

    \I__6300\ : Span4Mux_v
    port map (
            O => \N__32637\,
            I => \N__32634\
        );

    \I__6299\ : Odrv4
    port map (
            O => \N__32634\,
            I => \nx.n1876\
        );

    \I__6298\ : InMux
    port map (
            O => \N__32631\,
            I => \nx.n10628\
        );

    \I__6297\ : CascadeMux
    port map (
            O => \N__32628\,
            I => \N__32625\
        );

    \I__6296\ : InMux
    port map (
            O => \N__32625\,
            I => \N__32620\
        );

    \I__6295\ : InMux
    port map (
            O => \N__32624\,
            I => \N__32615\
        );

    \I__6294\ : InMux
    port map (
            O => \N__32623\,
            I => \N__32615\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__32620\,
            I => \N__32612\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__32615\,
            I => \nx.n1808\
        );

    \I__6291\ : Odrv12
    port map (
            O => \N__32612\,
            I => \nx.n1808\
        );

    \I__6290\ : InMux
    port map (
            O => \N__32607\,
            I => \N__32604\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__32604\,
            I => \N__32601\
        );

    \I__6288\ : Span4Mux_h
    port map (
            O => \N__32601\,
            I => \N__32598\
        );

    \I__6287\ : Odrv4
    port map (
            O => \N__32598\,
            I => \nx.n1875\
        );

    \I__6286\ : InMux
    port map (
            O => \N__32595\,
            I => \nx.n10629\
        );

    \I__6285\ : CascadeMux
    port map (
            O => \N__32592\,
            I => \N__32589\
        );

    \I__6284\ : InMux
    port map (
            O => \N__32589\,
            I => \N__32582\
        );

    \I__6283\ : InMux
    port map (
            O => \N__32588\,
            I => \N__32582\
        );

    \I__6282\ : CascadeMux
    port map (
            O => \N__32587\,
            I => \N__32579\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__32582\,
            I => \N__32576\
        );

    \I__6280\ : InMux
    port map (
            O => \N__32579\,
            I => \N__32573\
        );

    \I__6279\ : Odrv4
    port map (
            O => \N__32576\,
            I => \nx.n1807\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__32573\,
            I => \nx.n1807\
        );

    \I__6277\ : InMux
    port map (
            O => \N__32568\,
            I => \N__32565\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__32565\,
            I => \N__32562\
        );

    \I__6275\ : Span4Mux_h
    port map (
            O => \N__32562\,
            I => \N__32559\
        );

    \I__6274\ : Odrv4
    port map (
            O => \N__32559\,
            I => \nx.n1874\
        );

    \I__6273\ : InMux
    port map (
            O => \N__32556\,
            I => \nx.n10630\
        );

    \I__6272\ : CascadeMux
    port map (
            O => \N__32553\,
            I => \N__32550\
        );

    \I__6271\ : InMux
    port map (
            O => \N__32550\,
            I => \N__32547\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__32547\,
            I => \N__32544\
        );

    \I__6269\ : Odrv4
    port map (
            O => \N__32544\,
            I => \nx.n1873\
        );

    \I__6268\ : InMux
    port map (
            O => \N__32541\,
            I => \nx.n10631\
        );

    \I__6267\ : InMux
    port map (
            O => \N__32538\,
            I => \N__32534\
        );

    \I__6266\ : CascadeMux
    port map (
            O => \N__32537\,
            I => \N__32531\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__32534\,
            I => \N__32527\
        );

    \I__6264\ : InMux
    port map (
            O => \N__32531\,
            I => \N__32524\
        );

    \I__6263\ : InMux
    port map (
            O => \N__32530\,
            I => \N__32521\
        );

    \I__6262\ : Span4Mux_v
    port map (
            O => \N__32527\,
            I => \N__32516\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__32524\,
            I => \N__32516\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__32521\,
            I => \nx.n1805\
        );

    \I__6259\ : Odrv4
    port map (
            O => \N__32516\,
            I => \nx.n1805\
        );

    \I__6258\ : CascadeMux
    port map (
            O => \N__32511\,
            I => \N__32508\
        );

    \I__6257\ : InMux
    port map (
            O => \N__32508\,
            I => \N__32505\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__32505\,
            I => \N__32502\
        );

    \I__6255\ : Span4Mux_v
    port map (
            O => \N__32502\,
            I => \N__32499\
        );

    \I__6254\ : Span4Mux_h
    port map (
            O => \N__32499\,
            I => \N__32496\
        );

    \I__6253\ : Odrv4
    port map (
            O => \N__32496\,
            I => \nx.n1872\
        );

    \I__6252\ : InMux
    port map (
            O => \N__32493\,
            I => \nx.n10632\
        );

    \I__6251\ : CascadeMux
    port map (
            O => \N__32490\,
            I => \N__32487\
        );

    \I__6250\ : InMux
    port map (
            O => \N__32487\,
            I => \N__32483\
        );

    \I__6249\ : InMux
    port map (
            O => \N__32486\,
            I => \N__32480\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__32483\,
            I => \N__32477\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__32480\,
            I => \nx.n1804\
        );

    \I__6246\ : Odrv4
    port map (
            O => \N__32477\,
            I => \nx.n1804\
        );

    \I__6245\ : InMux
    port map (
            O => \N__32472\,
            I => \N__32469\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__32469\,
            I => \N__32466\
        );

    \I__6243\ : Span4Mux_h
    port map (
            O => \N__32466\,
            I => \N__32463\
        );

    \I__6242\ : Odrv4
    port map (
            O => \N__32463\,
            I => \nx.n1871\
        );

    \I__6241\ : InMux
    port map (
            O => \N__32460\,
            I => \nx.n10633\
        );

    \I__6240\ : InMux
    port map (
            O => \N__32457\,
            I => \N__32453\
        );

    \I__6239\ : InMux
    port map (
            O => \N__32456\,
            I => \N__32450\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__32453\,
            I => \N__32444\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__32450\,
            I => \N__32444\
        );

    \I__6236\ : InMux
    port map (
            O => \N__32449\,
            I => \N__32441\
        );

    \I__6235\ : Span4Mux_h
    port map (
            O => \N__32444\,
            I => \N__32438\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__32441\,
            I => \N__32435\
        );

    \I__6233\ : Odrv4
    port map (
            O => \N__32438\,
            I => \nx.n1901\
        );

    \I__6232\ : Odrv4
    port map (
            O => \N__32435\,
            I => \nx.n1901\
        );

    \I__6231\ : InMux
    port map (
            O => \N__32430\,
            I => \N__32426\
        );

    \I__6230\ : InMux
    port map (
            O => \N__32429\,
            I => \N__32423\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__32426\,
            I => \N__32417\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__32423\,
            I => \N__32417\
        );

    \I__6227\ : InMux
    port map (
            O => \N__32422\,
            I => \N__32414\
        );

    \I__6226\ : Odrv4
    port map (
            O => \N__32417\,
            I => \nx.n1905\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__32414\,
            I => \nx.n1905\
        );

    \I__6224\ : InMux
    port map (
            O => \N__32409\,
            I => \N__32406\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__32406\,
            I => \N__32403\
        );

    \I__6222\ : Odrv4
    port map (
            O => \N__32403\,
            I => \nx.n25_adj_606\
        );

    \I__6221\ : CascadeMux
    port map (
            O => \N__32400\,
            I => \N__32397\
        );

    \I__6220\ : InMux
    port map (
            O => \N__32397\,
            I => \N__32394\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__32394\,
            I => \N__32391\
        );

    \I__6218\ : Odrv12
    port map (
            O => \N__32391\,
            I => \nx.n22\
        );

    \I__6217\ : InMux
    port map (
            O => \N__32388\,
            I => \N__32384\
        );

    \I__6216\ : InMux
    port map (
            O => \N__32387\,
            I => \N__32381\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__32384\,
            I => \N__32375\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__32381\,
            I => \N__32375\
        );

    \I__6213\ : InMux
    port map (
            O => \N__32380\,
            I => \N__32372\
        );

    \I__6212\ : Odrv4
    port map (
            O => \N__32375\,
            I => \nx.n1900\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__32372\,
            I => \nx.n1900\
        );

    \I__6210\ : CascadeMux
    port map (
            O => \N__32367\,
            I => \nx.n1799_cascade_\
        );

    \I__6209\ : InMux
    port map (
            O => \N__32364\,
            I => \N__32360\
        );

    \I__6208\ : InMux
    port map (
            O => \N__32363\,
            I => \N__32357\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__32360\,
            I => \N__32351\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__32357\,
            I => \N__32351\
        );

    \I__6205\ : InMux
    port map (
            O => \N__32356\,
            I => \N__32348\
        );

    \I__6204\ : Span4Mux_h
    port map (
            O => \N__32351\,
            I => \N__32345\
        );

    \I__6203\ : LocalMux
    port map (
            O => \N__32348\,
            I => \N__32342\
        );

    \I__6202\ : Odrv4
    port map (
            O => \N__32345\,
            I => \nx.n1898\
        );

    \I__6201\ : Odrv12
    port map (
            O => \N__32342\,
            I => \nx.n1898\
        );

    \I__6200\ : CascadeMux
    port map (
            O => \N__32337\,
            I => \nx.n1797_cascade_\
        );

    \I__6199\ : CascadeMux
    port map (
            O => \N__32334\,
            I => \N__32329\
        );

    \I__6198\ : InMux
    port map (
            O => \N__32333\,
            I => \N__32324\
        );

    \I__6197\ : InMux
    port map (
            O => \N__32332\,
            I => \N__32324\
        );

    \I__6196\ : InMux
    port map (
            O => \N__32329\,
            I => \N__32321\
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__32324\,
            I => \N__32318\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__32321\,
            I => \N__32315\
        );

    \I__6193\ : Span4Mux_h
    port map (
            O => \N__32318\,
            I => \N__32312\
        );

    \I__6192\ : Span4Mux_h
    port map (
            O => \N__32315\,
            I => \N__32309\
        );

    \I__6191\ : Odrv4
    port map (
            O => \N__32312\,
            I => \nx.n2001\
        );

    \I__6190\ : Odrv4
    port map (
            O => \N__32309\,
            I => \nx.n2001\
        );

    \I__6189\ : InMux
    port map (
            O => \N__32304\,
            I => \N__32301\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__32301\,
            I => \N__32298\
        );

    \I__6187\ : Odrv4
    port map (
            O => \N__32298\,
            I => \nx.n2068\
        );

    \I__6186\ : InMux
    port map (
            O => \N__32295\,
            I => \nx.n10665\
        );

    \I__6185\ : CascadeMux
    port map (
            O => \N__32292\,
            I => \N__32288\
        );

    \I__6184\ : CascadeMux
    port map (
            O => \N__32291\,
            I => \N__32284\
        );

    \I__6183\ : InMux
    port map (
            O => \N__32288\,
            I => \N__32279\
        );

    \I__6182\ : InMux
    port map (
            O => \N__32287\,
            I => \N__32279\
        );

    \I__6181\ : InMux
    port map (
            O => \N__32284\,
            I => \N__32276\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__32279\,
            I => \N__32273\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__32276\,
            I => \N__32270\
        );

    \I__6178\ : Span4Mux_h
    port map (
            O => \N__32273\,
            I => \N__32267\
        );

    \I__6177\ : Span4Mux_h
    port map (
            O => \N__32270\,
            I => \N__32264\
        );

    \I__6176\ : Odrv4
    port map (
            O => \N__32267\,
            I => \nx.n2000\
        );

    \I__6175\ : Odrv4
    port map (
            O => \N__32264\,
            I => \nx.n2000\
        );

    \I__6174\ : InMux
    port map (
            O => \N__32259\,
            I => \N__32256\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__32256\,
            I => \N__32253\
        );

    \I__6172\ : Odrv4
    port map (
            O => \N__32253\,
            I => \nx.n2067\
        );

    \I__6171\ : InMux
    port map (
            O => \N__32250\,
            I => \nx.n10666\
        );

    \I__6170\ : CascadeMux
    port map (
            O => \N__32247\,
            I => \N__32242\
        );

    \I__6169\ : CascadeMux
    port map (
            O => \N__32246\,
            I => \N__32239\
        );

    \I__6168\ : InMux
    port map (
            O => \N__32245\,
            I => \N__32234\
        );

    \I__6167\ : InMux
    port map (
            O => \N__32242\,
            I => \N__32234\
        );

    \I__6166\ : InMux
    port map (
            O => \N__32239\,
            I => \N__32231\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__32234\,
            I => \N__32228\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__32231\,
            I => \N__32225\
        );

    \I__6163\ : Span4Mux_h
    port map (
            O => \N__32228\,
            I => \N__32222\
        );

    \I__6162\ : Span4Mux_v
    port map (
            O => \N__32225\,
            I => \N__32219\
        );

    \I__6161\ : Odrv4
    port map (
            O => \N__32222\,
            I => \nx.n1999\
        );

    \I__6160\ : Odrv4
    port map (
            O => \N__32219\,
            I => \nx.n1999\
        );

    \I__6159\ : InMux
    port map (
            O => \N__32214\,
            I => \N__32211\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__32211\,
            I => \N__32208\
        );

    \I__6157\ : Odrv4
    port map (
            O => \N__32208\,
            I => \nx.n2066\
        );

    \I__6156\ : InMux
    port map (
            O => \N__32205\,
            I => \nx.n10667\
        );

    \I__6155\ : InMux
    port map (
            O => \N__32202\,
            I => \nx.n10668\
        );

    \I__6154\ : InMux
    port map (
            O => \N__32199\,
            I => \nx.n10669\
        );

    \I__6153\ : InMux
    port map (
            O => \N__32196\,
            I => \N__32192\
        );

    \I__6152\ : CascadeMux
    port map (
            O => \N__32195\,
            I => \N__32189\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__32192\,
            I => \N__32186\
        );

    \I__6150\ : InMux
    port map (
            O => \N__32189\,
            I => \N__32183\
        );

    \I__6149\ : Span4Mux_h
    port map (
            O => \N__32186\,
            I => \N__32179\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__32183\,
            I => \N__32176\
        );

    \I__6147\ : InMux
    port map (
            O => \N__32182\,
            I => \N__32173\
        );

    \I__6146\ : Span4Mux_v
    port map (
            O => \N__32179\,
            I => \N__32170\
        );

    \I__6145\ : Span4Mux_h
    port map (
            O => \N__32176\,
            I => \N__32167\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__32173\,
            I => \N__32164\
        );

    \I__6143\ : Odrv4
    port map (
            O => \N__32170\,
            I => \nx.n1996\
        );

    \I__6142\ : Odrv4
    port map (
            O => \N__32167\,
            I => \nx.n1996\
        );

    \I__6141\ : Odrv12
    port map (
            O => \N__32164\,
            I => \nx.n1996\
        );

    \I__6140\ : CascadeMux
    port map (
            O => \N__32157\,
            I => \N__32154\
        );

    \I__6139\ : InMux
    port map (
            O => \N__32154\,
            I => \N__32151\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__32151\,
            I => \N__32148\
        );

    \I__6137\ : Span4Mux_h
    port map (
            O => \N__32148\,
            I => \N__32145\
        );

    \I__6136\ : Odrv4
    port map (
            O => \N__32145\,
            I => \nx.n2063\
        );

    \I__6135\ : InMux
    port map (
            O => \N__32142\,
            I => \nx.n10670\
        );

    \I__6134\ : InMux
    port map (
            O => \N__32139\,
            I => \nx.n10671\
        );

    \I__6133\ : CascadeMux
    port map (
            O => \N__32136\,
            I => \N__32133\
        );

    \I__6132\ : InMux
    port map (
            O => \N__32133\,
            I => \N__32130\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__32130\,
            I => \N__32126\
        );

    \I__6130\ : InMux
    port map (
            O => \N__32129\,
            I => \N__32123\
        );

    \I__6129\ : Span4Mux_h
    port map (
            O => \N__32126\,
            I => \N__32120\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__32123\,
            I => \N__32117\
        );

    \I__6127\ : Odrv4
    port map (
            O => \N__32120\,
            I => \nx.n1994\
        );

    \I__6126\ : Odrv12
    port map (
            O => \N__32117\,
            I => \nx.n1994\
        );

    \I__6125\ : InMux
    port map (
            O => \N__32112\,
            I => \bfn_9_25_0_\
        );

    \I__6124\ : InMux
    port map (
            O => \N__32109\,
            I => \bfn_9_23_0_\
        );

    \I__6123\ : InMux
    port map (
            O => \N__32106\,
            I => \nx.n10657\
        );

    \I__6122\ : InMux
    port map (
            O => \N__32103\,
            I => \nx.n10658\
        );

    \I__6121\ : InMux
    port map (
            O => \N__32100\,
            I => \nx.n10659\
        );

    \I__6120\ : InMux
    port map (
            O => \N__32097\,
            I => \N__32093\
        );

    \I__6119\ : CascadeMux
    port map (
            O => \N__32096\,
            I => \N__32090\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__32093\,
            I => \N__32086\
        );

    \I__6117\ : InMux
    port map (
            O => \N__32090\,
            I => \N__32083\
        );

    \I__6116\ : CascadeMux
    port map (
            O => \N__32089\,
            I => \N__32080\
        );

    \I__6115\ : Span4Mux_h
    port map (
            O => \N__32086\,
            I => \N__32077\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__32083\,
            I => \N__32074\
        );

    \I__6113\ : InMux
    port map (
            O => \N__32080\,
            I => \N__32071\
        );

    \I__6112\ : Span4Mux_v
    port map (
            O => \N__32077\,
            I => \N__32066\
        );

    \I__6111\ : Span4Mux_v
    port map (
            O => \N__32074\,
            I => \N__32066\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__32071\,
            I => \nx.n2006\
        );

    \I__6109\ : Odrv4
    port map (
            O => \N__32066\,
            I => \nx.n2006\
        );

    \I__6108\ : InMux
    port map (
            O => \N__32061\,
            I => \N__32058\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__32058\,
            I => \N__32055\
        );

    \I__6106\ : Odrv12
    port map (
            O => \N__32055\,
            I => \nx.n2073\
        );

    \I__6105\ : InMux
    port map (
            O => \N__32052\,
            I => \nx.n10660\
        );

    \I__6104\ : CascadeMux
    port map (
            O => \N__32049\,
            I => \N__32045\
        );

    \I__6103\ : CascadeMux
    port map (
            O => \N__32048\,
            I => \N__32042\
        );

    \I__6102\ : InMux
    port map (
            O => \N__32045\,
            I => \N__32039\
        );

    \I__6101\ : InMux
    port map (
            O => \N__32042\,
            I => \N__32036\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__32039\,
            I => \N__32033\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__32036\,
            I => \N__32029\
        );

    \I__6098\ : Span4Mux_h
    port map (
            O => \N__32033\,
            I => \N__32026\
        );

    \I__6097\ : InMux
    port map (
            O => \N__32032\,
            I => \N__32023\
        );

    \I__6096\ : Span4Mux_h
    port map (
            O => \N__32029\,
            I => \N__32020\
        );

    \I__6095\ : Odrv4
    port map (
            O => \N__32026\,
            I => \nx.n2005\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__32023\,
            I => \nx.n2005\
        );

    \I__6093\ : Odrv4
    port map (
            O => \N__32020\,
            I => \nx.n2005\
        );

    \I__6092\ : InMux
    port map (
            O => \N__32013\,
            I => \N__32010\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__32010\,
            I => \N__32007\
        );

    \I__6090\ : Odrv4
    port map (
            O => \N__32007\,
            I => \nx.n2072\
        );

    \I__6089\ : InMux
    port map (
            O => \N__32004\,
            I => \nx.n10661\
        );

    \I__6088\ : CascadeMux
    port map (
            O => \N__32001\,
            I => \N__31997\
        );

    \I__6087\ : CascadeMux
    port map (
            O => \N__32000\,
            I => \N__31994\
        );

    \I__6086\ : InMux
    port map (
            O => \N__31997\,
            I => \N__31991\
        );

    \I__6085\ : InMux
    port map (
            O => \N__31994\,
            I => \N__31988\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__31991\,
            I => \N__31985\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__31988\,
            I => \N__31981\
        );

    \I__6082\ : Span4Mux_v
    port map (
            O => \N__31985\,
            I => \N__31978\
        );

    \I__6081\ : InMux
    port map (
            O => \N__31984\,
            I => \N__31975\
        );

    \I__6080\ : Span4Mux_h
    port map (
            O => \N__31981\,
            I => \N__31972\
        );

    \I__6079\ : Odrv4
    port map (
            O => \N__31978\,
            I => \nx.n2004\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__31975\,
            I => \nx.n2004\
        );

    \I__6077\ : Odrv4
    port map (
            O => \N__31972\,
            I => \nx.n2004\
        );

    \I__6076\ : InMux
    port map (
            O => \N__31965\,
            I => \N__31962\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__31962\,
            I => \nx.n2071\
        );

    \I__6074\ : InMux
    port map (
            O => \N__31959\,
            I => \nx.n10662\
        );

    \I__6073\ : InMux
    port map (
            O => \N__31956\,
            I => \nx.n10663\
        );

    \I__6072\ : InMux
    port map (
            O => \N__31953\,
            I => \bfn_9_24_0_\
        );

    \I__6071\ : CascadeMux
    port map (
            O => \N__31950\,
            I => \nx.n2595_cascade_\
        );

    \I__6070\ : InMux
    port map (
            O => \N__31947\,
            I => \N__31944\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__31944\,
            I => \N__31941\
        );

    \I__6068\ : Span4Mux_h
    port map (
            O => \N__31941\,
            I => \N__31938\
        );

    \I__6067\ : Odrv4
    port map (
            O => \N__31938\,
            I => \nx.n28_adj_663\
        );

    \I__6066\ : CascadeMux
    port map (
            O => \N__31935\,
            I => \nx.n26_adj_664_cascade_\
        );

    \I__6065\ : InMux
    port map (
            O => \N__31932\,
            I => \N__31929\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__31929\,
            I => \N__31926\
        );

    \I__6063\ : Odrv4
    port map (
            O => \N__31926\,
            I => \nx.n25_adj_666\
        );

    \I__6062\ : CascadeMux
    port map (
            O => \N__31923\,
            I => \nx.n2027_cascade_\
        );

    \I__6061\ : CascadeMux
    port map (
            O => \N__31920\,
            I => \nx.n2099_cascade_\
        );

    \I__6060\ : InMux
    port map (
            O => \N__31917\,
            I => \N__31914\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__31914\,
            I => \N__31910\
        );

    \I__6058\ : CascadeMux
    port map (
            O => \N__31913\,
            I => \N__31907\
        );

    \I__6057\ : Span4Mux_h
    port map (
            O => \N__31910\,
            I => \N__31903\
        );

    \I__6056\ : InMux
    port map (
            O => \N__31907\,
            I => \N__31900\
        );

    \I__6055\ : InMux
    port map (
            O => \N__31906\,
            I => \N__31897\
        );

    \I__6054\ : Odrv4
    port map (
            O => \N__31903\,
            I => \nx.n2904\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__31900\,
            I => \nx.n2904\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__31897\,
            I => \nx.n2904\
        );

    \I__6051\ : CascadeMux
    port map (
            O => \N__31890\,
            I => \N__31887\
        );

    \I__6050\ : InMux
    port map (
            O => \N__31887\,
            I => \N__31884\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__31884\,
            I => \N__31881\
        );

    \I__6048\ : Odrv12
    port map (
            O => \N__31881\,
            I => \nx.n2971\
        );

    \I__6047\ : InMux
    port map (
            O => \N__31878\,
            I => \N__31871\
        );

    \I__6046\ : CascadeMux
    port map (
            O => \N__31877\,
            I => \N__31868\
        );

    \I__6045\ : CascadeMux
    port map (
            O => \N__31876\,
            I => \N__31860\
        );

    \I__6044\ : CascadeMux
    port map (
            O => \N__31875\,
            I => \N__31855\
        );

    \I__6043\ : InMux
    port map (
            O => \N__31874\,
            I => \N__31848\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__31871\,
            I => \N__31845\
        );

    \I__6041\ : InMux
    port map (
            O => \N__31868\,
            I => \N__31840\
        );

    \I__6040\ : InMux
    port map (
            O => \N__31867\,
            I => \N__31840\
        );

    \I__6039\ : CascadeMux
    port map (
            O => \N__31866\,
            I => \N__31830\
        );

    \I__6038\ : CascadeMux
    port map (
            O => \N__31865\,
            I => \N__31827\
        );

    \I__6037\ : CascadeMux
    port map (
            O => \N__31864\,
            I => \N__31823\
        );

    \I__6036\ : CascadeMux
    port map (
            O => \N__31863\,
            I => \N__31819\
        );

    \I__6035\ : InMux
    port map (
            O => \N__31860\,
            I => \N__31814\
        );

    \I__6034\ : InMux
    port map (
            O => \N__31859\,
            I => \N__31814\
        );

    \I__6033\ : InMux
    port map (
            O => \N__31858\,
            I => \N__31807\
        );

    \I__6032\ : InMux
    port map (
            O => \N__31855\,
            I => \N__31807\
        );

    \I__6031\ : InMux
    port map (
            O => \N__31854\,
            I => \N__31807\
        );

    \I__6030\ : InMux
    port map (
            O => \N__31853\,
            I => \N__31800\
        );

    \I__6029\ : InMux
    port map (
            O => \N__31852\,
            I => \N__31800\
        );

    \I__6028\ : InMux
    port map (
            O => \N__31851\,
            I => \N__31800\
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__31848\,
            I => \N__31797\
        );

    \I__6026\ : Span4Mux_v
    port map (
            O => \N__31845\,
            I => \N__31794\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__31840\,
            I => \N__31791\
        );

    \I__6024\ : InMux
    port map (
            O => \N__31839\,
            I => \N__31784\
        );

    \I__6023\ : InMux
    port map (
            O => \N__31838\,
            I => \N__31784\
        );

    \I__6022\ : InMux
    port map (
            O => \N__31837\,
            I => \N__31784\
        );

    \I__6021\ : InMux
    port map (
            O => \N__31836\,
            I => \N__31775\
        );

    \I__6020\ : InMux
    port map (
            O => \N__31835\,
            I => \N__31775\
        );

    \I__6019\ : InMux
    port map (
            O => \N__31834\,
            I => \N__31775\
        );

    \I__6018\ : InMux
    port map (
            O => \N__31833\,
            I => \N__31775\
        );

    \I__6017\ : InMux
    port map (
            O => \N__31830\,
            I => \N__31762\
        );

    \I__6016\ : InMux
    port map (
            O => \N__31827\,
            I => \N__31762\
        );

    \I__6015\ : InMux
    port map (
            O => \N__31826\,
            I => \N__31762\
        );

    \I__6014\ : InMux
    port map (
            O => \N__31823\,
            I => \N__31762\
        );

    \I__6013\ : InMux
    port map (
            O => \N__31822\,
            I => \N__31762\
        );

    \I__6012\ : InMux
    port map (
            O => \N__31819\,
            I => \N__31762\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__31814\,
            I => \N__31759\
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__31807\,
            I => \N__31756\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__31800\,
            I => \N__31749\
        );

    \I__6008\ : Span4Mux_s1_h
    port map (
            O => \N__31797\,
            I => \N__31749\
        );

    \I__6007\ : Span4Mux_h
    port map (
            O => \N__31794\,
            I => \N__31749\
        );

    \I__6006\ : Odrv4
    port map (
            O => \N__31791\,
            I => \nx.n2918\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__31784\,
            I => \nx.n2918\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__31775\,
            I => \nx.n2918\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__31762\,
            I => \nx.n2918\
        );

    \I__6002\ : Odrv4
    port map (
            O => \N__31759\,
            I => \nx.n2918\
        );

    \I__6001\ : Odrv4
    port map (
            O => \N__31756\,
            I => \nx.n2918\
        );

    \I__6000\ : Odrv4
    port map (
            O => \N__31749\,
            I => \nx.n2918\
        );

    \I__5999\ : CascadeMux
    port map (
            O => \N__31734\,
            I => \N__31729\
        );

    \I__5998\ : InMux
    port map (
            O => \N__31733\,
            I => \N__31726\
        );

    \I__5997\ : InMux
    port map (
            O => \N__31732\,
            I => \N__31723\
        );

    \I__5996\ : InMux
    port map (
            O => \N__31729\,
            I => \N__31720\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__31726\,
            I => \N__31717\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__31723\,
            I => \N__31714\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__31720\,
            I => \N__31711\
        );

    \I__5992\ : Span4Mux_h
    port map (
            O => \N__31717\,
            I => \N__31708\
        );

    \I__5991\ : Span4Mux_v
    port map (
            O => \N__31714\,
            I => \N__31703\
        );

    \I__5990\ : Span4Mux_v
    port map (
            O => \N__31711\,
            I => \N__31703\
        );

    \I__5989\ : Span4Mux_h
    port map (
            O => \N__31708\,
            I => \N__31700\
        );

    \I__5988\ : Span4Mux_h
    port map (
            O => \N__31703\,
            I => \N__31697\
        );

    \I__5987\ : Odrv4
    port map (
            O => \N__31700\,
            I => \nx.n3003\
        );

    \I__5986\ : Odrv4
    port map (
            O => \N__31697\,
            I => \nx.n3003\
        );

    \I__5985\ : CascadeMux
    port map (
            O => \N__31692\,
            I => \N__31689\
        );

    \I__5984\ : InMux
    port map (
            O => \N__31689\,
            I => \N__31685\
        );

    \I__5983\ : InMux
    port map (
            O => \N__31688\,
            I => \N__31682\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__31685\,
            I => \N__31679\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__31682\,
            I => \N__31676\
        );

    \I__5980\ : Span4Mux_v
    port map (
            O => \N__31679\,
            I => \N__31673\
        );

    \I__5979\ : Odrv4
    port map (
            O => \N__31676\,
            I => \nx.n2689\
        );

    \I__5978\ : Odrv4
    port map (
            O => \N__31673\,
            I => \nx.n2689\
        );

    \I__5977\ : CascadeMux
    port map (
            O => \N__31668\,
            I => \N__31664\
        );

    \I__5976\ : CascadeMux
    port map (
            O => \N__31667\,
            I => \N__31661\
        );

    \I__5975\ : InMux
    port map (
            O => \N__31664\,
            I => \N__31658\
        );

    \I__5974\ : InMux
    port map (
            O => \N__31661\,
            I => \N__31655\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__31658\,
            I => \N__31652\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__31655\,
            I => \N__31649\
        );

    \I__5971\ : Span4Mux_v
    port map (
            O => \N__31652\,
            I => \N__31645\
        );

    \I__5970\ : Span4Mux_h
    port map (
            O => \N__31649\,
            I => \N__31642\
        );

    \I__5969\ : InMux
    port map (
            O => \N__31648\,
            I => \N__31639\
        );

    \I__5968\ : Odrv4
    port map (
            O => \N__31645\,
            I => \nx.n2690\
        );

    \I__5967\ : Odrv4
    port map (
            O => \N__31642\,
            I => \nx.n2690\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__31639\,
            I => \nx.n2690\
        );

    \I__5965\ : CascadeMux
    port map (
            O => \N__31632\,
            I => \nx.n2689_cascade_\
        );

    \I__5964\ : CascadeMux
    port map (
            O => \N__31629\,
            I => \N__31625\
        );

    \I__5963\ : CascadeMux
    port map (
            O => \N__31628\,
            I => \N__31622\
        );

    \I__5962\ : InMux
    port map (
            O => \N__31625\,
            I => \N__31619\
        );

    \I__5961\ : InMux
    port map (
            O => \N__31622\,
            I => \N__31616\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__31619\,
            I => \N__31611\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__31616\,
            I => \N__31611\
        );

    \I__5958\ : Span4Mux_v
    port map (
            O => \N__31611\,
            I => \N__31607\
        );

    \I__5957\ : InMux
    port map (
            O => \N__31610\,
            I => \N__31604\
        );

    \I__5956\ : Odrv4
    port map (
            O => \N__31607\,
            I => \nx.n2691\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__31604\,
            I => \nx.n2691\
        );

    \I__5954\ : InMux
    port map (
            O => \N__31599\,
            I => \N__31595\
        );

    \I__5953\ : CascadeMux
    port map (
            O => \N__31598\,
            I => \N__31592\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__31595\,
            I => \N__31589\
        );

    \I__5951\ : InMux
    port map (
            O => \N__31592\,
            I => \N__31586\
        );

    \I__5950\ : Span4Mux_h
    port map (
            O => \N__31589\,
            I => \N__31580\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__31586\,
            I => \N__31580\
        );

    \I__5948\ : InMux
    port map (
            O => \N__31585\,
            I => \N__31577\
        );

    \I__5947\ : Odrv4
    port map (
            O => \N__31580\,
            I => \nx.n2701\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__31577\,
            I => \nx.n2701\
        );

    \I__5945\ : CascadeMux
    port map (
            O => \N__31572\,
            I => \nx.n2105_cascade_\
        );

    \I__5944\ : InMux
    port map (
            O => \N__31569\,
            I => \N__31565\
        );

    \I__5943\ : CascadeMux
    port map (
            O => \N__31568\,
            I => \N__31561\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__31565\,
            I => \N__31558\
        );

    \I__5941\ : InMux
    port map (
            O => \N__31564\,
            I => \N__31555\
        );

    \I__5940\ : InMux
    port map (
            O => \N__31561\,
            I => \N__31552\
        );

    \I__5939\ : Span4Mux_v
    port map (
            O => \N__31558\,
            I => \N__31545\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__31555\,
            I => \N__31545\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__31552\,
            I => \N__31545\
        );

    \I__5936\ : Odrv4
    port map (
            O => \N__31545\,
            I => \nx.n2704\
        );

    \I__5935\ : CascadeMux
    port map (
            O => \N__31542\,
            I => \N__31539\
        );

    \I__5934\ : InMux
    port map (
            O => \N__31539\,
            I => \N__31534\
        );

    \I__5933\ : InMux
    port map (
            O => \N__31538\,
            I => \N__31529\
        );

    \I__5932\ : InMux
    port map (
            O => \N__31537\,
            I => \N__31529\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__31534\,
            I => \N__31526\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__31529\,
            I => \N__31523\
        );

    \I__5929\ : Span4Mux_v
    port map (
            O => \N__31526\,
            I => \N__31518\
        );

    \I__5928\ : Span4Mux_h
    port map (
            O => \N__31523\,
            I => \N__31518\
        );

    \I__5927\ : Odrv4
    port map (
            O => \N__31518\,
            I => \nx.n2695\
        );

    \I__5926\ : CascadeMux
    port map (
            O => \N__31515\,
            I => \N__31512\
        );

    \I__5925\ : InMux
    port map (
            O => \N__31512\,
            I => \N__31508\
        );

    \I__5924\ : InMux
    port map (
            O => \N__31511\,
            I => \N__31505\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__31508\,
            I => \N__31500\
        );

    \I__5922\ : LocalMux
    port map (
            O => \N__31505\,
            I => \N__31500\
        );

    \I__5921\ : Span4Mux_v
    port map (
            O => \N__31500\,
            I => \N__31497\
        );

    \I__5920\ : Odrv4
    port map (
            O => \N__31497\,
            I => \nx.n2698\
        );

    \I__5919\ : CascadeMux
    port map (
            O => \N__31494\,
            I => \nx.n2698_cascade_\
        );

    \I__5918\ : InMux
    port map (
            O => \N__31491\,
            I => \N__31488\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__31488\,
            I => \N__31485\
        );

    \I__5916\ : Odrv4
    port map (
            O => \N__31485\,
            I => \nx.n39_adj_610\
        );

    \I__5915\ : InMux
    port map (
            O => \N__31482\,
            I => \N__31478\
        );

    \I__5914\ : CascadeMux
    port map (
            O => \N__31481\,
            I => \N__31475\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__31478\,
            I => \N__31471\
        );

    \I__5912\ : InMux
    port map (
            O => \N__31475\,
            I => \N__31468\
        );

    \I__5911\ : InMux
    port map (
            O => \N__31474\,
            I => \N__31465\
        );

    \I__5910\ : Span4Mux_h
    port map (
            O => \N__31471\,
            I => \N__31460\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__31468\,
            I => \N__31460\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__31465\,
            I => \nx.n2703\
        );

    \I__5907\ : Odrv4
    port map (
            O => \N__31460\,
            I => \nx.n2703\
        );

    \I__5906\ : InMux
    port map (
            O => \N__31455\,
            I => \N__31450\
        );

    \I__5905\ : InMux
    port map (
            O => \N__31454\,
            I => \N__31447\
        );

    \I__5904\ : CascadeMux
    port map (
            O => \N__31453\,
            I => \N__31444\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__31450\,
            I => \N__31441\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__31447\,
            I => \N__31438\
        );

    \I__5901\ : InMux
    port map (
            O => \N__31444\,
            I => \N__31435\
        );

    \I__5900\ : Span4Mux_v
    port map (
            O => \N__31441\,
            I => \N__31428\
        );

    \I__5899\ : Span4Mux_h
    port map (
            O => \N__31438\,
            I => \N__31428\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__31435\,
            I => \N__31428\
        );

    \I__5897\ : Odrv4
    port map (
            O => \N__31428\,
            I => \nx.n2709\
        );

    \I__5896\ : CascadeMux
    port map (
            O => \N__31425\,
            I => \nx.n2592_cascade_\
        );

    \I__5895\ : InMux
    port map (
            O => \N__31422\,
            I => \N__31419\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__31419\,
            I => \N__31416\
        );

    \I__5893\ : Span4Mux_h
    port map (
            O => \N__31416\,
            I => \N__31413\
        );

    \I__5892\ : Odrv4
    port map (
            O => \N__31413\,
            I => n13146
        );

    \I__5891\ : CascadeMux
    port map (
            O => \N__31410\,
            I => \n13462_cascade_\
        );

    \I__5890\ : InMux
    port map (
            O => \N__31407\,
            I => \N__31404\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__31404\,
            I => n13153
        );

    \I__5888\ : IoInMux
    port map (
            O => \N__31401\,
            I => \N__31398\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__31398\,
            I => \N__31395\
        );

    \I__5886\ : IoSpan4Mux
    port map (
            O => \N__31395\,
            I => \N__31392\
        );

    \I__5885\ : Span4Mux_s3_h
    port map (
            O => \N__31392\,
            I => \N__31389\
        );

    \I__5884\ : Span4Mux_h
    port map (
            O => \N__31389\,
            I => \N__31384\
        );

    \I__5883\ : InMux
    port map (
            O => \N__31388\,
            I => \N__31379\
        );

    \I__5882\ : InMux
    port map (
            O => \N__31387\,
            I => \N__31379\
        );

    \I__5881\ : Odrv4
    port map (
            O => \N__31384\,
            I => pin_out_3
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__31379\,
            I => pin_out_3
        );

    \I__5879\ : IoInMux
    port map (
            O => \N__31374\,
            I => \N__31371\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__31371\,
            I => \N__31368\
        );

    \I__5877\ : IoSpan4Mux
    port map (
            O => \N__31368\,
            I => \N__31365\
        );

    \I__5876\ : Span4Mux_s0_h
    port map (
            O => \N__31365\,
            I => \N__31362\
        );

    \I__5875\ : Span4Mux_h
    port map (
            O => \N__31362\,
            I => \N__31357\
        );

    \I__5874\ : InMux
    port map (
            O => \N__31361\,
            I => \N__31354\
        );

    \I__5873\ : InMux
    port map (
            O => \N__31360\,
            I => \N__31351\
        );

    \I__5872\ : Span4Mux_h
    port map (
            O => \N__31357\,
            I => \N__31346\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__31354\,
            I => \N__31346\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__31351\,
            I => pin_out_2
        );

    \I__5869\ : Odrv4
    port map (
            O => \N__31346\,
            I => pin_out_2
        );

    \I__5868\ : InMux
    port map (
            O => \N__31341\,
            I => \N__31338\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__31338\,
            I => n13147
        );

    \I__5866\ : InMux
    port map (
            O => \N__31335\,
            I => \N__31332\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__31332\,
            I => n13168
        );

    \I__5864\ : CascadeMux
    port map (
            O => \N__31329\,
            I => \n13167_cascade_\
        );

    \I__5863\ : InMux
    port map (
            O => \N__31326\,
            I => \N__31323\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__31323\,
            I => \N__31320\
        );

    \I__5861\ : Odrv12
    port map (
            O => \N__31320\,
            I => n13450
        );

    \I__5860\ : InMux
    port map (
            O => \N__31317\,
            I => \N__31313\
        );

    \I__5859\ : InMux
    port map (
            O => \N__31316\,
            I => \N__31309\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__31313\,
            I => \N__31306\
        );

    \I__5857\ : InMux
    port map (
            O => \N__31312\,
            I => \N__31303\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__31309\,
            I => \N__31300\
        );

    \I__5855\ : Span4Mux_v
    port map (
            O => \N__31306\,
            I => \N__31295\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__31303\,
            I => \N__31295\
        );

    \I__5853\ : Span4Mux_v
    port map (
            O => \N__31300\,
            I => \N__31290\
        );

    \I__5852\ : Span4Mux_h
    port map (
            O => \N__31295\,
            I => \N__31290\
        );

    \I__5851\ : Odrv4
    port map (
            O => \N__31290\,
            I => \nx.n2694\
        );

    \I__5850\ : CascadeMux
    port map (
            O => \N__31287\,
            I => \N__31283\
        );

    \I__5849\ : CascadeMux
    port map (
            O => \N__31286\,
            I => \N__31279\
        );

    \I__5848\ : InMux
    port map (
            O => \N__31283\,
            I => \N__31276\
        );

    \I__5847\ : InMux
    port map (
            O => \N__31282\,
            I => \N__31271\
        );

    \I__5846\ : InMux
    port map (
            O => \N__31279\,
            I => \N__31271\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__31276\,
            I => \N__31268\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__31271\,
            I => \N__31265\
        );

    \I__5843\ : Span4Mux_h
    port map (
            O => \N__31268\,
            I => \N__31262\
        );

    \I__5842\ : Odrv12
    port map (
            O => \N__31265\,
            I => \nx.n2697\
        );

    \I__5841\ : Odrv4
    port map (
            O => \N__31262\,
            I => \nx.n2697\
        );

    \I__5840\ : CascadeMux
    port map (
            O => \N__31257\,
            I => \n7258_cascade_\
        );

    \I__5839\ : InMux
    port map (
            O => \N__31254\,
            I => \N__31251\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__31251\,
            I => \N__31248\
        );

    \I__5837\ : Odrv4
    port map (
            O => \N__31248\,
            I => n7236
        );

    \I__5836\ : CascadeMux
    port map (
            O => \N__31245\,
            I => \n7270_cascade_\
        );

    \I__5835\ : InMux
    port map (
            O => \N__31242\,
            I => \N__31239\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__31239\,
            I => \N__31236\
        );

    \I__5833\ : Span4Mux_h
    port map (
            O => \N__31236\,
            I => \N__31233\
        );

    \I__5832\ : Odrv4
    port map (
            O => \N__31233\,
            I => n7254
        );

    \I__5831\ : IoInMux
    port map (
            O => \N__31230\,
            I => \N__31227\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__31227\,
            I => \N__31224\
        );

    \I__5829\ : IoSpan4Mux
    port map (
            O => \N__31224\,
            I => \N__31221\
        );

    \I__5828\ : Sp12to4
    port map (
            O => \N__31221\,
            I => \N__31218\
        );

    \I__5827\ : Span12Mux_s6_h
    port map (
            O => \N__31218\,
            I => \N__31215\
        );

    \I__5826\ : Span12Mux_v
    port map (
            O => \N__31215\,
            I => \N__31210\
        );

    \I__5825\ : InMux
    port map (
            O => \N__31214\,
            I => \N__31207\
        );

    \I__5824\ : InMux
    port map (
            O => \N__31213\,
            I => \N__31204\
        );

    \I__5823\ : Odrv12
    port map (
            O => \N__31210\,
            I => pin_out_5
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__31207\,
            I => pin_out_5
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__31204\,
            I => pin_out_5
        );

    \I__5820\ : CascadeMux
    port map (
            O => \N__31197\,
            I => \n13152_cascade_\
        );

    \I__5819\ : InMux
    port map (
            O => \N__31194\,
            I => \nx.n10608\
        );

    \I__5818\ : CascadeMux
    port map (
            O => \N__31191\,
            I => \N__31188\
        );

    \I__5817\ : InMux
    port map (
            O => \N__31188\,
            I => \N__31183\
        );

    \I__5816\ : InMux
    port map (
            O => \N__31187\,
            I => \N__31178\
        );

    \I__5815\ : InMux
    port map (
            O => \N__31186\,
            I => \N__31178\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__31183\,
            I => \nx.n1603\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__31178\,
            I => \nx.n1603\
        );

    \I__5812\ : CascadeMux
    port map (
            O => \N__31173\,
            I => \N__31170\
        );

    \I__5811\ : InMux
    port map (
            O => \N__31170\,
            I => \N__31167\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__31167\,
            I => \nx.n1670\
        );

    \I__5809\ : InMux
    port map (
            O => \N__31164\,
            I => \nx.n10609\
        );

    \I__5808\ : CascadeMux
    port map (
            O => \N__31161\,
            I => \N__31157\
        );

    \I__5807\ : CascadeMux
    port map (
            O => \N__31160\,
            I => \N__31153\
        );

    \I__5806\ : InMux
    port map (
            O => \N__31157\,
            I => \N__31150\
        );

    \I__5805\ : InMux
    port map (
            O => \N__31156\,
            I => \N__31147\
        );

    \I__5804\ : InMux
    port map (
            O => \N__31153\,
            I => \N__31144\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__31150\,
            I => \N__31141\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__31147\,
            I => \N__31138\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__31144\,
            I => \nx.n1602\
        );

    \I__5800\ : Odrv4
    port map (
            O => \N__31141\,
            I => \nx.n1602\
        );

    \I__5799\ : Odrv4
    port map (
            O => \N__31138\,
            I => \nx.n1602\
        );

    \I__5798\ : InMux
    port map (
            O => \N__31131\,
            I => \N__31128\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__31128\,
            I => \N__31125\
        );

    \I__5796\ : Odrv4
    port map (
            O => \N__31125\,
            I => \nx.n1669\
        );

    \I__5795\ : InMux
    port map (
            O => \N__31122\,
            I => \bfn_7_31_0_\
        );

    \I__5794\ : InMux
    port map (
            O => \N__31119\,
            I => \nx.n10611\
        );

    \I__5793\ : InMux
    port map (
            O => \N__31116\,
            I => \nx.n10612\
        );

    \I__5792\ : CascadeMux
    port map (
            O => \N__31113\,
            I => \N__31110\
        );

    \I__5791\ : InMux
    port map (
            O => \N__31110\,
            I => \N__31106\
        );

    \I__5790\ : InMux
    port map (
            O => \N__31109\,
            I => \N__31103\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__31106\,
            I => \nx.n1599\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__31103\,
            I => \nx.n1599\
        );

    \I__5787\ : InMux
    port map (
            O => \N__31098\,
            I => \N__31095\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__31095\,
            I => \nx.n1666\
        );

    \I__5785\ : InMux
    port map (
            O => \N__31092\,
            I => \nx.n10613\
        );

    \I__5784\ : InMux
    port map (
            O => \N__31089\,
            I => \N__31085\
        );

    \I__5783\ : InMux
    port map (
            O => \N__31088\,
            I => \N__31082\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__31085\,
            I => \N__31079\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__31082\,
            I => \nx.n1598\
        );

    \I__5780\ : Odrv4
    port map (
            O => \N__31079\,
            I => \nx.n1598\
        );

    \I__5779\ : InMux
    port map (
            O => \N__31074\,
            I => \nx.n10614\
        );

    \I__5778\ : CascadeMux
    port map (
            O => \N__31071\,
            I => \N__31066\
        );

    \I__5777\ : CascadeMux
    port map (
            O => \N__31070\,
            I => \N__31063\
        );

    \I__5776\ : InMux
    port map (
            O => \N__31069\,
            I => \N__31058\
        );

    \I__5775\ : InMux
    port map (
            O => \N__31066\,
            I => \N__31058\
        );

    \I__5774\ : InMux
    port map (
            O => \N__31063\,
            I => \N__31055\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__31058\,
            I => \nx.n1600\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__31055\,
            I => \nx.n1600\
        );

    \I__5771\ : CascadeMux
    port map (
            O => \N__31050\,
            I => \N__31047\
        );

    \I__5770\ : InMux
    port map (
            O => \N__31047\,
            I => \N__31044\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__31044\,
            I => \nx.n1667\
        );

    \I__5768\ : InMux
    port map (
            O => \N__31041\,
            I => \N__31038\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__31038\,
            I => \N__31035\
        );

    \I__5766\ : Odrv4
    port map (
            O => \N__31035\,
            I => \nx.n1570\
        );

    \I__5765\ : CascadeMux
    port map (
            O => \N__31032\,
            I => \N__31028\
        );

    \I__5764\ : InMux
    port map (
            O => \N__31031\,
            I => \N__31025\
        );

    \I__5763\ : InMux
    port map (
            O => \N__31028\,
            I => \N__31022\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__31025\,
            I => \N__31017\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__31022\,
            I => \N__31017\
        );

    \I__5760\ : Span4Mux_v
    port map (
            O => \N__31017\,
            I => \N__31013\
        );

    \I__5759\ : InMux
    port map (
            O => \N__31016\,
            I => \N__31010\
        );

    \I__5758\ : Odrv4
    port map (
            O => \N__31013\,
            I => \nx.n1503\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__31010\,
            I => \nx.n1503\
        );

    \I__5756\ : InMux
    port map (
            O => \N__31005\,
            I => \N__31000\
        );

    \I__5755\ : InMux
    port map (
            O => \N__31004\,
            I => \N__30996\
        );

    \I__5754\ : InMux
    port map (
            O => \N__31003\,
            I => \N__30992\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__31000\,
            I => \N__30989\
        );

    \I__5752\ : InMux
    port map (
            O => \N__30999\,
            I => \N__30986\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__30996\,
            I => \N__30983\
        );

    \I__5750\ : InMux
    port map (
            O => \N__30995\,
            I => \N__30980\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__30992\,
            I => \N__30977\
        );

    \I__5748\ : Span4Mux_h
    port map (
            O => \N__30989\,
            I => \N__30974\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__30986\,
            I => \N__30971\
        );

    \I__5746\ : Span4Mux_h
    port map (
            O => \N__30983\,
            I => \N__30968\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__30980\,
            I => \nx.bit_ctr_19\
        );

    \I__5744\ : Odrv4
    port map (
            O => \N__30977\,
            I => \nx.bit_ctr_19\
        );

    \I__5743\ : Odrv4
    port map (
            O => \N__30974\,
            I => \nx.bit_ctr_19\
        );

    \I__5742\ : Odrv4
    port map (
            O => \N__30971\,
            I => \nx.bit_ctr_19\
        );

    \I__5741\ : Odrv4
    port map (
            O => \N__30968\,
            I => \nx.bit_ctr_19\
        );

    \I__5740\ : InMux
    port map (
            O => \N__30957\,
            I => \N__30954\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__30954\,
            I => \N__30951\
        );

    \I__5738\ : Span4Mux_h
    port map (
            O => \N__30951\,
            I => \N__30948\
        );

    \I__5737\ : Odrv4
    port map (
            O => \N__30948\,
            I => \nx.n1677\
        );

    \I__5736\ : InMux
    port map (
            O => \N__30945\,
            I => \bfn_7_30_0_\
        );

    \I__5735\ : CascadeMux
    port map (
            O => \N__30942\,
            I => \N__30938\
        );

    \I__5734\ : InMux
    port map (
            O => \N__30941\,
            I => \N__30935\
        );

    \I__5733\ : InMux
    port map (
            O => \N__30938\,
            I => \N__30932\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__30935\,
            I => \nx.n1609\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__30932\,
            I => \nx.n1609\
        );

    \I__5730\ : InMux
    port map (
            O => \N__30927\,
            I => \N__30924\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__30924\,
            I => \nx.n1676\
        );

    \I__5728\ : InMux
    port map (
            O => \N__30921\,
            I => \nx.n10603\
        );

    \I__5727\ : InMux
    port map (
            O => \N__30918\,
            I => \nx.n10604\
        );

    \I__5726\ : CascadeMux
    port map (
            O => \N__30915\,
            I => \N__30911\
        );

    \I__5725\ : CascadeMux
    port map (
            O => \N__30914\,
            I => \N__30907\
        );

    \I__5724\ : InMux
    port map (
            O => \N__30911\,
            I => \N__30904\
        );

    \I__5723\ : InMux
    port map (
            O => \N__30910\,
            I => \N__30901\
        );

    \I__5722\ : InMux
    port map (
            O => \N__30907\,
            I => \N__30898\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__30904\,
            I => \nx.n1607\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__30901\,
            I => \nx.n1607\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__30898\,
            I => \nx.n1607\
        );

    \I__5718\ : InMux
    port map (
            O => \N__30891\,
            I => \N__30888\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__30888\,
            I => \N__30885\
        );

    \I__5716\ : Odrv4
    port map (
            O => \N__30885\,
            I => \nx.n1674\
        );

    \I__5715\ : InMux
    port map (
            O => \N__30882\,
            I => \nx.n10605\
        );

    \I__5714\ : InMux
    port map (
            O => \N__30879\,
            I => \nx.n10606\
        );

    \I__5713\ : InMux
    port map (
            O => \N__30876\,
            I => \N__30873\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__30873\,
            I => \nx.n1672\
        );

    \I__5711\ : InMux
    port map (
            O => \N__30870\,
            I => \nx.n10607\
        );

    \I__5710\ : CascadeMux
    port map (
            O => \N__30867\,
            I => \nx.n1701_cascade_\
        );

    \I__5709\ : CascadeMux
    port map (
            O => \N__30864\,
            I => \nx.n1801_cascade_\
        );

    \I__5708\ : InMux
    port map (
            O => \N__30861\,
            I => \N__30858\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__30858\,
            I => \nx.n23\
        );

    \I__5706\ : InMux
    port map (
            O => \N__30855\,
            I => \N__30852\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__30852\,
            I => \N__30849\
        );

    \I__5704\ : Odrv4
    port map (
            O => \N__30849\,
            I => \nx.n1577\
        );

    \I__5703\ : InMux
    port map (
            O => \N__30846\,
            I => \N__30841\
        );

    \I__5702\ : InMux
    port map (
            O => \N__30845\,
            I => \N__30838\
        );

    \I__5701\ : InMux
    port map (
            O => \N__30844\,
            I => \N__30833\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__30841\,
            I => \N__30828\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__30838\,
            I => \N__30828\
        );

    \I__5698\ : InMux
    port map (
            O => \N__30837\,
            I => \N__30825\
        );

    \I__5697\ : InMux
    port map (
            O => \N__30836\,
            I => \N__30822\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__30833\,
            I => \N__30819\
        );

    \I__5695\ : Span4Mux_h
    port map (
            O => \N__30828\,
            I => \N__30816\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__30825\,
            I => \N__30813\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__30822\,
            I => \nx.bit_ctr_20\
        );

    \I__5692\ : Odrv4
    port map (
            O => \N__30819\,
            I => \nx.bit_ctr_20\
        );

    \I__5691\ : Odrv4
    port map (
            O => \N__30816\,
            I => \nx.bit_ctr_20\
        );

    \I__5690\ : Odrv12
    port map (
            O => \N__30813\,
            I => \nx.bit_ctr_20\
        );

    \I__5689\ : CascadeMux
    port map (
            O => \N__30804\,
            I => \nx.n1609_cascade_\
        );

    \I__5688\ : InMux
    port map (
            O => \N__30801\,
            I => \N__30798\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__30798\,
            I => \nx.n16_adj_646\
        );

    \I__5686\ : InMux
    port map (
            O => \N__30795\,
            I => \nx.n10653\
        );

    \I__5685\ : InMux
    port map (
            O => \N__30792\,
            I => \nx.n10654\
        );

    \I__5684\ : InMux
    port map (
            O => \N__30789\,
            I => \nx.n10655\
        );

    \I__5683\ : CascadeMux
    port map (
            O => \N__30786\,
            I => \N__30770\
        );

    \I__5682\ : CascadeMux
    port map (
            O => \N__30785\,
            I => \N__30767\
        );

    \I__5681\ : CascadeMux
    port map (
            O => \N__30784\,
            I => \N__30764\
        );

    \I__5680\ : CascadeMux
    port map (
            O => \N__30783\,
            I => \N__30761\
        );

    \I__5679\ : CascadeMux
    port map (
            O => \N__30782\,
            I => \N__30758\
        );

    \I__5678\ : CascadeMux
    port map (
            O => \N__30781\,
            I => \N__30755\
        );

    \I__5677\ : CascadeMux
    port map (
            O => \N__30780\,
            I => \N__30752\
        );

    \I__5676\ : CascadeMux
    port map (
            O => \N__30779\,
            I => \N__30749\
        );

    \I__5675\ : CascadeMux
    port map (
            O => \N__30778\,
            I => \N__30746\
        );

    \I__5674\ : CascadeMux
    port map (
            O => \N__30777\,
            I => \N__30743\
        );

    \I__5673\ : CascadeMux
    port map (
            O => \N__30776\,
            I => \N__30740\
        );

    \I__5672\ : CascadeMux
    port map (
            O => \N__30775\,
            I => \N__30737\
        );

    \I__5671\ : CascadeMux
    port map (
            O => \N__30774\,
            I => \N__30734\
        );

    \I__5670\ : CascadeMux
    port map (
            O => \N__30773\,
            I => \N__30731\
        );

    \I__5669\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30722\
        );

    \I__5668\ : InMux
    port map (
            O => \N__30767\,
            I => \N__30722\
        );

    \I__5667\ : InMux
    port map (
            O => \N__30764\,
            I => \N__30722\
        );

    \I__5666\ : InMux
    port map (
            O => \N__30761\,
            I => \N__30722\
        );

    \I__5665\ : InMux
    port map (
            O => \N__30758\,
            I => \N__30713\
        );

    \I__5664\ : InMux
    port map (
            O => \N__30755\,
            I => \N__30713\
        );

    \I__5663\ : InMux
    port map (
            O => \N__30752\,
            I => \N__30713\
        );

    \I__5662\ : InMux
    port map (
            O => \N__30749\,
            I => \N__30713\
        );

    \I__5661\ : InMux
    port map (
            O => \N__30746\,
            I => \N__30706\
        );

    \I__5660\ : InMux
    port map (
            O => \N__30743\,
            I => \N__30706\
        );

    \I__5659\ : InMux
    port map (
            O => \N__30740\,
            I => \N__30706\
        );

    \I__5658\ : InMux
    port map (
            O => \N__30737\,
            I => \N__30699\
        );

    \I__5657\ : InMux
    port map (
            O => \N__30734\,
            I => \N__30699\
        );

    \I__5656\ : InMux
    port map (
            O => \N__30731\,
            I => \N__30699\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__30722\,
            I => \nx.n1928\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__30713\,
            I => \nx.n1928\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__30706\,
            I => \nx.n1928\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__30699\,
            I => \nx.n1928\
        );

    \I__5651\ : InMux
    port map (
            O => \N__30690\,
            I => \nx.n10656\
        );

    \I__5650\ : InMux
    port map (
            O => \N__30687\,
            I => \N__30682\
        );

    \I__5649\ : InMux
    port map (
            O => \N__30686\,
            I => \N__30679\
        );

    \I__5648\ : InMux
    port map (
            O => \N__30685\,
            I => \N__30676\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__30682\,
            I => \N__30673\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__30679\,
            I => \nx.n1897\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__30676\,
            I => \nx.n1897\
        );

    \I__5644\ : Odrv4
    port map (
            O => \N__30673\,
            I => \nx.n1897\
        );

    \I__5643\ : InMux
    port map (
            O => \N__30666\,
            I => \N__30662\
        );

    \I__5642\ : InMux
    port map (
            O => \N__30665\,
            I => \N__30659\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__30662\,
            I => \N__30653\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__30659\,
            I => \N__30653\
        );

    \I__5639\ : InMux
    port map (
            O => \N__30658\,
            I => \N__30650\
        );

    \I__5638\ : Odrv4
    port map (
            O => \N__30653\,
            I => \nx.n1902\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__30650\,
            I => \nx.n1902\
        );

    \I__5636\ : CascadeMux
    port map (
            O => \N__30645\,
            I => \N__30640\
        );

    \I__5635\ : InMux
    port map (
            O => \N__30644\,
            I => \N__30636\
        );

    \I__5634\ : InMux
    port map (
            O => \N__30643\,
            I => \N__30633\
        );

    \I__5633\ : InMux
    port map (
            O => \N__30640\,
            I => \N__30628\
        );

    \I__5632\ : InMux
    port map (
            O => \N__30639\,
            I => \N__30628\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__30636\,
            I => \N__30622\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__30633\,
            I => \N__30619\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__30628\,
            I => \N__30616\
        );

    \I__5628\ : InMux
    port map (
            O => \N__30627\,
            I => \N__30609\
        );

    \I__5627\ : InMux
    port map (
            O => \N__30626\,
            I => \N__30609\
        );

    \I__5626\ : InMux
    port map (
            O => \N__30625\,
            I => \N__30609\
        );

    \I__5625\ : Span4Mux_h
    port map (
            O => \N__30622\,
            I => \N__30606\
        );

    \I__5624\ : Odrv4
    port map (
            O => \N__30619\,
            I => \nx.n10994\
        );

    \I__5623\ : Odrv4
    port map (
            O => \N__30616\,
            I => \nx.n10994\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__30609\,
            I => \nx.n10994\
        );

    \I__5621\ : Odrv4
    port map (
            O => \N__30606\,
            I => \nx.n10994\
        );

    \I__5620\ : InMux
    port map (
            O => \N__30597\,
            I => \N__30594\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__30594\,
            I => \nx.n13425\
        );

    \I__5618\ : InMux
    port map (
            O => \N__30591\,
            I => \N__30587\
        );

    \I__5617\ : InMux
    port map (
            O => \N__30590\,
            I => \N__30584\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__30587\,
            I => \nx.n1906\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__30584\,
            I => \nx.n1906\
        );

    \I__5614\ : InMux
    port map (
            O => \N__30579\,
            I => \nx.n10645\
        );

    \I__5613\ : InMux
    port map (
            O => \N__30576\,
            I => \nx.n10646\
        );

    \I__5612\ : CascadeMux
    port map (
            O => \N__30573\,
            I => \N__30568\
        );

    \I__5611\ : InMux
    port map (
            O => \N__30572\,
            I => \N__30565\
        );

    \I__5610\ : InMux
    port map (
            O => \N__30571\,
            I => \N__30562\
        );

    \I__5609\ : InMux
    port map (
            O => \N__30568\,
            I => \N__30559\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__30565\,
            I => \nx.n1904\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__30562\,
            I => \nx.n1904\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__30559\,
            I => \nx.n1904\
        );

    \I__5605\ : InMux
    port map (
            O => \N__30552\,
            I => \nx.n10647\
        );

    \I__5604\ : InMux
    port map (
            O => \N__30549\,
            I => \N__30544\
        );

    \I__5603\ : InMux
    port map (
            O => \N__30548\,
            I => \N__30541\
        );

    \I__5602\ : InMux
    port map (
            O => \N__30547\,
            I => \N__30538\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__30544\,
            I => \nx.n1903\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__30541\,
            I => \nx.n1903\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__30538\,
            I => \nx.n1903\
        );

    \I__5598\ : InMux
    port map (
            O => \N__30531\,
            I => \nx.n10648\
        );

    \I__5597\ : InMux
    port map (
            O => \N__30528\,
            I => \bfn_7_26_0_\
        );

    \I__5596\ : InMux
    port map (
            O => \N__30525\,
            I => \nx.n10650\
        );

    \I__5595\ : InMux
    port map (
            O => \N__30522\,
            I => \nx.n10651\
        );

    \I__5594\ : InMux
    port map (
            O => \N__30519\,
            I => \N__30514\
        );

    \I__5593\ : InMux
    port map (
            O => \N__30518\,
            I => \N__30511\
        );

    \I__5592\ : InMux
    port map (
            O => \N__30517\,
            I => \N__30508\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__30514\,
            I => \N__30505\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__30511\,
            I => \nx.n1899\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__30508\,
            I => \nx.n1899\
        );

    \I__5588\ : Odrv4
    port map (
            O => \N__30505\,
            I => \nx.n1899\
        );

    \I__5587\ : InMux
    port map (
            O => \N__30498\,
            I => \nx.n10652\
        );

    \I__5586\ : CascadeMux
    port map (
            O => \N__30495\,
            I => \N__30492\
        );

    \I__5585\ : InMux
    port map (
            O => \N__30492\,
            I => \N__30489\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__30489\,
            I => \N__30485\
        );

    \I__5583\ : CascadeMux
    port map (
            O => \N__30488\,
            I => \N__30482\
        );

    \I__5582\ : Span4Mux_v
    port map (
            O => \N__30485\,
            I => \N__30478\
        );

    \I__5581\ : InMux
    port map (
            O => \N__30482\,
            I => \N__30475\
        );

    \I__5580\ : InMux
    port map (
            O => \N__30481\,
            I => \N__30472\
        );

    \I__5579\ : Odrv4
    port map (
            O => \N__30478\,
            I => \nx.n2888\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__30475\,
            I => \nx.n2888\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__30472\,
            I => \nx.n2888\
        );

    \I__5576\ : CascadeMux
    port map (
            O => \N__30465\,
            I => \nx.n2887_cascade_\
        );

    \I__5575\ : InMux
    port map (
            O => \N__30462\,
            I => \N__30459\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__30459\,
            I => \N__30456\
        );

    \I__5573\ : Span4Mux_h
    port map (
            O => \N__30456\,
            I => \N__30453\
        );

    \I__5572\ : Odrv4
    port map (
            O => \N__30453\,
            I => \nx.n39_adj_679\
        );

    \I__5571\ : InMux
    port map (
            O => \N__30450\,
            I => \N__30447\
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__30447\,
            I => \N__30443\
        );

    \I__5569\ : CascadeMux
    port map (
            O => \N__30446\,
            I => \N__30439\
        );

    \I__5568\ : Span4Mux_v
    port map (
            O => \N__30443\,
            I => \N__30436\
        );

    \I__5567\ : InMux
    port map (
            O => \N__30442\,
            I => \N__30433\
        );

    \I__5566\ : InMux
    port map (
            O => \N__30439\,
            I => \N__30430\
        );

    \I__5565\ : Odrv4
    port map (
            O => \N__30436\,
            I => \nx.n2803\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__30433\,
            I => \nx.n2803\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__30430\,
            I => \nx.n2803\
        );

    \I__5562\ : InMux
    port map (
            O => \N__30423\,
            I => \N__30420\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__30420\,
            I => \N__30417\
        );

    \I__5560\ : Span4Mux_h
    port map (
            O => \N__30417\,
            I => \N__30414\
        );

    \I__5559\ : Odrv4
    port map (
            O => \N__30414\,
            I => \nx.n2870\
        );

    \I__5558\ : InMux
    port map (
            O => \N__30411\,
            I => \N__30406\
        );

    \I__5557\ : CascadeMux
    port map (
            O => \N__30410\,
            I => \N__30403\
        );

    \I__5556\ : CascadeMux
    port map (
            O => \N__30409\,
            I => \N__30400\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__30406\,
            I => \N__30397\
        );

    \I__5554\ : InMux
    port map (
            O => \N__30403\,
            I => \N__30394\
        );

    \I__5553\ : InMux
    port map (
            O => \N__30400\,
            I => \N__30391\
        );

    \I__5552\ : Span4Mux_s2_h
    port map (
            O => \N__30397\,
            I => \N__30384\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__30394\,
            I => \N__30384\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__30391\,
            I => \N__30384\
        );

    \I__5549\ : Span4Mux_h
    port map (
            O => \N__30384\,
            I => \N__30381\
        );

    \I__5548\ : Odrv4
    port map (
            O => \N__30381\,
            I => \nx.n2902\
        );

    \I__5547\ : InMux
    port map (
            O => \N__30378\,
            I => \N__30375\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__30375\,
            I => \N__30372\
        );

    \I__5545\ : Odrv4
    port map (
            O => \N__30372\,
            I => \nx.n2871\
        );

    \I__5544\ : CascadeMux
    port map (
            O => \N__30369\,
            I => \N__30365\
        );

    \I__5543\ : CascadeMux
    port map (
            O => \N__30368\,
            I => \N__30362\
        );

    \I__5542\ : InMux
    port map (
            O => \N__30365\,
            I => \N__30358\
        );

    \I__5541\ : InMux
    port map (
            O => \N__30362\,
            I => \N__30355\
        );

    \I__5540\ : InMux
    port map (
            O => \N__30361\,
            I => \N__30352\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__30358\,
            I => \N__30349\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__30355\,
            I => \N__30346\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__30352\,
            I => \N__30343\
        );

    \I__5536\ : Span4Mux_h
    port map (
            O => \N__30349\,
            I => \N__30340\
        );

    \I__5535\ : Span4Mux_h
    port map (
            O => \N__30346\,
            I => \N__30337\
        );

    \I__5534\ : Odrv4
    port map (
            O => \N__30343\,
            I => \nx.n2903\
        );

    \I__5533\ : Odrv4
    port map (
            O => \N__30340\,
            I => \nx.n2903\
        );

    \I__5532\ : Odrv4
    port map (
            O => \N__30337\,
            I => \nx.n2903\
        );

    \I__5531\ : InMux
    port map (
            O => \N__30330\,
            I => \N__30326\
        );

    \I__5530\ : CascadeMux
    port map (
            O => \N__30329\,
            I => \N__30323\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__30326\,
            I => \N__30319\
        );

    \I__5528\ : InMux
    port map (
            O => \N__30323\,
            I => \N__30316\
        );

    \I__5527\ : InMux
    port map (
            O => \N__30322\,
            I => \N__30313\
        );

    \I__5526\ : Odrv4
    port map (
            O => \N__30319\,
            I => \nx.n2790\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__30316\,
            I => \nx.n2790\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__30313\,
            I => \nx.n2790\
        );

    \I__5523\ : CascadeMux
    port map (
            O => \N__30306\,
            I => \N__30298\
        );

    \I__5522\ : CascadeMux
    port map (
            O => \N__30305\,
            I => \N__30295\
        );

    \I__5521\ : CascadeMux
    port map (
            O => \N__30304\,
            I => \N__30290\
        );

    \I__5520\ : CascadeMux
    port map (
            O => \N__30303\,
            I => \N__30287\
        );

    \I__5519\ : InMux
    port map (
            O => \N__30302\,
            I => \N__30278\
        );

    \I__5518\ : InMux
    port map (
            O => \N__30301\,
            I => \N__30278\
        );

    \I__5517\ : InMux
    port map (
            O => \N__30298\,
            I => \N__30263\
        );

    \I__5516\ : InMux
    port map (
            O => \N__30295\,
            I => \N__30263\
        );

    \I__5515\ : InMux
    port map (
            O => \N__30294\,
            I => \N__30263\
        );

    \I__5514\ : InMux
    port map (
            O => \N__30293\,
            I => \N__30263\
        );

    \I__5513\ : InMux
    port map (
            O => \N__30290\,
            I => \N__30263\
        );

    \I__5512\ : InMux
    port map (
            O => \N__30287\,
            I => \N__30258\
        );

    \I__5511\ : InMux
    port map (
            O => \N__30286\,
            I => \N__30258\
        );

    \I__5510\ : CascadeMux
    port map (
            O => \N__30285\,
            I => \N__30252\
        );

    \I__5509\ : CascadeMux
    port map (
            O => \N__30284\,
            I => \N__30247\
        );

    \I__5508\ : CascadeMux
    port map (
            O => \N__30283\,
            I => \N__30243\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__30278\,
            I => \N__30240\
        );

    \I__5506\ : CascadeMux
    port map (
            O => \N__30277\,
            I => \N__30237\
        );

    \I__5505\ : CascadeMux
    port map (
            O => \N__30276\,
            I => \N__30234\
        );

    \I__5504\ : CascadeMux
    port map (
            O => \N__30275\,
            I => \N__30231\
        );

    \I__5503\ : CascadeMux
    port map (
            O => \N__30274\,
            I => \N__30228\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__30263\,
            I => \N__30224\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__30258\,
            I => \N__30221\
        );

    \I__5500\ : InMux
    port map (
            O => \N__30257\,
            I => \N__30218\
        );

    \I__5499\ : CascadeMux
    port map (
            O => \N__30256\,
            I => \N__30215\
        );

    \I__5498\ : CascadeMux
    port map (
            O => \N__30255\,
            I => \N__30212\
        );

    \I__5497\ : InMux
    port map (
            O => \N__30252\,
            I => \N__30206\
        );

    \I__5496\ : InMux
    port map (
            O => \N__30251\,
            I => \N__30206\
        );

    \I__5495\ : InMux
    port map (
            O => \N__30250\,
            I => \N__30197\
        );

    \I__5494\ : InMux
    port map (
            O => \N__30247\,
            I => \N__30197\
        );

    \I__5493\ : InMux
    port map (
            O => \N__30246\,
            I => \N__30197\
        );

    \I__5492\ : InMux
    port map (
            O => \N__30243\,
            I => \N__30197\
        );

    \I__5491\ : Span4Mux_h
    port map (
            O => \N__30240\,
            I => \N__30194\
        );

    \I__5490\ : InMux
    port map (
            O => \N__30237\,
            I => \N__30183\
        );

    \I__5489\ : InMux
    port map (
            O => \N__30234\,
            I => \N__30183\
        );

    \I__5488\ : InMux
    port map (
            O => \N__30231\,
            I => \N__30183\
        );

    \I__5487\ : InMux
    port map (
            O => \N__30228\,
            I => \N__30183\
        );

    \I__5486\ : InMux
    port map (
            O => \N__30227\,
            I => \N__30183\
        );

    \I__5485\ : Span4Mux_v
    port map (
            O => \N__30224\,
            I => \N__30180\
        );

    \I__5484\ : Span4Mux_h
    port map (
            O => \N__30221\,
            I => \N__30177\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__30218\,
            I => \N__30174\
        );

    \I__5482\ : InMux
    port map (
            O => \N__30215\,
            I => \N__30167\
        );

    \I__5481\ : InMux
    port map (
            O => \N__30212\,
            I => \N__30167\
        );

    \I__5480\ : InMux
    port map (
            O => \N__30211\,
            I => \N__30167\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__30206\,
            I => \nx.n2819\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__30197\,
            I => \nx.n2819\
        );

    \I__5477\ : Odrv4
    port map (
            O => \N__30194\,
            I => \nx.n2819\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__30183\,
            I => \nx.n2819\
        );

    \I__5475\ : Odrv4
    port map (
            O => \N__30180\,
            I => \nx.n2819\
        );

    \I__5474\ : Odrv4
    port map (
            O => \N__30177\,
            I => \nx.n2819\
        );

    \I__5473\ : Odrv12
    port map (
            O => \N__30174\,
            I => \nx.n2819\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__30167\,
            I => \nx.n2819\
        );

    \I__5471\ : InMux
    port map (
            O => \N__30150\,
            I => \N__30147\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__30147\,
            I => \nx.n2857\
        );

    \I__5469\ : InMux
    port map (
            O => \N__30144\,
            I => \N__30140\
        );

    \I__5468\ : CascadeMux
    port map (
            O => \N__30143\,
            I => \N__30137\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__30140\,
            I => \N__30134\
        );

    \I__5466\ : InMux
    port map (
            O => \N__30137\,
            I => \N__30131\
        );

    \I__5465\ : Span4Mux_v
    port map (
            O => \N__30134\,
            I => \N__30125\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__30131\,
            I => \N__30125\
        );

    \I__5463\ : InMux
    port map (
            O => \N__30130\,
            I => \N__30122\
        );

    \I__5462\ : Odrv4
    port map (
            O => \N__30125\,
            I => \nx.n2889\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__30122\,
            I => \nx.n2889\
        );

    \I__5460\ : InMux
    port map (
            O => \N__30117\,
            I => \N__30112\
        );

    \I__5459\ : InMux
    port map (
            O => \N__30116\,
            I => \N__30109\
        );

    \I__5458\ : CascadeMux
    port map (
            O => \N__30115\,
            I => \N__30105\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__30112\,
            I => \N__30100\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__30109\,
            I => \N__30100\
        );

    \I__5455\ : InMux
    port map (
            O => \N__30108\,
            I => \N__30097\
        );

    \I__5454\ : InMux
    port map (
            O => \N__30105\,
            I => \N__30093\
        );

    \I__5453\ : Span4Mux_h
    port map (
            O => \N__30100\,
            I => \N__30090\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__30097\,
            I => \N__30087\
        );

    \I__5451\ : InMux
    port map (
            O => \N__30096\,
            I => \N__30084\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__30093\,
            I => \N__30081\
        );

    \I__5449\ : Span4Mux_s3_h
    port map (
            O => \N__30090\,
            I => \N__30078\
        );

    \I__5448\ : Span4Mux_v
    port map (
            O => \N__30087\,
            I => \N__30075\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__30084\,
            I => \nx.bit_ctr_16\
        );

    \I__5446\ : Odrv4
    port map (
            O => \N__30081\,
            I => \nx.bit_ctr_16\
        );

    \I__5445\ : Odrv4
    port map (
            O => \N__30078\,
            I => \nx.bit_ctr_16\
        );

    \I__5444\ : Odrv4
    port map (
            O => \N__30075\,
            I => \nx.bit_ctr_16\
        );

    \I__5443\ : InMux
    port map (
            O => \N__30066\,
            I => \bfn_7_25_0_\
        );

    \I__5442\ : InMux
    port map (
            O => \N__30063\,
            I => \N__30058\
        );

    \I__5441\ : InMux
    port map (
            O => \N__30062\,
            I => \N__30055\
        );

    \I__5440\ : InMux
    port map (
            O => \N__30061\,
            I => \N__30052\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__30058\,
            I => \nx.n1909\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__30055\,
            I => \nx.n1909\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__30052\,
            I => \nx.n1909\
        );

    \I__5436\ : CascadeMux
    port map (
            O => \N__30045\,
            I => \N__30041\
        );

    \I__5435\ : CascadeMux
    port map (
            O => \N__30044\,
            I => \N__30038\
        );

    \I__5434\ : InMux
    port map (
            O => \N__30041\,
            I => \N__30035\
        );

    \I__5433\ : InMux
    port map (
            O => \N__30038\,
            I => \N__30032\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__30035\,
            I => \nx.n13435\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__30032\,
            I => \nx.n13435\
        );

    \I__5430\ : InMux
    port map (
            O => \N__30027\,
            I => \nx.n10642\
        );

    \I__5429\ : InMux
    port map (
            O => \N__30024\,
            I => \N__30020\
        );

    \I__5428\ : InMux
    port map (
            O => \N__30023\,
            I => \N__30017\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__30020\,
            I => \nx.n1908\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__30017\,
            I => \nx.n1908\
        );

    \I__5425\ : InMux
    port map (
            O => \N__30012\,
            I => \nx.n10643\
        );

    \I__5424\ : InMux
    port map (
            O => \N__30009\,
            I => \N__30004\
        );

    \I__5423\ : InMux
    port map (
            O => \N__30008\,
            I => \N__30001\
        );

    \I__5422\ : InMux
    port map (
            O => \N__30007\,
            I => \N__29998\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__30004\,
            I => \nx.n1907\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__30001\,
            I => \nx.n1907\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__29998\,
            I => \nx.n1907\
        );

    \I__5418\ : InMux
    port map (
            O => \N__29991\,
            I => \nx.n10644\
        );

    \I__5417\ : InMux
    port map (
            O => \N__29988\,
            I => \N__29985\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__29985\,
            I => \N__29982\
        );

    \I__5415\ : Span4Mux_h
    port map (
            O => \N__29982\,
            I => \N__29979\
        );

    \I__5414\ : Odrv4
    port map (
            O => \N__29979\,
            I => \nx.n44\
        );

    \I__5413\ : InMux
    port map (
            O => \N__29976\,
            I => \N__29973\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__29973\,
            I => \nx.n2854\
        );

    \I__5411\ : CascadeMux
    port map (
            O => \N__29970\,
            I => \nx.n2819_cascade_\
        );

    \I__5410\ : CascadeMux
    port map (
            O => \N__29967\,
            I => \N__29963\
        );

    \I__5409\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29960\
        );

    \I__5408\ : InMux
    port map (
            O => \N__29963\,
            I => \N__29957\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__29960\,
            I => \N__29953\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__29957\,
            I => \N__29950\
        );

    \I__5405\ : InMux
    port map (
            O => \N__29956\,
            I => \N__29947\
        );

    \I__5404\ : Span4Mux_v
    port map (
            O => \N__29953\,
            I => \N__29944\
        );

    \I__5403\ : Span4Mux_v
    port map (
            O => \N__29950\,
            I => \N__29939\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__29947\,
            I => \N__29939\
        );

    \I__5401\ : Odrv4
    port map (
            O => \N__29944\,
            I => \nx.n2886\
        );

    \I__5400\ : Odrv4
    port map (
            O => \N__29939\,
            I => \nx.n2886\
        );

    \I__5399\ : CascadeMux
    port map (
            O => \N__29934\,
            I => \N__29930\
        );

    \I__5398\ : CascadeMux
    port map (
            O => \N__29933\,
            I => \N__29927\
        );

    \I__5397\ : InMux
    port map (
            O => \N__29930\,
            I => \N__29924\
        );

    \I__5396\ : InMux
    port map (
            O => \N__29927\,
            I => \N__29921\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__29924\,
            I => \nx.n2789\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__29921\,
            I => \nx.n2789\
        );

    \I__5393\ : InMux
    port map (
            O => \N__29916\,
            I => \N__29913\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__29913\,
            I => \nx.n26_adj_615\
        );

    \I__5391\ : InMux
    port map (
            O => \N__29910\,
            I => \N__29907\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__29907\,
            I => \nx.n2863\
        );

    \I__5389\ : InMux
    port map (
            O => \N__29904\,
            I => \N__29900\
        );

    \I__5388\ : CascadeMux
    port map (
            O => \N__29903\,
            I => \N__29897\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__29900\,
            I => \N__29894\
        );

    \I__5386\ : InMux
    port map (
            O => \N__29897\,
            I => \N__29891\
        );

    \I__5385\ : Span4Mux_v
    port map (
            O => \N__29894\,
            I => \N__29887\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__29891\,
            I => \N__29884\
        );

    \I__5383\ : InMux
    port map (
            O => \N__29890\,
            I => \N__29881\
        );

    \I__5382\ : Odrv4
    port map (
            O => \N__29887\,
            I => \nx.n2796\
        );

    \I__5381\ : Odrv12
    port map (
            O => \N__29884\,
            I => \nx.n2796\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__29881\,
            I => \nx.n2796\
        );

    \I__5379\ : InMux
    port map (
            O => \N__29874\,
            I => \N__29869\
        );

    \I__5378\ : CascadeMux
    port map (
            O => \N__29873\,
            I => \N__29866\
        );

    \I__5377\ : InMux
    port map (
            O => \N__29872\,
            I => \N__29863\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__29869\,
            I => \N__29860\
        );

    \I__5375\ : InMux
    port map (
            O => \N__29866\,
            I => \N__29857\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__29863\,
            I => \N__29854\
        );

    \I__5373\ : Span4Mux_v
    port map (
            O => \N__29860\,
            I => \N__29849\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__29857\,
            I => \N__29849\
        );

    \I__5371\ : Span4Mux_h
    port map (
            O => \N__29854\,
            I => \N__29846\
        );

    \I__5370\ : Odrv4
    port map (
            O => \N__29849\,
            I => \nx.n2895\
        );

    \I__5369\ : Odrv4
    port map (
            O => \N__29846\,
            I => \nx.n2895\
        );

    \I__5368\ : InMux
    port map (
            O => \N__29841\,
            I => \N__29838\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__29838\,
            I => \N__29835\
        );

    \I__5366\ : Span4Mux_v
    port map (
            O => \N__29835\,
            I => \N__29832\
        );

    \I__5365\ : Odrv4
    port map (
            O => \N__29832\,
            I => \nx.n2877\
        );

    \I__5364\ : InMux
    port map (
            O => \N__29829\,
            I => \N__29823\
        );

    \I__5363\ : InMux
    port map (
            O => \N__29828\,
            I => \N__29820\
        );

    \I__5362\ : InMux
    port map (
            O => \N__29827\,
            I => \N__29817\
        );

    \I__5361\ : InMux
    port map (
            O => \N__29826\,
            I => \N__29814\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__29823\,
            I => \N__29809\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__29820\,
            I => \N__29809\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__29817\,
            I => \N__29805\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__29814\,
            I => \N__29802\
        );

    \I__5356\ : Span4Mux_v
    port map (
            O => \N__29809\,
            I => \N__29799\
        );

    \I__5355\ : InMux
    port map (
            O => \N__29808\,
            I => \N__29796\
        );

    \I__5354\ : Span12Mux_s5_v
    port map (
            O => \N__29805\,
            I => \N__29791\
        );

    \I__5353\ : Span12Mux_v
    port map (
            O => \N__29802\,
            I => \N__29791\
        );

    \I__5352\ : Span4Mux_v
    port map (
            O => \N__29799\,
            I => \N__29788\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__29796\,
            I => \nx.bit_ctr_7\
        );

    \I__5350\ : Odrv12
    port map (
            O => \N__29791\,
            I => \nx.bit_ctr_7\
        );

    \I__5349\ : Odrv4
    port map (
            O => \N__29788\,
            I => \nx.bit_ctr_7\
        );

    \I__5348\ : CascadeMux
    port map (
            O => \N__29781\,
            I => \N__29778\
        );

    \I__5347\ : InMux
    port map (
            O => \N__29778\,
            I => \N__29773\
        );

    \I__5346\ : InMux
    port map (
            O => \N__29777\,
            I => \N__29770\
        );

    \I__5345\ : InMux
    port map (
            O => \N__29776\,
            I => \N__29767\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__29773\,
            I => \N__29764\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__29770\,
            I => \N__29761\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__29767\,
            I => \N__29758\
        );

    \I__5341\ : Span4Mux_h
    port map (
            O => \N__29764\,
            I => \N__29755\
        );

    \I__5340\ : Span4Mux_h
    port map (
            O => \N__29761\,
            I => \N__29752\
        );

    \I__5339\ : Odrv12
    port map (
            O => \N__29758\,
            I => \nx.n2909\
        );

    \I__5338\ : Odrv4
    port map (
            O => \N__29755\,
            I => \nx.n2909\
        );

    \I__5337\ : Odrv4
    port map (
            O => \N__29752\,
            I => \nx.n2909\
        );

    \I__5336\ : InMux
    port map (
            O => \N__29745\,
            I => \N__29742\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__29742\,
            I => \nx.n2868\
        );

    \I__5334\ : InMux
    port map (
            O => \N__29739\,
            I => \N__29735\
        );

    \I__5333\ : CascadeMux
    port map (
            O => \N__29738\,
            I => \N__29732\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__29735\,
            I => \N__29729\
        );

    \I__5331\ : InMux
    port map (
            O => \N__29732\,
            I => \N__29726\
        );

    \I__5330\ : Span4Mux_v
    port map (
            O => \N__29729\,
            I => \N__29723\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__29726\,
            I => \N__29720\
        );

    \I__5328\ : Odrv4
    port map (
            O => \N__29723\,
            I => \nx.n2801\
        );

    \I__5327\ : Odrv12
    port map (
            O => \N__29720\,
            I => \nx.n2801\
        );

    \I__5326\ : InMux
    port map (
            O => \N__29715\,
            I => \N__29711\
        );

    \I__5325\ : CascadeMux
    port map (
            O => \N__29714\,
            I => \N__29708\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__29711\,
            I => \N__29704\
        );

    \I__5323\ : InMux
    port map (
            O => \N__29708\,
            I => \N__29701\
        );

    \I__5322\ : InMux
    port map (
            O => \N__29707\,
            I => \N__29698\
        );

    \I__5321\ : Span4Mux_s3_h
    port map (
            O => \N__29704\,
            I => \N__29691\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__29701\,
            I => \N__29691\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__29698\,
            I => \N__29691\
        );

    \I__5318\ : Odrv4
    port map (
            O => \N__29691\,
            I => \nx.n2900\
        );

    \I__5317\ : InMux
    port map (
            O => \N__29688\,
            I => \N__29685\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__29685\,
            I => \nx.n2861\
        );

    \I__5315\ : InMux
    port map (
            O => \N__29682\,
            I => \N__29678\
        );

    \I__5314\ : CascadeMux
    port map (
            O => \N__29681\,
            I => \N__29675\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__29678\,
            I => \N__29672\
        );

    \I__5312\ : InMux
    port map (
            O => \N__29675\,
            I => \N__29669\
        );

    \I__5311\ : Span4Mux_v
    port map (
            O => \N__29672\,
            I => \N__29665\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__29669\,
            I => \N__29662\
        );

    \I__5309\ : InMux
    port map (
            O => \N__29668\,
            I => \N__29659\
        );

    \I__5308\ : Odrv4
    port map (
            O => \N__29665\,
            I => \nx.n2794\
        );

    \I__5307\ : Odrv12
    port map (
            O => \N__29662\,
            I => \nx.n2794\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__29659\,
            I => \nx.n2794\
        );

    \I__5305\ : InMux
    port map (
            O => \N__29652\,
            I => \N__29647\
        );

    \I__5304\ : CascadeMux
    port map (
            O => \N__29651\,
            I => \N__29644\
        );

    \I__5303\ : InMux
    port map (
            O => \N__29650\,
            I => \N__29641\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__29647\,
            I => \N__29638\
        );

    \I__5301\ : InMux
    port map (
            O => \N__29644\,
            I => \N__29635\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__29641\,
            I => \N__29632\
        );

    \I__5299\ : Span4Mux_v
    port map (
            O => \N__29638\,
            I => \N__29627\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__29635\,
            I => \N__29627\
        );

    \I__5297\ : Span4Mux_h
    port map (
            O => \N__29632\,
            I => \N__29624\
        );

    \I__5296\ : Odrv4
    port map (
            O => \N__29627\,
            I => \nx.n2893\
        );

    \I__5295\ : Odrv4
    port map (
            O => \N__29624\,
            I => \nx.n2893\
        );

    \I__5294\ : InMux
    port map (
            O => \N__29619\,
            I => \N__29614\
        );

    \I__5293\ : InMux
    port map (
            O => \N__29618\,
            I => \N__29611\
        );

    \I__5292\ : InMux
    port map (
            O => \N__29617\,
            I => \N__29608\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__29614\,
            I => \N__29601\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__29611\,
            I => \N__29601\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__29608\,
            I => \N__29601\
        );

    \I__5288\ : Span4Mux_v
    port map (
            O => \N__29601\,
            I => \N__29598\
        );

    \I__5287\ : Odrv4
    port map (
            O => \N__29598\,
            I => \nx.n2788\
        );

    \I__5286\ : InMux
    port map (
            O => \N__29595\,
            I => \N__29592\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__29592\,
            I => \nx.n2855\
        );

    \I__5284\ : InMux
    port map (
            O => \N__29589\,
            I => \N__29586\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__29586\,
            I => \N__29582\
        );

    \I__5282\ : InMux
    port map (
            O => \N__29585\,
            I => \N__29579\
        );

    \I__5281\ : Span4Mux_v
    port map (
            O => \N__29582\,
            I => \N__29574\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__29579\,
            I => \N__29574\
        );

    \I__5279\ : Odrv4
    port map (
            O => \N__29574\,
            I => \nx.n2887\
        );

    \I__5278\ : InMux
    port map (
            O => \N__29571\,
            I => \N__29567\
        );

    \I__5277\ : CascadeMux
    port map (
            O => \N__29570\,
            I => \N__29564\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__29567\,
            I => \N__29560\
        );

    \I__5275\ : InMux
    port map (
            O => \N__29564\,
            I => \N__29557\
        );

    \I__5274\ : InMux
    port map (
            O => \N__29563\,
            I => \N__29554\
        );

    \I__5273\ : Odrv4
    port map (
            O => \N__29560\,
            I => \nx.n2890\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__29557\,
            I => \nx.n2890\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__29554\,
            I => \nx.n2890\
        );

    \I__5270\ : CascadeMux
    port map (
            O => \N__29547\,
            I => \N__29544\
        );

    \I__5269\ : InMux
    port map (
            O => \N__29544\,
            I => \N__29541\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__29541\,
            I => \nx.n2761\
        );

    \I__5267\ : InMux
    port map (
            O => \N__29538\,
            I => \N__29535\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__29535\,
            I => \nx.n2860\
        );

    \I__5265\ : CascadeMux
    port map (
            O => \N__29532\,
            I => \nx.n2793_cascade_\
        );

    \I__5264\ : CascadeMux
    port map (
            O => \N__29529\,
            I => \N__29525\
        );

    \I__5263\ : InMux
    port map (
            O => \N__29528\,
            I => \N__29522\
        );

    \I__5262\ : InMux
    port map (
            O => \N__29525\,
            I => \N__29519\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__29522\,
            I => \N__29515\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__29519\,
            I => \N__29512\
        );

    \I__5259\ : InMux
    port map (
            O => \N__29518\,
            I => \N__29509\
        );

    \I__5258\ : Span4Mux_h
    port map (
            O => \N__29515\,
            I => \N__29506\
        );

    \I__5257\ : Span4Mux_v
    port map (
            O => \N__29512\,
            I => \N__29503\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__29509\,
            I => \N__29500\
        );

    \I__5255\ : Odrv4
    port map (
            O => \N__29506\,
            I => \nx.n2892\
        );

    \I__5254\ : Odrv4
    port map (
            O => \N__29503\,
            I => \nx.n2892\
        );

    \I__5253\ : Odrv4
    port map (
            O => \N__29500\,
            I => \nx.n2892\
        );

    \I__5252\ : InMux
    port map (
            O => \N__29493\,
            I => \N__29490\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__29490\,
            I => \nx.n2758\
        );

    \I__5250\ : InMux
    port map (
            O => \N__29487\,
            I => \N__29484\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__29484\,
            I => \nx.n2760\
        );

    \I__5248\ : InMux
    port map (
            O => \N__29481\,
            I => \N__29478\
        );

    \I__5247\ : LocalMux
    port map (
            O => \N__29478\,
            I => \nx.n2873\
        );

    \I__5246\ : InMux
    port map (
            O => \N__29475\,
            I => \N__29471\
        );

    \I__5245\ : CascadeMux
    port map (
            O => \N__29474\,
            I => \N__29467\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__29471\,
            I => \N__29464\
        );

    \I__5243\ : InMux
    port map (
            O => \N__29470\,
            I => \N__29461\
        );

    \I__5242\ : InMux
    port map (
            O => \N__29467\,
            I => \N__29458\
        );

    \I__5241\ : Odrv4
    port map (
            O => \N__29464\,
            I => \nx.n2806\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__29461\,
            I => \nx.n2806\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__29458\,
            I => \nx.n2806\
        );

    \I__5238\ : InMux
    port map (
            O => \N__29451\,
            I => \N__29447\
        );

    \I__5237\ : InMux
    port map (
            O => \N__29450\,
            I => \N__29444\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__29447\,
            I => \N__29438\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__29444\,
            I => \N__29438\
        );

    \I__5234\ : InMux
    port map (
            O => \N__29443\,
            I => \N__29435\
        );

    \I__5233\ : Span4Mux_v
    port map (
            O => \N__29438\,
            I => \N__29430\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__29435\,
            I => \N__29430\
        );

    \I__5231\ : Odrv4
    port map (
            O => \N__29430\,
            I => \nx.n2905\
        );

    \I__5230\ : CascadeMux
    port map (
            O => \N__29427\,
            I => \N__29424\
        );

    \I__5229\ : InMux
    port map (
            O => \N__29424\,
            I => \N__29420\
        );

    \I__5228\ : InMux
    port map (
            O => \N__29423\,
            I => \N__29417\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__29420\,
            I => \nx.n2793\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__29417\,
            I => \nx.n2793\
        );

    \I__5225\ : CascadeMux
    port map (
            O => \N__29412\,
            I => \N__29409\
        );

    \I__5224\ : InMux
    port map (
            O => \N__29409\,
            I => \N__29405\
        );

    \I__5223\ : InMux
    port map (
            O => \N__29408\,
            I => \N__29402\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__29405\,
            I => \nx.n2791\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__29402\,
            I => \nx.n2791\
        );

    \I__5220\ : InMux
    port map (
            O => \N__29397\,
            I => \N__29392\
        );

    \I__5219\ : CascadeMux
    port map (
            O => \N__29396\,
            I => \N__29389\
        );

    \I__5218\ : CascadeMux
    port map (
            O => \N__29395\,
            I => \N__29386\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__29392\,
            I => \N__29383\
        );

    \I__5216\ : InMux
    port map (
            O => \N__29389\,
            I => \N__29380\
        );

    \I__5215\ : InMux
    port map (
            O => \N__29386\,
            I => \N__29377\
        );

    \I__5214\ : Odrv4
    port map (
            O => \N__29383\,
            I => \nx.n2792\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__29380\,
            I => \nx.n2792\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__29377\,
            I => \nx.n2792\
        );

    \I__5211\ : InMux
    port map (
            O => \N__29370\,
            I => \N__29366\
        );

    \I__5210\ : InMux
    port map (
            O => \N__29369\,
            I => \N__29363\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__29366\,
            I => \N__29358\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__29363\,
            I => \N__29358\
        );

    \I__5207\ : Odrv4
    port map (
            O => \N__29358\,
            I => \nx.n2786\
        );

    \I__5206\ : CascadeMux
    port map (
            O => \N__29355\,
            I => \nx.n38_adj_625_cascade_\
        );

    \I__5205\ : InMux
    port map (
            O => \N__29352\,
            I => \N__29349\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__29349\,
            I => \N__29346\
        );

    \I__5203\ : Span4Mux_v
    port map (
            O => \N__29346\,
            I => \N__29343\
        );

    \I__5202\ : Odrv4
    port map (
            O => \N__29343\,
            I => \nx.n42_adj_635\
        );

    \I__5201\ : InMux
    port map (
            O => \N__29340\,
            I => \N__29337\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__29337\,
            I => \N__29334\
        );

    \I__5199\ : Odrv4
    port map (
            O => \N__29334\,
            I => \nx.n41_adj_643\
        );

    \I__5198\ : CascadeMux
    port map (
            O => \N__29331\,
            I => \nx.n43_cascade_\
        );

    \I__5197\ : InMux
    port map (
            O => \N__29328\,
            I => \nx.n10806\
        );

    \I__5196\ : InMux
    port map (
            O => \N__29325\,
            I => \N__29322\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__29322\,
            I => \N__29319\
        );

    \I__5194\ : Odrv4
    port map (
            O => \N__29319\,
            I => \nx.n2759\
        );

    \I__5193\ : InMux
    port map (
            O => \N__29316\,
            I => \nx.n10807\
        );

    \I__5192\ : InMux
    port map (
            O => \N__29313\,
            I => \nx.n10808\
        );

    \I__5191\ : InMux
    port map (
            O => \N__29310\,
            I => \N__29307\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__29307\,
            I => \N__29304\
        );

    \I__5189\ : Odrv4
    port map (
            O => \N__29304\,
            I => \nx.n2757\
        );

    \I__5188\ : InMux
    port map (
            O => \N__29301\,
            I => \nx.n10809\
        );

    \I__5187\ : InMux
    port map (
            O => \N__29298\,
            I => \N__29295\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__29295\,
            I => \nx.n2756\
        );

    \I__5185\ : InMux
    port map (
            O => \N__29292\,
            I => \nx.n10810\
        );

    \I__5184\ : InMux
    port map (
            O => \N__29289\,
            I => \nx.n10811\
        );

    \I__5183\ : InMux
    port map (
            O => \N__29286\,
            I => \nx.n10812\
        );

    \I__5182\ : InMux
    port map (
            O => \N__29283\,
            I => \N__29280\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__29280\,
            I => \N__29277\
        );

    \I__5180\ : Span4Mux_v
    port map (
            O => \N__29277\,
            I => \N__29273\
        );

    \I__5179\ : InMux
    port map (
            O => \N__29276\,
            I => \N__29270\
        );

    \I__5178\ : Span4Mux_v
    port map (
            O => \N__29273\,
            I => \N__29267\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__29270\,
            I => neo_pixel_transmitter_t0_22
        );

    \I__5176\ : Odrv4
    port map (
            O => \N__29267\,
            I => neo_pixel_transmitter_t0_22
        );

    \I__5175\ : CascadeMux
    port map (
            O => \N__29262\,
            I => \N__29259\
        );

    \I__5174\ : InMux
    port map (
            O => \N__29259\,
            I => \N__29256\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__29256\,
            I => \N__29253\
        );

    \I__5172\ : Span4Mux_v
    port map (
            O => \N__29253\,
            I => \N__29250\
        );

    \I__5171\ : Span4Mux_h
    port map (
            O => \N__29250\,
            I => \N__29247\
        );

    \I__5170\ : Odrv4
    port map (
            O => \N__29247\,
            I => \nx.n11\
        );

    \I__5169\ : InMux
    port map (
            O => \N__29244\,
            I => \N__29241\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__29241\,
            I => \N__29238\
        );

    \I__5167\ : Odrv4
    port map (
            O => \N__29238\,
            I => \nx.n2768\
        );

    \I__5166\ : InMux
    port map (
            O => \N__29235\,
            I => \nx.n10798\
        );

    \I__5165\ : CascadeMux
    port map (
            O => \N__29232\,
            I => \N__29228\
        );

    \I__5164\ : CascadeMux
    port map (
            O => \N__29231\,
            I => \N__29225\
        );

    \I__5163\ : InMux
    port map (
            O => \N__29228\,
            I => \N__29222\
        );

    \I__5162\ : InMux
    port map (
            O => \N__29225\,
            I => \N__29219\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__29222\,
            I => \N__29214\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__29219\,
            I => \N__29214\
        );

    \I__5159\ : Odrv4
    port map (
            O => \N__29214\,
            I => \nx.n2700\
        );

    \I__5158\ : InMux
    port map (
            O => \N__29211\,
            I => \N__29208\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__29208\,
            I => \nx.n2767\
        );

    \I__5156\ : InMux
    port map (
            O => \N__29205\,
            I => \nx.n10799\
        );

    \I__5155\ : InMux
    port map (
            O => \N__29202\,
            I => \N__29199\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__29199\,
            I => \nx.n2766\
        );

    \I__5153\ : InMux
    port map (
            O => \N__29196\,
            I => \nx.n10800\
        );

    \I__5152\ : InMux
    port map (
            O => \N__29193\,
            I => \N__29190\
        );

    \I__5151\ : LocalMux
    port map (
            O => \N__29190\,
            I => \nx.n2765\
        );

    \I__5150\ : InMux
    port map (
            O => \N__29187\,
            I => \nx.n10801\
        );

    \I__5149\ : CascadeMux
    port map (
            O => \N__29184\,
            I => \N__29181\
        );

    \I__5148\ : InMux
    port map (
            O => \N__29181\,
            I => \N__29178\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__29178\,
            I => \nx.n2764\
        );

    \I__5146\ : InMux
    port map (
            O => \N__29175\,
            I => \nx.n10802\
        );

    \I__5145\ : CascadeMux
    port map (
            O => \N__29172\,
            I => \N__29168\
        );

    \I__5144\ : InMux
    port map (
            O => \N__29171\,
            I => \N__29164\
        );

    \I__5143\ : InMux
    port map (
            O => \N__29168\,
            I => \N__29161\
        );

    \I__5142\ : InMux
    port map (
            O => \N__29167\,
            I => \N__29158\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__29164\,
            I => \N__29153\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__29161\,
            I => \N__29153\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__29158\,
            I => \N__29150\
        );

    \I__5138\ : Span4Mux_h
    port map (
            O => \N__29153\,
            I => \N__29147\
        );

    \I__5137\ : Odrv12
    port map (
            O => \N__29150\,
            I => \nx.n2696\
        );

    \I__5136\ : Odrv4
    port map (
            O => \N__29147\,
            I => \nx.n2696\
        );

    \I__5135\ : CascadeMux
    port map (
            O => \N__29142\,
            I => \N__29139\
        );

    \I__5134\ : InMux
    port map (
            O => \N__29139\,
            I => \N__29136\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__29136\,
            I => \nx.n2763\
        );

    \I__5132\ : InMux
    port map (
            O => \N__29133\,
            I => \nx.n10803\
        );

    \I__5131\ : InMux
    port map (
            O => \N__29130\,
            I => \N__29127\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__29127\,
            I => \nx.n2762\
        );

    \I__5129\ : InMux
    port map (
            O => \N__29124\,
            I => \nx.n10804\
        );

    \I__5128\ : InMux
    port map (
            O => \N__29121\,
            I => \bfn_7_21_0_\
        );

    \I__5127\ : CascadeMux
    port map (
            O => \N__29118\,
            I => \N__29115\
        );

    \I__5126\ : InMux
    port map (
            O => \N__29115\,
            I => \N__29112\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__29112\,
            I => \nx.n2776\
        );

    \I__5124\ : InMux
    port map (
            O => \N__29109\,
            I => \nx.n10790\
        );

    \I__5123\ : CascadeMux
    port map (
            O => \N__29106\,
            I => \N__29102\
        );

    \I__5122\ : CascadeMux
    port map (
            O => \N__29105\,
            I => \N__29098\
        );

    \I__5121\ : InMux
    port map (
            O => \N__29102\,
            I => \N__29095\
        );

    \I__5120\ : InMux
    port map (
            O => \N__29101\,
            I => \N__29092\
        );

    \I__5119\ : InMux
    port map (
            O => \N__29098\,
            I => \N__29089\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__29095\,
            I => \nx.n2708\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__29092\,
            I => \nx.n2708\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__29089\,
            I => \nx.n2708\
        );

    \I__5115\ : InMux
    port map (
            O => \N__29082\,
            I => \N__29079\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__29079\,
            I => \nx.n2775\
        );

    \I__5113\ : InMux
    port map (
            O => \N__29076\,
            I => \nx.n10791\
        );

    \I__5112\ : CascadeMux
    port map (
            O => \N__29073\,
            I => \N__29070\
        );

    \I__5111\ : InMux
    port map (
            O => \N__29070\,
            I => \N__29065\
        );

    \I__5110\ : CascadeMux
    port map (
            O => \N__29069\,
            I => \N__29062\
        );

    \I__5109\ : CascadeMux
    port map (
            O => \N__29068\,
            I => \N__29059\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__29065\,
            I => \N__29056\
        );

    \I__5107\ : InMux
    port map (
            O => \N__29062\,
            I => \N__29053\
        );

    \I__5106\ : InMux
    port map (
            O => \N__29059\,
            I => \N__29050\
        );

    \I__5105\ : Odrv4
    port map (
            O => \N__29056\,
            I => \nx.n2707\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__29053\,
            I => \nx.n2707\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__29050\,
            I => \nx.n2707\
        );

    \I__5102\ : InMux
    port map (
            O => \N__29043\,
            I => \N__29040\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__29040\,
            I => \nx.n2774\
        );

    \I__5100\ : InMux
    port map (
            O => \N__29037\,
            I => \nx.n10792\
        );

    \I__5099\ : CascadeMux
    port map (
            O => \N__29034\,
            I => \N__29029\
        );

    \I__5098\ : InMux
    port map (
            O => \N__29033\,
            I => \N__29026\
        );

    \I__5097\ : InMux
    port map (
            O => \N__29032\,
            I => \N__29023\
        );

    \I__5096\ : InMux
    port map (
            O => \N__29029\,
            I => \N__29020\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__29026\,
            I => \nx.n2706\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__29023\,
            I => \nx.n2706\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__29020\,
            I => \nx.n2706\
        );

    \I__5092\ : CascadeMux
    port map (
            O => \N__29013\,
            I => \N__29010\
        );

    \I__5091\ : InMux
    port map (
            O => \N__29010\,
            I => \N__29007\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__29007\,
            I => \N__29004\
        );

    \I__5089\ : Odrv4
    port map (
            O => \N__29004\,
            I => \nx.n2773\
        );

    \I__5088\ : InMux
    port map (
            O => \N__29001\,
            I => \nx.n10793\
        );

    \I__5087\ : InMux
    port map (
            O => \N__28998\,
            I => \nx.n10794\
        );

    \I__5086\ : InMux
    port map (
            O => \N__28995\,
            I => \N__28992\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__28992\,
            I => \nx.n2771\
        );

    \I__5084\ : InMux
    port map (
            O => \N__28989\,
            I => \nx.n10795\
        );

    \I__5083\ : InMux
    port map (
            O => \N__28986\,
            I => \N__28983\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__28983\,
            I => \nx.n2770\
        );

    \I__5081\ : InMux
    port map (
            O => \N__28980\,
            I => \nx.n10796\
        );

    \I__5080\ : CascadeMux
    port map (
            O => \N__28977\,
            I => \N__28973\
        );

    \I__5079\ : CascadeMux
    port map (
            O => \N__28976\,
            I => \N__28970\
        );

    \I__5078\ : InMux
    port map (
            O => \N__28973\,
            I => \N__28966\
        );

    \I__5077\ : InMux
    port map (
            O => \N__28970\,
            I => \N__28961\
        );

    \I__5076\ : InMux
    port map (
            O => \N__28969\,
            I => \N__28961\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__28966\,
            I => \N__28958\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__28961\,
            I => \nx.n2702\
        );

    \I__5073\ : Odrv12
    port map (
            O => \N__28958\,
            I => \nx.n2702\
        );

    \I__5072\ : InMux
    port map (
            O => \N__28953\,
            I => \N__28950\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__28950\,
            I => \N__28947\
        );

    \I__5070\ : Odrv4
    port map (
            O => \N__28947\,
            I => \nx.n2769\
        );

    \I__5069\ : InMux
    port map (
            O => \N__28944\,
            I => \bfn_7_20_0_\
        );

    \I__5068\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28938\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__28938\,
            I => \N__28934\
        );

    \I__5066\ : InMux
    port map (
            O => \N__28937\,
            I => \N__28931\
        );

    \I__5065\ : Span4Mux_s1_v
    port map (
            O => \N__28934\,
            I => \N__28926\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__28931\,
            I => \N__28926\
        );

    \I__5063\ : Span4Mux_h
    port map (
            O => \N__28926\,
            I => \N__28923\
        );

    \I__5062\ : Odrv4
    port map (
            O => \N__28923\,
            I => \nx.n1499\
        );

    \I__5061\ : InMux
    port map (
            O => \N__28920\,
            I => \nx.n10602\
        );

    \I__5060\ : InMux
    port map (
            O => \N__28917\,
            I => \N__28912\
        );

    \I__5059\ : InMux
    port map (
            O => \N__28916\,
            I => \N__28909\
        );

    \I__5058\ : InMux
    port map (
            O => \N__28915\,
            I => \N__28906\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__28912\,
            I => \N__28901\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__28909\,
            I => \N__28901\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__28906\,
            I => \N__28898\
        );

    \I__5054\ : Span4Mux_v
    port map (
            O => \N__28901\,
            I => \N__28894\
        );

    \I__5053\ : Span4Mux_h
    port map (
            O => \N__28898\,
            I => \N__28891\
        );

    \I__5052\ : InMux
    port map (
            O => \N__28897\,
            I => \N__28888\
        );

    \I__5051\ : Span4Mux_h
    port map (
            O => \N__28894\,
            I => \N__28885\
        );

    \I__5050\ : Odrv4
    port map (
            O => \N__28891\,
            I => neopxl_color_13
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__28888\,
            I => neopxl_color_13
        );

    \I__5048\ : Odrv4
    port map (
            O => \N__28885\,
            I => neopxl_color_13
        );

    \I__5047\ : InMux
    port map (
            O => \N__28878\,
            I => \N__28870\
        );

    \I__5046\ : InMux
    port map (
            O => \N__28877\,
            I => \N__28867\
        );

    \I__5045\ : InMux
    port map (
            O => \N__28876\,
            I => \N__28859\
        );

    \I__5044\ : CascadeMux
    port map (
            O => \N__28875\,
            I => \N__28852\
        );

    \I__5043\ : InMux
    port map (
            O => \N__28874\,
            I => \N__28847\
        );

    \I__5042\ : CascadeMux
    port map (
            O => \N__28873\,
            I => \N__28844\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__28870\,
            I => \N__28828\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__28867\,
            I => \N__28828\
        );

    \I__5039\ : InMux
    port map (
            O => \N__28866\,
            I => \N__28825\
        );

    \I__5038\ : InMux
    port map (
            O => \N__28865\,
            I => \N__28822\
        );

    \I__5037\ : InMux
    port map (
            O => \N__28864\,
            I => \N__28815\
        );

    \I__5036\ : InMux
    port map (
            O => \N__28863\,
            I => \N__28815\
        );

    \I__5035\ : InMux
    port map (
            O => \N__28862\,
            I => \N__28815\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__28859\,
            I => \N__28812\
        );

    \I__5033\ : InMux
    port map (
            O => \N__28858\,
            I => \N__28807\
        );

    \I__5032\ : InMux
    port map (
            O => \N__28857\,
            I => \N__28807\
        );

    \I__5031\ : InMux
    port map (
            O => \N__28856\,
            I => \N__28802\
        );

    \I__5030\ : InMux
    port map (
            O => \N__28855\,
            I => \N__28802\
        );

    \I__5029\ : InMux
    port map (
            O => \N__28852\,
            I => \N__28797\
        );

    \I__5028\ : InMux
    port map (
            O => \N__28851\,
            I => \N__28797\
        );

    \I__5027\ : InMux
    port map (
            O => \N__28850\,
            I => \N__28794\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__28847\,
            I => \N__28791\
        );

    \I__5025\ : InMux
    port map (
            O => \N__28844\,
            I => \N__28786\
        );

    \I__5024\ : InMux
    port map (
            O => \N__28843\,
            I => \N__28786\
        );

    \I__5023\ : InMux
    port map (
            O => \N__28842\,
            I => \N__28783\
        );

    \I__5022\ : InMux
    port map (
            O => \N__28841\,
            I => \N__28778\
        );

    \I__5021\ : InMux
    port map (
            O => \N__28840\,
            I => \N__28778\
        );

    \I__5020\ : InMux
    port map (
            O => \N__28839\,
            I => \N__28769\
        );

    \I__5019\ : InMux
    port map (
            O => \N__28838\,
            I => \N__28769\
        );

    \I__5018\ : InMux
    port map (
            O => \N__28837\,
            I => \N__28764\
        );

    \I__5017\ : InMux
    port map (
            O => \N__28836\,
            I => \N__28764\
        );

    \I__5016\ : InMux
    port map (
            O => \N__28835\,
            I => \N__28757\
        );

    \I__5015\ : InMux
    port map (
            O => \N__28834\,
            I => \N__28757\
        );

    \I__5014\ : InMux
    port map (
            O => \N__28833\,
            I => \N__28757\
        );

    \I__5013\ : Span4Mux_v
    port map (
            O => \N__28828\,
            I => \N__28750\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__28825\,
            I => \N__28750\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__28822\,
            I => \N__28750\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__28815\,
            I => \N__28745\
        );

    \I__5009\ : Span4Mux_h
    port map (
            O => \N__28812\,
            I => \N__28745\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__28807\,
            I => \N__28742\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__28802\,
            I => \N__28735\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__28797\,
            I => \N__28735\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__28794\,
            I => \N__28735\
        );

    \I__5004\ : Span4Mux_v
    port map (
            O => \N__28791\,
            I => \N__28732\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__28786\,
            I => \N__28725\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__28783\,
            I => \N__28725\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__28778\,
            I => \N__28725\
        );

    \I__5000\ : InMux
    port map (
            O => \N__28777\,
            I => \N__28722\
        );

    \I__4999\ : InMux
    port map (
            O => \N__28776\,
            I => \N__28717\
        );

    \I__4998\ : InMux
    port map (
            O => \N__28775\,
            I => \N__28717\
        );

    \I__4997\ : InMux
    port map (
            O => \N__28774\,
            I => \N__28714\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__28769\,
            I => \N__28709\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__28764\,
            I => \N__28709\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__28757\,
            I => \N__28704\
        );

    \I__4993\ : Span4Mux_v
    port map (
            O => \N__28750\,
            I => \N__28704\
        );

    \I__4992\ : Span4Mux_v
    port map (
            O => \N__28745\,
            I => \N__28701\
        );

    \I__4991\ : Span4Mux_v
    port map (
            O => \N__28742\,
            I => \N__28692\
        );

    \I__4990\ : Span4Mux_v
    port map (
            O => \N__28735\,
            I => \N__28692\
        );

    \I__4989\ : Span4Mux_h
    port map (
            O => \N__28732\,
            I => \N__28692\
        );

    \I__4988\ : Span4Mux_v
    port map (
            O => \N__28725\,
            I => \N__28692\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__28722\,
            I => n11683
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__28717\,
            I => n11683
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__28714\,
            I => n11683
        );

    \I__4984\ : Odrv4
    port map (
            O => \N__28709\,
            I => n11683
        );

    \I__4983\ : Odrv4
    port map (
            O => \N__28704\,
            I => n11683
        );

    \I__4982\ : Odrv4
    port map (
            O => \N__28701\,
            I => n11683
        );

    \I__4981\ : Odrv4
    port map (
            O => \N__28692\,
            I => n11683
        );

    \I__4980\ : CascadeMux
    port map (
            O => \N__28677\,
            I => \N__28674\
        );

    \I__4979\ : InMux
    port map (
            O => \N__28674\,
            I => \N__28670\
        );

    \I__4978\ : InMux
    port map (
            O => \N__28673\,
            I => \N__28667\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__28670\,
            I => \N__28663\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__28667\,
            I => \N__28660\
        );

    \I__4975\ : InMux
    port map (
            O => \N__28666\,
            I => \N__28657\
        );

    \I__4974\ : Span4Mux_v
    port map (
            O => \N__28663\,
            I => \N__28654\
        );

    \I__4973\ : Odrv12
    port map (
            O => \N__28660\,
            I => timer_0
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__28657\,
            I => timer_0
        );

    \I__4971\ : Odrv4
    port map (
            O => \N__28654\,
            I => timer_0
        );

    \I__4970\ : InMux
    port map (
            O => \N__28647\,
            I => \N__28643\
        );

    \I__4969\ : InMux
    port map (
            O => \N__28646\,
            I => \N__28640\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__28643\,
            I => neo_pixel_transmitter_t0_0
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__28640\,
            I => neo_pixel_transmitter_t0_0
        );

    \I__4966\ : InMux
    port map (
            O => \N__28635\,
            I => \N__28632\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__28632\,
            I => \N__28629\
        );

    \I__4964\ : Span12Mux_v
    port map (
            O => \N__28629\,
            I => \N__28626\
        );

    \I__4963\ : Odrv12
    port map (
            O => \N__28626\,
            I => \nx.n33_adj_652\
        );

    \I__4962\ : IoInMux
    port map (
            O => \N__28623\,
            I => \N__28620\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__28620\,
            I => \N__28617\
        );

    \I__4960\ : Span12Mux_s4_v
    port map (
            O => \N__28617\,
            I => \N__28614\
        );

    \I__4959\ : Span12Mux_h
    port map (
            O => \N__28614\,
            I => \N__28609\
        );

    \I__4958\ : CascadeMux
    port map (
            O => \N__28613\,
            I => \N__28606\
        );

    \I__4957\ : InMux
    port map (
            O => \N__28612\,
            I => \N__28603\
        );

    \I__4956\ : Span12Mux_v
    port map (
            O => \N__28609\,
            I => \N__28600\
        );

    \I__4955\ : InMux
    port map (
            O => \N__28606\,
            I => \N__28597\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__28603\,
            I => \N__28594\
        );

    \I__4953\ : Odrv12
    port map (
            O => \N__28600\,
            I => pin_out_0
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__28597\,
            I => pin_out_0
        );

    \I__4951\ : Odrv4
    port map (
            O => \N__28594\,
            I => pin_out_0
        );

    \I__4950\ : IoInMux
    port map (
            O => \N__28587\,
            I => \N__28584\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__28584\,
            I => \N__28581\
        );

    \I__4948\ : IoSpan4Mux
    port map (
            O => \N__28581\,
            I => \N__28578\
        );

    \I__4947\ : Span4Mux_s3_v
    port map (
            O => \N__28578\,
            I => \N__28575\
        );

    \I__4946\ : Span4Mux_v
    port map (
            O => \N__28575\,
            I => \N__28572\
        );

    \I__4945\ : Span4Mux_v
    port map (
            O => \N__28572\,
            I => \N__28568\
        );

    \I__4944\ : CascadeMux
    port map (
            O => \N__28571\,
            I => \N__28565\
        );

    \I__4943\ : Span4Mux_v
    port map (
            O => \N__28568\,
            I => \N__28561\
        );

    \I__4942\ : InMux
    port map (
            O => \N__28565\,
            I => \N__28558\
        );

    \I__4941\ : InMux
    port map (
            O => \N__28564\,
            I => \N__28555\
        );

    \I__4940\ : Odrv4
    port map (
            O => \N__28561\,
            I => pin_out_1
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__28558\,
            I => pin_out_1
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__28555\,
            I => pin_out_1
        );

    \I__4937\ : InMux
    port map (
            O => \N__28548\,
            I => \N__28545\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__28545\,
            I => \N__28540\
        );

    \I__4935\ : InMux
    port map (
            O => \N__28544\,
            I => \N__28537\
        );

    \I__4934\ : InMux
    port map (
            O => \N__28543\,
            I => \N__28534\
        );

    \I__4933\ : Span4Mux_v
    port map (
            O => \N__28540\,
            I => \N__28530\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__28537\,
            I => \N__28527\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__28534\,
            I => \N__28524\
        );

    \I__4930\ : InMux
    port map (
            O => \N__28533\,
            I => \N__28520\
        );

    \I__4929\ : Span4Mux_v
    port map (
            O => \N__28530\,
            I => \N__28517\
        );

    \I__4928\ : Span4Mux_v
    port map (
            O => \N__28527\,
            I => \N__28512\
        );

    \I__4927\ : Span4Mux_v
    port map (
            O => \N__28524\,
            I => \N__28512\
        );

    \I__4926\ : InMux
    port map (
            O => \N__28523\,
            I => \N__28509\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__28520\,
            I => \N__28506\
        );

    \I__4924\ : Span4Mux_h
    port map (
            O => \N__28517\,
            I => \N__28503\
        );

    \I__4923\ : Span4Mux_v
    port map (
            O => \N__28512\,
            I => \N__28500\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__28509\,
            I => \nx.bit_ctr_8\
        );

    \I__4921\ : Odrv4
    port map (
            O => \N__28506\,
            I => \nx.bit_ctr_8\
        );

    \I__4920\ : Odrv4
    port map (
            O => \N__28503\,
            I => \nx.bit_ctr_8\
        );

    \I__4919\ : Odrv4
    port map (
            O => \N__28500\,
            I => \nx.bit_ctr_8\
        );

    \I__4918\ : InMux
    port map (
            O => \N__28491\,
            I => \N__28488\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__28488\,
            I => \N__28485\
        );

    \I__4916\ : Span4Mux_h
    port map (
            O => \N__28485\,
            I => \N__28482\
        );

    \I__4915\ : Odrv4
    port map (
            O => \N__28482\,
            I => \nx.n2777\
        );

    \I__4914\ : InMux
    port map (
            O => \N__28479\,
            I => \bfn_7_19_0_\
        );

    \I__4913\ : InMux
    port map (
            O => \N__28476\,
            I => \N__28469\
        );

    \I__4912\ : InMux
    port map (
            O => \N__28475\,
            I => \N__28469\
        );

    \I__4911\ : CascadeMux
    port map (
            O => \N__28474\,
            I => \N__28466\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__28469\,
            I => \N__28463\
        );

    \I__4909\ : InMux
    port map (
            O => \N__28466\,
            I => \N__28460\
        );

    \I__4908\ : Odrv4
    port map (
            O => \N__28463\,
            I => \nx.n1507\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__28460\,
            I => \nx.n1507\
        );

    \I__4906\ : CascadeMux
    port map (
            O => \N__28455\,
            I => \N__28452\
        );

    \I__4905\ : InMux
    port map (
            O => \N__28452\,
            I => \N__28449\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__28449\,
            I => \N__28446\
        );

    \I__4903\ : Odrv4
    port map (
            O => \N__28446\,
            I => \nx.n1574\
        );

    \I__4902\ : InMux
    port map (
            O => \N__28443\,
            I => \nx.n10594\
        );

    \I__4901\ : InMux
    port map (
            O => \N__28440\,
            I => \nx.n10595\
        );

    \I__4900\ : InMux
    port map (
            O => \N__28437\,
            I => \N__28434\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__28434\,
            I => \N__28429\
        );

    \I__4898\ : InMux
    port map (
            O => \N__28433\,
            I => \N__28426\
        );

    \I__4897\ : CascadeMux
    port map (
            O => \N__28432\,
            I => \N__28423\
        );

    \I__4896\ : Span4Mux_h
    port map (
            O => \N__28429\,
            I => \N__28418\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__28426\,
            I => \N__28418\
        );

    \I__4894\ : InMux
    port map (
            O => \N__28423\,
            I => \N__28415\
        );

    \I__4893\ : Odrv4
    port map (
            O => \N__28418\,
            I => \nx.n1505\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__28415\,
            I => \nx.n1505\
        );

    \I__4891\ : InMux
    port map (
            O => \N__28410\,
            I => \N__28407\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__28407\,
            I => \N__28404\
        );

    \I__4889\ : Odrv4
    port map (
            O => \N__28404\,
            I => \nx.n1572\
        );

    \I__4888\ : InMux
    port map (
            O => \N__28401\,
            I => \nx.n10596\
        );

    \I__4887\ : CascadeMux
    port map (
            O => \N__28398\,
            I => \N__28394\
        );

    \I__4886\ : InMux
    port map (
            O => \N__28397\,
            I => \N__28388\
        );

    \I__4885\ : InMux
    port map (
            O => \N__28394\,
            I => \N__28388\
        );

    \I__4884\ : CascadeMux
    port map (
            O => \N__28393\,
            I => \N__28385\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__28388\,
            I => \N__28382\
        );

    \I__4882\ : InMux
    port map (
            O => \N__28385\,
            I => \N__28379\
        );

    \I__4881\ : Span4Mux_h
    port map (
            O => \N__28382\,
            I => \N__28376\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__28379\,
            I => \nx.n1504\
        );

    \I__4879\ : Odrv4
    port map (
            O => \N__28376\,
            I => \nx.n1504\
        );

    \I__4878\ : InMux
    port map (
            O => \N__28371\,
            I => \N__28368\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__28368\,
            I => \N__28365\
        );

    \I__4876\ : Odrv4
    port map (
            O => \N__28365\,
            I => \nx.n1571\
        );

    \I__4875\ : InMux
    port map (
            O => \N__28362\,
            I => \nx.n10597\
        );

    \I__4874\ : InMux
    port map (
            O => \N__28359\,
            I => \nx.n10598\
        );

    \I__4873\ : CascadeMux
    port map (
            O => \N__28356\,
            I => \N__28352\
        );

    \I__4872\ : InMux
    port map (
            O => \N__28355\,
            I => \N__28348\
        );

    \I__4871\ : InMux
    port map (
            O => \N__28352\,
            I => \N__28345\
        );

    \I__4870\ : InMux
    port map (
            O => \N__28351\,
            I => \N__28342\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__28348\,
            I => \nx.n1502\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__28345\,
            I => \nx.n1502\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__28342\,
            I => \nx.n1502\
        );

    \I__4866\ : InMux
    port map (
            O => \N__28335\,
            I => \N__28332\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__28332\,
            I => \N__28329\
        );

    \I__4864\ : Odrv4
    port map (
            O => \N__28329\,
            I => \nx.n1569\
        );

    \I__4863\ : InMux
    port map (
            O => \N__28326\,
            I => \bfn_6_32_0_\
        );

    \I__4862\ : InMux
    port map (
            O => \N__28323\,
            I => \N__28319\
        );

    \I__4861\ : CascadeMux
    port map (
            O => \N__28322\,
            I => \N__28316\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__28319\,
            I => \N__28313\
        );

    \I__4859\ : InMux
    port map (
            O => \N__28316\,
            I => \N__28310\
        );

    \I__4858\ : Span4Mux_v
    port map (
            O => \N__28313\,
            I => \N__28305\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__28310\,
            I => \N__28305\
        );

    \I__4856\ : Odrv4
    port map (
            O => \N__28305\,
            I => \nx.n1501\
        );

    \I__4855\ : CascadeMux
    port map (
            O => \N__28302\,
            I => \N__28299\
        );

    \I__4854\ : InMux
    port map (
            O => \N__28299\,
            I => \N__28296\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__28296\,
            I => \N__28293\
        );

    \I__4852\ : Odrv4
    port map (
            O => \N__28293\,
            I => \nx.n1568\
        );

    \I__4851\ : InMux
    port map (
            O => \N__28290\,
            I => \nx.n10600\
        );

    \I__4850\ : InMux
    port map (
            O => \N__28287\,
            I => \N__28283\
        );

    \I__4849\ : CascadeMux
    port map (
            O => \N__28286\,
            I => \N__28280\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__28283\,
            I => \N__28276\
        );

    \I__4847\ : InMux
    port map (
            O => \N__28280\,
            I => \N__28273\
        );

    \I__4846\ : InMux
    port map (
            O => \N__28279\,
            I => \N__28270\
        );

    \I__4845\ : Odrv4
    port map (
            O => \N__28276\,
            I => \nx.n1500\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__28273\,
            I => \nx.n1500\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__28270\,
            I => \nx.n1500\
        );

    \I__4842\ : CascadeMux
    port map (
            O => \N__28263\,
            I => \N__28260\
        );

    \I__4841\ : InMux
    port map (
            O => \N__28260\,
            I => \N__28257\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__28257\,
            I => \N__28254\
        );

    \I__4839\ : Odrv4
    port map (
            O => \N__28254\,
            I => \nx.n1567\
        );

    \I__4838\ : InMux
    port map (
            O => \N__28251\,
            I => \nx.n10601\
        );

    \I__4837\ : InMux
    port map (
            O => \N__28248\,
            I => \N__28244\
        );

    \I__4836\ : CascadeMux
    port map (
            O => \N__28247\,
            I => \N__28240\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__28244\,
            I => \N__28237\
        );

    \I__4834\ : InMux
    port map (
            O => \N__28243\,
            I => \N__28234\
        );

    \I__4833\ : InMux
    port map (
            O => \N__28240\,
            I => \N__28231\
        );

    \I__4832\ : Odrv12
    port map (
            O => \N__28237\,
            I => \nx.n1409\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__28234\,
            I => \nx.n1409\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__28231\,
            I => \nx.n1409\
        );

    \I__4829\ : CascadeMux
    port map (
            O => \N__28224\,
            I => \N__28221\
        );

    \I__4828\ : InMux
    port map (
            O => \N__28221\,
            I => \N__28218\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__28218\,
            I => \N__28215\
        );

    \I__4826\ : Span4Mux_v
    port map (
            O => \N__28215\,
            I => \N__28212\
        );

    \I__4825\ : Odrv4
    port map (
            O => \N__28212\,
            I => \nx.n1476\
        );

    \I__4824\ : InMux
    port map (
            O => \N__28209\,
            I => \N__28204\
        );

    \I__4823\ : CascadeMux
    port map (
            O => \N__28208\,
            I => \N__28199\
        );

    \I__4822\ : CascadeMux
    port map (
            O => \N__28207\,
            I => \N__28196\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__28204\,
            I => \N__28192\
        );

    \I__4820\ : CascadeMux
    port map (
            O => \N__28203\,
            I => \N__28189\
        );

    \I__4819\ : CascadeMux
    port map (
            O => \N__28202\,
            I => \N__28183\
        );

    \I__4818\ : InMux
    port map (
            O => \N__28199\,
            I => \N__28175\
        );

    \I__4817\ : InMux
    port map (
            O => \N__28196\,
            I => \N__28175\
        );

    \I__4816\ : InMux
    port map (
            O => \N__28195\,
            I => \N__28175\
        );

    \I__4815\ : Span4Mux_h
    port map (
            O => \N__28192\,
            I => \N__28172\
        );

    \I__4814\ : InMux
    port map (
            O => \N__28189\,
            I => \N__28169\
        );

    \I__4813\ : InMux
    port map (
            O => \N__28188\,
            I => \N__28162\
        );

    \I__4812\ : InMux
    port map (
            O => \N__28187\,
            I => \N__28162\
        );

    \I__4811\ : InMux
    port map (
            O => \N__28186\,
            I => \N__28162\
        );

    \I__4810\ : InMux
    port map (
            O => \N__28183\,
            I => \N__28157\
        );

    \I__4809\ : InMux
    port map (
            O => \N__28182\,
            I => \N__28157\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__28175\,
            I => \nx.n1433\
        );

    \I__4807\ : Odrv4
    port map (
            O => \N__28172\,
            I => \nx.n1433\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__28169\,
            I => \nx.n1433\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__28162\,
            I => \nx.n1433\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__28157\,
            I => \nx.n1433\
        );

    \I__4803\ : CascadeMux
    port map (
            O => \N__28146\,
            I => \nx.n1508_cascade_\
        );

    \I__4802\ : InMux
    port map (
            O => \N__28143\,
            I => \N__28140\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__28140\,
            I => \nx.n16_adj_633\
        );

    \I__4800\ : CascadeMux
    port map (
            O => \N__28137\,
            I => \nx.n1599_cascade_\
        );

    \I__4799\ : InMux
    port map (
            O => \N__28134\,
            I => \bfn_6_31_0_\
        );

    \I__4798\ : InMux
    port map (
            O => \N__28131\,
            I => \nx.n10592\
        );

    \I__4797\ : CascadeMux
    port map (
            O => \N__28128\,
            I => \N__28124\
        );

    \I__4796\ : CascadeMux
    port map (
            O => \N__28127\,
            I => \N__28121\
        );

    \I__4795\ : InMux
    port map (
            O => \N__28124\,
            I => \N__28118\
        );

    \I__4794\ : InMux
    port map (
            O => \N__28121\,
            I => \N__28115\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__28118\,
            I => \nx.n1508\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__28115\,
            I => \nx.n1508\
        );

    \I__4791\ : InMux
    port map (
            O => \N__28110\,
            I => \N__28107\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__28107\,
            I => \N__28104\
        );

    \I__4789\ : Odrv4
    port map (
            O => \N__28104\,
            I => \nx.n1575\
        );

    \I__4788\ : InMux
    port map (
            O => \N__28101\,
            I => \nx.n10593\
        );

    \I__4787\ : InMux
    port map (
            O => \N__28098\,
            I => \N__28095\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__28095\,
            I => \N__28092\
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__28092\,
            I => \nx.n20_adj_634\
        );

    \I__4784\ : CascadeMux
    port map (
            O => \N__28089\,
            I => \nx.n1532_cascade_\
        );

    \I__4783\ : CascadeMux
    port map (
            O => \N__28086\,
            I => \nx.n1606_cascade_\
        );

    \I__4782\ : CascadeMux
    port map (
            O => \N__28083\,
            I => \nx.n22_adj_647_cascade_\
        );

    \I__4781\ : CascadeMux
    port map (
            O => \N__28080\,
            I => \nx.n1631_cascade_\
        );

    \I__4780\ : InMux
    port map (
            O => \N__28077\,
            I => \N__28074\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__28074\,
            I => \nx.n19_adj_602\
        );

    \I__4778\ : CascadeMux
    port map (
            O => \N__28071\,
            I => \N__28066\
        );

    \I__4777\ : CascadeMux
    port map (
            O => \N__28070\,
            I => \N__28063\
        );

    \I__4776\ : InMux
    port map (
            O => \N__28069\,
            I => \N__28060\
        );

    \I__4775\ : InMux
    port map (
            O => \N__28066\,
            I => \N__28057\
        );

    \I__4774\ : InMux
    port map (
            O => \N__28063\,
            I => \N__28053\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__28060\,
            I => \N__28049\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__28057\,
            I => \N__28046\
        );

    \I__4771\ : InMux
    port map (
            O => \N__28056\,
            I => \N__28043\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__28053\,
            I => \N__28040\
        );

    \I__4769\ : InMux
    port map (
            O => \N__28052\,
            I => \N__28037\
        );

    \I__4768\ : Span4Mux_v
    port map (
            O => \N__28049\,
            I => \N__28032\
        );

    \I__4767\ : Span4Mux_v
    port map (
            O => \N__28046\,
            I => \N__28032\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__28043\,
            I => \nx.bit_ctr_26\
        );

    \I__4765\ : Odrv4
    port map (
            O => \N__28040\,
            I => \nx.bit_ctr_26\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__28037\,
            I => \nx.bit_ctr_26\
        );

    \I__4763\ : Odrv4
    port map (
            O => \N__28032\,
            I => \nx.bit_ctr_26\
        );

    \I__4762\ : InMux
    port map (
            O => \N__28023\,
            I => \N__28020\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__28020\,
            I => \nx.n977\
        );

    \I__4760\ : InMux
    port map (
            O => \N__28017\,
            I => \bfn_6_28_0_\
        );

    \I__4759\ : CascadeMux
    port map (
            O => \N__28014\,
            I => \N__28010\
        );

    \I__4758\ : InMux
    port map (
            O => \N__28013\,
            I => \N__28007\
        );

    \I__4757\ : InMux
    port map (
            O => \N__28010\,
            I => \N__28004\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__28007\,
            I => \nx.n7082\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__28004\,
            I => \nx.n7082\
        );

    \I__4754\ : CascadeMux
    port map (
            O => \N__27999\,
            I => \N__27996\
        );

    \I__4753\ : InMux
    port map (
            O => \N__27996\,
            I => \N__27993\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__27993\,
            I => \nx.n976\
        );

    \I__4751\ : InMux
    port map (
            O => \N__27990\,
            I => \nx.n10474\
        );

    \I__4750\ : CascadeMux
    port map (
            O => \N__27987\,
            I => \N__27984\
        );

    \I__4749\ : InMux
    port map (
            O => \N__27984\,
            I => \N__27980\
        );

    \I__4748\ : InMux
    port map (
            O => \N__27983\,
            I => \N__27977\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__27980\,
            I => \nx.n7342\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__27977\,
            I => \nx.n7342\
        );

    \I__4745\ : CascadeMux
    port map (
            O => \N__27972\,
            I => \N__27968\
        );

    \I__4744\ : InMux
    port map (
            O => \N__27971\,
            I => \N__27963\
        );

    \I__4743\ : InMux
    port map (
            O => \N__27968\,
            I => \N__27963\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__27963\,
            I => \nx.n975\
        );

    \I__4741\ : InMux
    port map (
            O => \N__27960\,
            I => \nx.n10475\
        );

    \I__4740\ : CascadeMux
    port map (
            O => \N__27957\,
            I => \N__27953\
        );

    \I__4739\ : InMux
    port map (
            O => \N__27956\,
            I => \N__27950\
        );

    \I__4738\ : InMux
    port map (
            O => \N__27953\,
            I => \N__27947\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__27950\,
            I => \nx.n974\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__27947\,
            I => \nx.n974\
        );

    \I__4735\ : InMux
    port map (
            O => \N__27942\,
            I => \nx.n10476\
        );

    \I__4734\ : CascadeMux
    port map (
            O => \N__27939\,
            I => \N__27935\
        );

    \I__4733\ : CascadeMux
    port map (
            O => \N__27938\,
            I => \N__27932\
        );

    \I__4732\ : InMux
    port map (
            O => \N__27935\,
            I => \N__27928\
        );

    \I__4731\ : InMux
    port map (
            O => \N__27932\,
            I => \N__27925\
        );

    \I__4730\ : InMux
    port map (
            O => \N__27931\,
            I => \N__27922\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__27928\,
            I => \nx.n906\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__27925\,
            I => \nx.n906\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__27922\,
            I => \nx.n906\
        );

    \I__4726\ : InMux
    port map (
            O => \N__27915\,
            I => \N__27912\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__27912\,
            I => \nx.n973\
        );

    \I__4724\ : InMux
    port map (
            O => \N__27909\,
            I => \nx.n10477\
        );

    \I__4723\ : InMux
    port map (
            O => \N__27906\,
            I => \N__27902\
        );

    \I__4722\ : InMux
    port map (
            O => \N__27905\,
            I => \N__27899\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__27902\,
            I => \nx.n13064\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__27899\,
            I => \nx.n13064\
        );

    \I__4719\ : InMux
    port map (
            O => \N__27894\,
            I => \nx.n10478\
        );

    \I__4718\ : CascadeMux
    port map (
            O => \N__27891\,
            I => \N__27888\
        );

    \I__4717\ : InMux
    port map (
            O => \N__27888\,
            I => \N__27885\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__27885\,
            I => \N__27881\
        );

    \I__4715\ : InMux
    port map (
            O => \N__27884\,
            I => \N__27878\
        );

    \I__4714\ : Odrv4
    port map (
            O => \N__27881\,
            I => \nx.n4_adj_596\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__27878\,
            I => \nx.n4_adj_596\
        );

    \I__4712\ : InMux
    port map (
            O => \N__27873\,
            I => \N__27866\
        );

    \I__4711\ : InMux
    port map (
            O => \N__27872\,
            I => \N__27866\
        );

    \I__4710\ : InMux
    port map (
            O => \N__27871\,
            I => \N__27863\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__27866\,
            I => \N__27860\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__27863\,
            I => \nx.n5260\
        );

    \I__4707\ : Odrv4
    port map (
            O => \N__27860\,
            I => \nx.n5260\
        );

    \I__4706\ : CascadeMux
    port map (
            O => \N__27855\,
            I => \N__27850\
        );

    \I__4705\ : InMux
    port map (
            O => \N__27854\,
            I => \N__27845\
        );

    \I__4704\ : InMux
    port map (
            O => \N__27853\,
            I => \N__27845\
        );

    \I__4703\ : InMux
    port map (
            O => \N__27850\,
            I => \N__27842\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__27845\,
            I => \N__27838\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__27842\,
            I => \N__27835\
        );

    \I__4700\ : InMux
    port map (
            O => \N__27841\,
            I => \N__27832\
        );

    \I__4699\ : Odrv12
    port map (
            O => \N__27838\,
            I => \nx.n11559\
        );

    \I__4698\ : Odrv4
    port map (
            O => \N__27835\,
            I => \nx.n11559\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__27832\,
            I => \nx.n11559\
        );

    \I__4696\ : CascadeMux
    port map (
            O => \N__27825\,
            I => \N__27820\
        );

    \I__4695\ : CascadeMux
    port map (
            O => \N__27824\,
            I => \N__27817\
        );

    \I__4694\ : InMux
    port map (
            O => \N__27823\,
            I => \N__27812\
        );

    \I__4693\ : InMux
    port map (
            O => \N__27820\,
            I => \N__27803\
        );

    \I__4692\ : InMux
    port map (
            O => \N__27817\,
            I => \N__27803\
        );

    \I__4691\ : InMux
    port map (
            O => \N__27816\,
            I => \N__27803\
        );

    \I__4690\ : InMux
    port map (
            O => \N__27815\,
            I => \N__27803\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__27812\,
            I => \nx.n838\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__27803\,
            I => \nx.n838\
        );

    \I__4687\ : CascadeMux
    port map (
            O => \N__27798\,
            I => \N__27795\
        );

    \I__4686\ : InMux
    port map (
            O => \N__27795\,
            I => \N__27791\
        );

    \I__4685\ : InMux
    port map (
            O => \N__27794\,
            I => \N__27788\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__27791\,
            I => \nx.n11674\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__27788\,
            I => \nx.n11674\
        );

    \I__4682\ : CascadeMux
    port map (
            O => \N__27783\,
            I => \nx.n1829_cascade_\
        );

    \I__4681\ : CascadeMux
    port map (
            O => \N__27780\,
            I => \nx.n1906_cascade_\
        );

    \I__4680\ : CascadeMux
    port map (
            O => \N__27777\,
            I => \N__27774\
        );

    \I__4679\ : InMux
    port map (
            O => \N__27774\,
            I => \N__27771\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__27771\,
            I => \nx.n22_adj_605\
        );

    \I__4677\ : CascadeMux
    port map (
            O => \N__27768\,
            I => \N__27764\
        );

    \I__4676\ : CascadeMux
    port map (
            O => \N__27767\,
            I => \N__27761\
        );

    \I__4675\ : InMux
    port map (
            O => \N__27764\,
            I => \N__27758\
        );

    \I__4674\ : InMux
    port map (
            O => \N__27761\,
            I => \N__27755\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__27758\,
            I => \nx.n1006\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__27755\,
            I => \nx.n1006\
        );

    \I__4671\ : CascadeMux
    port map (
            O => \N__27750\,
            I => \nx.n1804_cascade_\
        );

    \I__4670\ : CascadeMux
    port map (
            O => \N__27747\,
            I => \nx.n19_cascade_\
        );

    \I__4669\ : InMux
    port map (
            O => \N__27744\,
            I => \N__27741\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__27741\,
            I => \nx.n26_adj_600\
        );

    \I__4667\ : InMux
    port map (
            O => \N__27738\,
            I => \N__27733\
        );

    \I__4666\ : InMux
    port map (
            O => \N__27737\,
            I => \N__27729\
        );

    \I__4665\ : CascadeMux
    port map (
            O => \N__27736\,
            I => \N__27725\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__27733\,
            I => \N__27720\
        );

    \I__4663\ : InMux
    port map (
            O => \N__27732\,
            I => \N__27717\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__27729\,
            I => \N__27714\
        );

    \I__4661\ : InMux
    port map (
            O => \N__27728\,
            I => \N__27711\
        );

    \I__4660\ : InMux
    port map (
            O => \N__27725\,
            I => \N__27704\
        );

    \I__4659\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27704\
        );

    \I__4658\ : InMux
    port map (
            O => \N__27723\,
            I => \N__27704\
        );

    \I__4657\ : Span4Mux_h
    port map (
            O => \N__27720\,
            I => \N__27701\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__27717\,
            I => \nx.bit_ctr_27\
        );

    \I__4655\ : Odrv4
    port map (
            O => \N__27714\,
            I => \nx.bit_ctr_27\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__27711\,
            I => \nx.bit_ctr_27\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__27704\,
            I => \nx.bit_ctr_27\
        );

    \I__4652\ : Odrv4
    port map (
            O => \N__27701\,
            I => \nx.bit_ctr_27\
        );

    \I__4651\ : CascadeMux
    port map (
            O => \N__27690\,
            I => \N__27686\
        );

    \I__4650\ : InMux
    port map (
            O => \N__27689\,
            I => \N__27683\
        );

    \I__4649\ : InMux
    port map (
            O => \N__27686\,
            I => \N__27679\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__27683\,
            I => \N__27675\
        );

    \I__4647\ : CascadeMux
    port map (
            O => \N__27682\,
            I => \N__27671\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__27679\,
            I => \N__27668\
        );

    \I__4645\ : InMux
    port map (
            O => \N__27678\,
            I => \N__27663\
        );

    \I__4644\ : Span4Mux_h
    port map (
            O => \N__27675\,
            I => \N__27660\
        );

    \I__4643\ : InMux
    port map (
            O => \N__27674\,
            I => \N__27655\
        );

    \I__4642\ : InMux
    port map (
            O => \N__27671\,
            I => \N__27655\
        );

    \I__4641\ : Span4Mux_v
    port map (
            O => \N__27668\,
            I => \N__27652\
        );

    \I__4640\ : InMux
    port map (
            O => \N__27667\,
            I => \N__27647\
        );

    \I__4639\ : InMux
    port map (
            O => \N__27666\,
            I => \N__27647\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__27663\,
            I => \nx.bit_ctr_28\
        );

    \I__4637\ : Odrv4
    port map (
            O => \N__27660\,
            I => \nx.bit_ctr_28\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__27655\,
            I => \nx.bit_ctr_28\
        );

    \I__4635\ : Odrv4
    port map (
            O => \N__27652\,
            I => \nx.bit_ctr_28\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__27647\,
            I => \nx.bit_ctr_28\
        );

    \I__4633\ : CascadeMux
    port map (
            O => \N__27636\,
            I => \N__27632\
        );

    \I__4632\ : InMux
    port map (
            O => \N__27635\,
            I => \N__27628\
        );

    \I__4631\ : InMux
    port map (
            O => \N__27632\,
            I => \N__27622\
        );

    \I__4630\ : InMux
    port map (
            O => \N__27631\,
            I => \N__27622\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__27628\,
            I => \N__27619\
        );

    \I__4628\ : InMux
    port map (
            O => \N__27627\,
            I => \N__27616\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__27622\,
            I => \nx.n739\
        );

    \I__4626\ : Odrv4
    port map (
            O => \N__27619\,
            I => \nx.n739\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__27616\,
            I => \nx.n739\
        );

    \I__4624\ : CascadeMux
    port map (
            O => \N__27609\,
            I => \nx.n28_adj_660_cascade_\
        );

    \I__4623\ : InMux
    port map (
            O => \N__27606\,
            I => \N__27603\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__27603\,
            I => \nx.n16\
        );

    \I__4621\ : CascadeMux
    port map (
            O => \N__27600\,
            I => \nx.n1928_cascade_\
        );

    \I__4620\ : CascadeMux
    port map (
            O => \N__27597\,
            I => \nx.n1908_cascade_\
        );

    \I__4619\ : InMux
    port map (
            O => \N__27594\,
            I => \N__27591\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__27591\,
            I => \nx.n24_adj_648\
        );

    \I__4617\ : InMux
    port map (
            O => \N__27588\,
            I => \N__27585\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__27585\,
            I => \nx.n1877\
        );

    \I__4615\ : InMux
    port map (
            O => \N__27582\,
            I => \bfn_6_24_0_\
        );

    \I__4614\ : InMux
    port map (
            O => \N__27579\,
            I => \N__27575\
        );

    \I__4613\ : CascadeMux
    port map (
            O => \N__27578\,
            I => \N__27572\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__27575\,
            I => \N__27569\
        );

    \I__4611\ : InMux
    port map (
            O => \N__27572\,
            I => \N__27566\
        );

    \I__4610\ : Span4Mux_v
    port map (
            O => \N__27569\,
            I => \N__27563\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__27566\,
            I => \nx.n2885\
        );

    \I__4608\ : Odrv4
    port map (
            O => \N__27563\,
            I => \nx.n2885\
        );

    \I__4607\ : InMux
    port map (
            O => \N__27558\,
            I => \N__27555\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__27555\,
            I => \nx.n2858\
        );

    \I__4605\ : CascadeMux
    port map (
            O => \N__27552\,
            I => \nx.n2791_cascade_\
        );

    \I__4604\ : InMux
    port map (
            O => \N__27549\,
            I => \N__27546\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__27546\,
            I => \nx.n2859\
        );

    \I__4602\ : InMux
    port map (
            O => \N__27543\,
            I => \N__27538\
        );

    \I__4601\ : InMux
    port map (
            O => \N__27542\,
            I => \N__27535\
        );

    \I__4600\ : CascadeMux
    port map (
            O => \N__27541\,
            I => \N__27532\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__27538\,
            I => \N__27529\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__27535\,
            I => \N__27526\
        );

    \I__4597\ : InMux
    port map (
            O => \N__27532\,
            I => \N__27523\
        );

    \I__4596\ : Span4Mux_h
    port map (
            O => \N__27529\,
            I => \N__27520\
        );

    \I__4595\ : Odrv4
    port map (
            O => \N__27526\,
            I => \nx.n2891\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__27523\,
            I => \nx.n2891\
        );

    \I__4593\ : Odrv4
    port map (
            O => \N__27520\,
            I => \nx.n2891\
        );

    \I__4592\ : InMux
    port map (
            O => \N__27513\,
            I => \N__27510\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__27510\,
            I => \nx.n2856\
        );

    \I__4590\ : CascadeMux
    port map (
            O => \N__27507\,
            I => \nx.n2789_cascade_\
        );

    \I__4589\ : InMux
    port map (
            O => \N__27504\,
            I => \N__27500\
        );

    \I__4588\ : InMux
    port map (
            O => \N__27503\,
            I => \N__27497\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__27500\,
            I => \N__27494\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__27497\,
            I => \N__27491\
        );

    \I__4585\ : Span4Mux_v
    port map (
            O => \N__27494\,
            I => \N__27488\
        );

    \I__4584\ : Span4Mux_v
    port map (
            O => \N__27491\,
            I => \N__27485\
        );

    \I__4583\ : Odrv4
    port map (
            O => \N__27488\,
            I => \nx.n2995\
        );

    \I__4582\ : Odrv4
    port map (
            O => \N__27485\,
            I => \nx.n2995\
        );

    \I__4581\ : CascadeMux
    port map (
            O => \N__27480\,
            I => \N__27477\
        );

    \I__4580\ : InMux
    port map (
            O => \N__27477\,
            I => \N__27474\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__27474\,
            I => \N__27471\
        );

    \I__4578\ : Span4Mux_h
    port map (
            O => \N__27471\,
            I => \N__27468\
        );

    \I__4577\ : Odrv4
    port map (
            O => \N__27468\,
            I => \nx.n3062\
        );

    \I__4576\ : CascadeMux
    port map (
            O => \N__27465\,
            I => \N__27460\
        );

    \I__4575\ : CascadeMux
    port map (
            O => \N__27464\,
            I => \N__27453\
        );

    \I__4574\ : InMux
    port map (
            O => \N__27463\,
            I => \N__27448\
        );

    \I__4573\ : InMux
    port map (
            O => \N__27460\,
            I => \N__27445\
        );

    \I__4572\ : InMux
    port map (
            O => \N__27459\,
            I => \N__27442\
        );

    \I__4571\ : InMux
    port map (
            O => \N__27458\,
            I => \N__27433\
        );

    \I__4570\ : InMux
    port map (
            O => \N__27457\,
            I => \N__27430\
        );

    \I__4569\ : InMux
    port map (
            O => \N__27456\,
            I => \N__27423\
        );

    \I__4568\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27423\
        );

    \I__4567\ : InMux
    port map (
            O => \N__27452\,
            I => \N__27423\
        );

    \I__4566\ : CascadeMux
    port map (
            O => \N__27451\,
            I => \N__27416\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__27448\,
            I => \N__27412\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__27445\,
            I => \N__27407\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__27442\,
            I => \N__27407\
        );

    \I__4562\ : InMux
    port map (
            O => \N__27441\,
            I => \N__27402\
        );

    \I__4561\ : InMux
    port map (
            O => \N__27440\,
            I => \N__27402\
        );

    \I__4560\ : CascadeMux
    port map (
            O => \N__27439\,
            I => \N__27396\
        );

    \I__4559\ : CascadeMux
    port map (
            O => \N__27438\,
            I => \N__27393\
        );

    \I__4558\ : CascadeMux
    port map (
            O => \N__27437\,
            I => \N__27390\
        );

    \I__4557\ : CascadeMux
    port map (
            O => \N__27436\,
            I => \N__27384\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__27433\,
            I => \N__27377\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__27430\,
            I => \N__27377\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__27423\,
            I => \N__27377\
        );

    \I__4553\ : InMux
    port map (
            O => \N__27422\,
            I => \N__27372\
        );

    \I__4552\ : InMux
    port map (
            O => \N__27421\,
            I => \N__27372\
        );

    \I__4551\ : InMux
    port map (
            O => \N__27420\,
            I => \N__27363\
        );

    \I__4550\ : InMux
    port map (
            O => \N__27419\,
            I => \N__27363\
        );

    \I__4549\ : InMux
    port map (
            O => \N__27416\,
            I => \N__27363\
        );

    \I__4548\ : InMux
    port map (
            O => \N__27415\,
            I => \N__27363\
        );

    \I__4547\ : Span4Mux_v
    port map (
            O => \N__27412\,
            I => \N__27360\
        );

    \I__4546\ : Span4Mux_v
    port map (
            O => \N__27407\,
            I => \N__27355\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__27402\,
            I => \N__27355\
        );

    \I__4544\ : InMux
    port map (
            O => \N__27401\,
            I => \N__27350\
        );

    \I__4543\ : InMux
    port map (
            O => \N__27400\,
            I => \N__27350\
        );

    \I__4542\ : InMux
    port map (
            O => \N__27399\,
            I => \N__27339\
        );

    \I__4541\ : InMux
    port map (
            O => \N__27396\,
            I => \N__27339\
        );

    \I__4540\ : InMux
    port map (
            O => \N__27393\,
            I => \N__27339\
        );

    \I__4539\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27339\
        );

    \I__4538\ : InMux
    port map (
            O => \N__27389\,
            I => \N__27339\
        );

    \I__4537\ : InMux
    port map (
            O => \N__27388\,
            I => \N__27332\
        );

    \I__4536\ : InMux
    port map (
            O => \N__27387\,
            I => \N__27332\
        );

    \I__4535\ : InMux
    port map (
            O => \N__27384\,
            I => \N__27332\
        );

    \I__4534\ : Span4Mux_h
    port map (
            O => \N__27377\,
            I => \N__27329\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__27372\,
            I => \nx.n3017\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__27363\,
            I => \nx.n3017\
        );

    \I__4531\ : Odrv4
    port map (
            O => \N__27360\,
            I => \nx.n3017\
        );

    \I__4530\ : Odrv4
    port map (
            O => \N__27355\,
            I => \nx.n3017\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__27350\,
            I => \nx.n3017\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__27339\,
            I => \nx.n3017\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__27332\,
            I => \nx.n3017\
        );

    \I__4526\ : Odrv4
    port map (
            O => \N__27329\,
            I => \nx.n3017\
        );

    \I__4525\ : InMux
    port map (
            O => \N__27312\,
            I => \N__27308\
        );

    \I__4524\ : InMux
    port map (
            O => \N__27311\,
            I => \N__27304\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__27308\,
            I => \N__27301\
        );

    \I__4522\ : CascadeMux
    port map (
            O => \N__27307\,
            I => \N__27298\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__27304\,
            I => \N__27293\
        );

    \I__4520\ : Span12Mux_s7_v
    port map (
            O => \N__27301\,
            I => \N__27293\
        );

    \I__4519\ : InMux
    port map (
            O => \N__27298\,
            I => \N__27290\
        );

    \I__4518\ : Odrv12
    port map (
            O => \N__27293\,
            I => \nx.n3094\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__27290\,
            I => \nx.n3094\
        );

    \I__4516\ : InMux
    port map (
            O => \N__27285\,
            I => \N__27281\
        );

    \I__4515\ : CascadeMux
    port map (
            O => \N__27284\,
            I => \N__27278\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__27281\,
            I => \N__27275\
        );

    \I__4513\ : InMux
    port map (
            O => \N__27278\,
            I => \N__27272\
        );

    \I__4512\ : Span4Mux_h
    port map (
            O => \N__27275\,
            I => \N__27266\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__27272\,
            I => \N__27266\
        );

    \I__4510\ : InMux
    port map (
            O => \N__27271\,
            I => \N__27263\
        );

    \I__4509\ : Odrv4
    port map (
            O => \N__27266\,
            I => \nx.n2795\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__27263\,
            I => \nx.n2795\
        );

    \I__4507\ : CascadeMux
    port map (
            O => \N__27258\,
            I => \N__27255\
        );

    \I__4506\ : InMux
    port map (
            O => \N__27255\,
            I => \N__27252\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__27252\,
            I => \N__27249\
        );

    \I__4504\ : Odrv4
    port map (
            O => \N__27249\,
            I => \nx.n2862\
        );

    \I__4503\ : InMux
    port map (
            O => \N__27246\,
            I => \nx.n10827\
        );

    \I__4502\ : InMux
    port map (
            O => \N__27243\,
            I => \bfn_6_23_0_\
        );

    \I__4501\ : InMux
    port map (
            O => \N__27240\,
            I => \nx.n10829\
        );

    \I__4500\ : InMux
    port map (
            O => \N__27237\,
            I => \nx.n10830\
        );

    \I__4499\ : InMux
    port map (
            O => \N__27234\,
            I => \nx.n10831\
        );

    \I__4498\ : InMux
    port map (
            O => \N__27231\,
            I => \nx.n10832\
        );

    \I__4497\ : InMux
    port map (
            O => \N__27228\,
            I => \nx.n10833\
        );

    \I__4496\ : InMux
    port map (
            O => \N__27225\,
            I => \nx.n10834\
        );

    \I__4495\ : InMux
    port map (
            O => \N__27222\,
            I => \nx.n10835\
        );

    \I__4494\ : InMux
    port map (
            O => \N__27219\,
            I => \nx.n10819\
        );

    \I__4493\ : CascadeMux
    port map (
            O => \N__27216\,
            I => \N__27212\
        );

    \I__4492\ : CascadeMux
    port map (
            O => \N__27215\,
            I => \N__27209\
        );

    \I__4491\ : InMux
    port map (
            O => \N__27212\,
            I => \N__27206\
        );

    \I__4490\ : InMux
    port map (
            O => \N__27209\,
            I => \N__27203\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__27206\,
            I => \N__27199\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__27203\,
            I => \N__27196\
        );

    \I__4487\ : InMux
    port map (
            O => \N__27202\,
            I => \N__27193\
        );

    \I__4486\ : Odrv4
    port map (
            O => \N__27199\,
            I => \nx.n2802\
        );

    \I__4485\ : Odrv12
    port map (
            O => \N__27196\,
            I => \nx.n2802\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__27193\,
            I => \nx.n2802\
        );

    \I__4483\ : InMux
    port map (
            O => \N__27186\,
            I => \N__27183\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__27183\,
            I => \nx.n2869\
        );

    \I__4481\ : InMux
    port map (
            O => \N__27180\,
            I => \bfn_6_22_0_\
        );

    \I__4480\ : InMux
    port map (
            O => \N__27177\,
            I => \nx.n10821\
        );

    \I__4479\ : CascadeMux
    port map (
            O => \N__27174\,
            I => \N__27170\
        );

    \I__4478\ : InMux
    port map (
            O => \N__27173\,
            I => \N__27167\
        );

    \I__4477\ : InMux
    port map (
            O => \N__27170\,
            I => \N__27164\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__27167\,
            I => \N__27160\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__27164\,
            I => \N__27157\
        );

    \I__4474\ : InMux
    port map (
            O => \N__27163\,
            I => \N__27154\
        );

    \I__4473\ : Odrv4
    port map (
            O => \N__27160\,
            I => \nx.n2800\
        );

    \I__4472\ : Odrv4
    port map (
            O => \N__27157\,
            I => \nx.n2800\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__27154\,
            I => \nx.n2800\
        );

    \I__4470\ : CascadeMux
    port map (
            O => \N__27147\,
            I => \N__27144\
        );

    \I__4469\ : InMux
    port map (
            O => \N__27144\,
            I => \N__27141\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__27141\,
            I => \N__27138\
        );

    \I__4467\ : Odrv4
    port map (
            O => \N__27138\,
            I => \nx.n2867\
        );

    \I__4466\ : InMux
    port map (
            O => \N__27135\,
            I => \nx.n10822\
        );

    \I__4465\ : CascadeMux
    port map (
            O => \N__27132\,
            I => \N__27128\
        );

    \I__4464\ : InMux
    port map (
            O => \N__27131\,
            I => \N__27125\
        );

    \I__4463\ : InMux
    port map (
            O => \N__27128\,
            I => \N__27122\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__27125\,
            I => \N__27116\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__27122\,
            I => \N__27116\
        );

    \I__4460\ : InMux
    port map (
            O => \N__27121\,
            I => \N__27113\
        );

    \I__4459\ : Odrv4
    port map (
            O => \N__27116\,
            I => \nx.n2799\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__27113\,
            I => \nx.n2799\
        );

    \I__4457\ : InMux
    port map (
            O => \N__27108\,
            I => \N__27105\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__27105\,
            I => \nx.n2866\
        );

    \I__4455\ : InMux
    port map (
            O => \N__27102\,
            I => \nx.n10823\
        );

    \I__4454\ : CascadeMux
    port map (
            O => \N__27099\,
            I => \N__27096\
        );

    \I__4453\ : InMux
    port map (
            O => \N__27096\,
            I => \N__27091\
        );

    \I__4452\ : InMux
    port map (
            O => \N__27095\,
            I => \N__27088\
        );

    \I__4451\ : InMux
    port map (
            O => \N__27094\,
            I => \N__27085\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__27091\,
            I => \N__27082\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__27088\,
            I => \N__27079\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__27085\,
            I => \nx.n2798\
        );

    \I__4447\ : Odrv4
    port map (
            O => \N__27082\,
            I => \nx.n2798\
        );

    \I__4446\ : Odrv4
    port map (
            O => \N__27079\,
            I => \nx.n2798\
        );

    \I__4445\ : InMux
    port map (
            O => \N__27072\,
            I => \N__27069\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__27069\,
            I => \N__27066\
        );

    \I__4443\ : Odrv4
    port map (
            O => \N__27066\,
            I => \nx.n2865\
        );

    \I__4442\ : InMux
    port map (
            O => \N__27063\,
            I => \nx.n10824\
        );

    \I__4441\ : CascadeMux
    port map (
            O => \N__27060\,
            I => \N__27056\
        );

    \I__4440\ : InMux
    port map (
            O => \N__27059\,
            I => \N__27053\
        );

    \I__4439\ : InMux
    port map (
            O => \N__27056\,
            I => \N__27050\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__27053\,
            I => \N__27045\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__27050\,
            I => \N__27045\
        );

    \I__4436\ : Odrv4
    port map (
            O => \N__27045\,
            I => \nx.n2797\
        );

    \I__4435\ : InMux
    port map (
            O => \N__27042\,
            I => \N__27039\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__27039\,
            I => \nx.n2864\
        );

    \I__4433\ : InMux
    port map (
            O => \N__27036\,
            I => \nx.n10825\
        );

    \I__4432\ : InMux
    port map (
            O => \N__27033\,
            I => \nx.n10826\
        );

    \I__4431\ : InMux
    port map (
            O => \N__27030\,
            I => \bfn_6_21_0_\
        );

    \I__4430\ : CascadeMux
    port map (
            O => \N__27027\,
            I => \N__27024\
        );

    \I__4429\ : InMux
    port map (
            O => \N__27024\,
            I => \N__27021\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__27021\,
            I => \N__27017\
        );

    \I__4427\ : CascadeMux
    port map (
            O => \N__27020\,
            I => \N__27014\
        );

    \I__4426\ : Span4Mux_h
    port map (
            O => \N__27017\,
            I => \N__27011\
        );

    \I__4425\ : InMux
    port map (
            O => \N__27014\,
            I => \N__27008\
        );

    \I__4424\ : Odrv4
    port map (
            O => \N__27011\,
            I => \nx.n2809\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__27008\,
            I => \nx.n2809\
        );

    \I__4422\ : InMux
    port map (
            O => \N__27003\,
            I => \N__27000\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__27000\,
            I => \N__26997\
        );

    \I__4420\ : Span12Mux_s11_v
    port map (
            O => \N__26997\,
            I => \N__26994\
        );

    \I__4419\ : Odrv12
    port map (
            O => \N__26994\,
            I => \nx.n2876\
        );

    \I__4418\ : InMux
    port map (
            O => \N__26991\,
            I => \nx.n10813\
        );

    \I__4417\ : CascadeMux
    port map (
            O => \N__26988\,
            I => \N__26983\
        );

    \I__4416\ : InMux
    port map (
            O => \N__26987\,
            I => \N__26978\
        );

    \I__4415\ : InMux
    port map (
            O => \N__26986\,
            I => \N__26978\
        );

    \I__4414\ : InMux
    port map (
            O => \N__26983\,
            I => \N__26975\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__26978\,
            I => \nx.n2808\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__26975\,
            I => \nx.n2808\
        );

    \I__4411\ : CascadeMux
    port map (
            O => \N__26970\,
            I => \N__26967\
        );

    \I__4410\ : InMux
    port map (
            O => \N__26967\,
            I => \N__26964\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__26964\,
            I => \nx.n2875\
        );

    \I__4408\ : InMux
    port map (
            O => \N__26961\,
            I => \nx.n10814\
        );

    \I__4407\ : CascadeMux
    port map (
            O => \N__26958\,
            I => \N__26954\
        );

    \I__4406\ : InMux
    port map (
            O => \N__26957\,
            I => \N__26950\
        );

    \I__4405\ : InMux
    port map (
            O => \N__26954\,
            I => \N__26947\
        );

    \I__4404\ : CascadeMux
    port map (
            O => \N__26953\,
            I => \N__26944\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__26950\,
            I => \N__26939\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__26947\,
            I => \N__26939\
        );

    \I__4401\ : InMux
    port map (
            O => \N__26944\,
            I => \N__26936\
        );

    \I__4400\ : Odrv4
    port map (
            O => \N__26939\,
            I => \nx.n2807\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__26936\,
            I => \nx.n2807\
        );

    \I__4398\ : InMux
    port map (
            O => \N__26931\,
            I => \N__26928\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__26928\,
            I => \nx.n2874\
        );

    \I__4396\ : InMux
    port map (
            O => \N__26925\,
            I => \nx.n10815\
        );

    \I__4395\ : InMux
    port map (
            O => \N__26922\,
            I => \nx.n10816\
        );

    \I__4394\ : CascadeMux
    port map (
            O => \N__26919\,
            I => \N__26915\
        );

    \I__4393\ : CascadeMux
    port map (
            O => \N__26918\,
            I => \N__26912\
        );

    \I__4392\ : InMux
    port map (
            O => \N__26915\,
            I => \N__26908\
        );

    \I__4391\ : InMux
    port map (
            O => \N__26912\,
            I => \N__26905\
        );

    \I__4390\ : InMux
    port map (
            O => \N__26911\,
            I => \N__26902\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__26908\,
            I => \N__26897\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__26905\,
            I => \N__26897\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__26902\,
            I => \nx.n2805\
        );

    \I__4386\ : Odrv4
    port map (
            O => \N__26897\,
            I => \nx.n2805\
        );

    \I__4385\ : InMux
    port map (
            O => \N__26892\,
            I => \N__26889\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__26889\,
            I => \nx.n2872\
        );

    \I__4383\ : InMux
    port map (
            O => \N__26886\,
            I => \nx.n10817\
        );

    \I__4382\ : InMux
    port map (
            O => \N__26883\,
            I => \nx.n10818\
        );

    \I__4381\ : InMux
    port map (
            O => \N__26880\,
            I => \N__26877\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__26877\,
            I => \nx.n29_adj_607\
        );

    \I__4379\ : CascadeMux
    port map (
            O => \N__26874\,
            I => \nx.n37_adj_608_cascade_\
        );

    \I__4378\ : InMux
    port map (
            O => \N__26871\,
            I => \N__26868\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__26868\,
            I => \nx.n40_adj_609\
        );

    \I__4376\ : CascadeMux
    port map (
            O => \N__26865\,
            I => \nx.n42_cascade_\
        );

    \I__4375\ : CascadeMux
    port map (
            O => \N__26862\,
            I => \nx.n2720_cascade_\
        );

    \I__4374\ : CascadeMux
    port map (
            O => \N__26859\,
            I => \nx.n2797_cascade_\
        );

    \I__4373\ : CascadeMux
    port map (
            O => \N__26856\,
            I => \nx.n2700_cascade_\
        );

    \I__4372\ : CascadeMux
    port map (
            O => \N__26853\,
            I => \nx.n2801_cascade_\
        );

    \I__4371\ : CascadeMux
    port map (
            O => \N__26850\,
            I => \N__26845\
        );

    \I__4370\ : InMux
    port map (
            O => \N__26849\,
            I => \N__26842\
        );

    \I__4369\ : InMux
    port map (
            O => \N__26848\,
            I => \N__26839\
        );

    \I__4368\ : InMux
    port map (
            O => \N__26845\,
            I => \N__26836\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__26842\,
            I => \nx.n1407\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__26839\,
            I => \nx.n1407\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__26836\,
            I => \nx.n1407\
        );

    \I__4364\ : CascadeMux
    port map (
            O => \N__26829\,
            I => \N__26826\
        );

    \I__4363\ : InMux
    port map (
            O => \N__26826\,
            I => \N__26823\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__26823\,
            I => \N__26820\
        );

    \I__4361\ : Odrv4
    port map (
            O => \N__26820\,
            I => \nx.n1474\
        );

    \I__4360\ : CascadeMux
    port map (
            O => \N__26817\,
            I => \nx.n1506_cascade_\
        );

    \I__4359\ : InMux
    port map (
            O => \N__26814\,
            I => \N__26811\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__26811\,
            I => \nx.n18_adj_632\
        );

    \I__4357\ : InMux
    port map (
            O => \N__26808\,
            I => \N__26805\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__26805\,
            I => \N__26802\
        );

    \I__4355\ : Odrv4
    port map (
            O => \N__26802\,
            I => \nx.n1475\
        );

    \I__4354\ : CascadeMux
    port map (
            O => \N__26799\,
            I => \N__26796\
        );

    \I__4353\ : InMux
    port map (
            O => \N__26796\,
            I => \N__26793\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__26793\,
            I => \N__26788\
        );

    \I__4351\ : InMux
    port map (
            O => \N__26792\,
            I => \N__26785\
        );

    \I__4350\ : CascadeMux
    port map (
            O => \N__26791\,
            I => \N__26782\
        );

    \I__4349\ : Span4Mux_s2_v
    port map (
            O => \N__26788\,
            I => \N__26779\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__26785\,
            I => \N__26776\
        );

    \I__4347\ : InMux
    port map (
            O => \N__26782\,
            I => \N__26773\
        );

    \I__4346\ : Odrv4
    port map (
            O => \N__26779\,
            I => \nx.n1408\
        );

    \I__4345\ : Odrv4
    port map (
            O => \N__26776\,
            I => \nx.n1408\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__26773\,
            I => \nx.n1408\
        );

    \I__4343\ : InMux
    port map (
            O => \N__26766\,
            I => \N__26762\
        );

    \I__4342\ : CascadeMux
    port map (
            O => \N__26765\,
            I => \N__26758\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__26762\,
            I => \N__26755\
        );

    \I__4340\ : InMux
    port map (
            O => \N__26761\,
            I => \N__26752\
        );

    \I__4339\ : InMux
    port map (
            O => \N__26758\,
            I => \N__26749\
        );

    \I__4338\ : Odrv4
    port map (
            O => \N__26755\,
            I => \nx.n1401\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__26752\,
            I => \nx.n1401\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__26749\,
            I => \nx.n1401\
        );

    \I__4335\ : InMux
    port map (
            O => \N__26742\,
            I => \N__26739\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__26739\,
            I => \N__26736\
        );

    \I__4333\ : Odrv4
    port map (
            O => \N__26736\,
            I => \nx.n1468\
        );

    \I__4332\ : InMux
    port map (
            O => \N__26733\,
            I => \N__26730\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__26730\,
            I => \N__26727\
        );

    \I__4330\ : Span4Mux_s1_v
    port map (
            O => \N__26727\,
            I => \N__26724\
        );

    \I__4329\ : Odrv4
    port map (
            O => \N__26724\,
            I => \nx.n1472\
        );

    \I__4328\ : CascadeMux
    port map (
            O => \N__26721\,
            I => \N__26716\
        );

    \I__4327\ : InMux
    port map (
            O => \N__26720\,
            I => \N__26713\
        );

    \I__4326\ : InMux
    port map (
            O => \N__26719\,
            I => \N__26710\
        );

    \I__4325\ : InMux
    port map (
            O => \N__26716\,
            I => \N__26707\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__26713\,
            I => \nx.n1405\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__26710\,
            I => \nx.n1405\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__26707\,
            I => \nx.n1405\
        );

    \I__4321\ : InMux
    port map (
            O => \N__26700\,
            I => \N__26697\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__26697\,
            I => \N__26694\
        );

    \I__4319\ : Span4Mux_s1_v
    port map (
            O => \N__26694\,
            I => \N__26691\
        );

    \I__4318\ : Odrv4
    port map (
            O => \N__26691\,
            I => \nx.n1473\
        );

    \I__4317\ : CascadeMux
    port map (
            O => \N__26688\,
            I => \N__26685\
        );

    \I__4316\ : InMux
    port map (
            O => \N__26685\,
            I => \N__26681\
        );

    \I__4315\ : CascadeMux
    port map (
            O => \N__26684\,
            I => \N__26678\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__26681\,
            I => \N__26674\
        );

    \I__4313\ : InMux
    port map (
            O => \N__26678\,
            I => \N__26671\
        );

    \I__4312\ : CascadeMux
    port map (
            O => \N__26677\,
            I => \N__26668\
        );

    \I__4311\ : Span4Mux_s2_v
    port map (
            O => \N__26674\,
            I => \N__26665\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__26671\,
            I => \N__26662\
        );

    \I__4309\ : InMux
    port map (
            O => \N__26668\,
            I => \N__26659\
        );

    \I__4308\ : Odrv4
    port map (
            O => \N__26665\,
            I => \nx.n1406\
        );

    \I__4307\ : Odrv4
    port map (
            O => \N__26662\,
            I => \nx.n1406\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__26659\,
            I => \nx.n1406\
        );

    \I__4305\ : CascadeMux
    port map (
            O => \N__26652\,
            I => \N__26648\
        );

    \I__4304\ : InMux
    port map (
            O => \N__26651\,
            I => \N__26643\
        );

    \I__4303\ : InMux
    port map (
            O => \N__26648\,
            I => \N__26640\
        );

    \I__4302\ : InMux
    port map (
            O => \N__26647\,
            I => \N__26637\
        );

    \I__4301\ : InMux
    port map (
            O => \N__26646\,
            I => \N__26634\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__26643\,
            I => \N__26629\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__26640\,
            I => \N__26629\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__26637\,
            I => \N__26626\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__26634\,
            I => \N__26621\
        );

    \I__4296\ : Span4Mux_v
    port map (
            O => \N__26629\,
            I => \N__26621\
        );

    \I__4295\ : Span4Mux_v
    port map (
            O => \N__26626\,
            I => \N__26618\
        );

    \I__4294\ : Odrv4
    port map (
            O => \N__26621\,
            I => neopxl_color_15
        );

    \I__4293\ : Odrv4
    port map (
            O => \N__26618\,
            I => neopxl_color_15
        );

    \I__4292\ : CascadeMux
    port map (
            O => \N__26613\,
            I => \nx.n9618_cascade_\
        );

    \I__4291\ : CascadeMux
    port map (
            O => \N__26610\,
            I => \N__26606\
        );

    \I__4290\ : InMux
    port map (
            O => \N__26609\,
            I => \N__26603\
        );

    \I__4289\ : InMux
    port map (
            O => \N__26606\,
            I => \N__26600\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__26603\,
            I => \nx.n608\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__26600\,
            I => \nx.n608\
        );

    \I__4286\ : CascadeMux
    port map (
            O => \N__26595\,
            I => \nx.n11738_cascade_\
        );

    \I__4285\ : InMux
    port map (
            O => \N__26592\,
            I => \N__26586\
        );

    \I__4284\ : InMux
    port map (
            O => \N__26591\,
            I => \N__26586\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__26586\,
            I => \nx.n708\
        );

    \I__4282\ : CascadeMux
    port map (
            O => \N__26583\,
            I => \nx.n739_cascade_\
        );

    \I__4281\ : InMux
    port map (
            O => \N__26580\,
            I => \N__26577\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__26577\,
            I => \nx.n11738\
        );

    \I__4279\ : InMux
    port map (
            O => \N__26574\,
            I => \N__26567\
        );

    \I__4278\ : InMux
    port map (
            O => \N__26573\,
            I => \N__26567\
        );

    \I__4277\ : InMux
    port map (
            O => \N__26572\,
            I => \N__26564\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__26567\,
            I => \nx.n807\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__26564\,
            I => \nx.n807\
        );

    \I__4274\ : CascadeMux
    port map (
            O => \N__26559\,
            I => \N__26554\
        );

    \I__4273\ : CascadeMux
    port map (
            O => \N__26558\,
            I => \N__26549\
        );

    \I__4272\ : InMux
    port map (
            O => \N__26557\,
            I => \N__26545\
        );

    \I__4271\ : InMux
    port map (
            O => \N__26554\,
            I => \N__26542\
        );

    \I__4270\ : InMux
    port map (
            O => \N__26553\,
            I => \N__26537\
        );

    \I__4269\ : InMux
    port map (
            O => \N__26552\,
            I => \N__26537\
        );

    \I__4268\ : InMux
    port map (
            O => \N__26549\,
            I => \N__26532\
        );

    \I__4267\ : InMux
    port map (
            O => \N__26548\,
            I => \N__26532\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__26545\,
            I => \nx.bit_ctr_31\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__26542\,
            I => \nx.bit_ctr_31\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__26537\,
            I => \nx.bit_ctr_31\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__26532\,
            I => \nx.bit_ctr_31\
        );

    \I__4262\ : CascadeMux
    port map (
            O => \N__26523\,
            I => \N__26519\
        );

    \I__4261\ : InMux
    port map (
            O => \N__26522\,
            I => \N__26515\
        );

    \I__4260\ : InMux
    port map (
            O => \N__26519\,
            I => \N__26510\
        );

    \I__4259\ : InMux
    port map (
            O => \N__26518\,
            I => \N__26510\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__26515\,
            I => \nx.n9618\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__26510\,
            I => \nx.n9618\
        );

    \I__4256\ : CascadeMux
    port map (
            O => \N__26505\,
            I => \N__26501\
        );

    \I__4255\ : InMux
    port map (
            O => \N__26504\,
            I => \N__26494\
        );

    \I__4254\ : InMux
    port map (
            O => \N__26501\,
            I => \N__26491\
        );

    \I__4253\ : InMux
    port map (
            O => \N__26500\,
            I => \N__26482\
        );

    \I__4252\ : InMux
    port map (
            O => \N__26499\,
            I => \N__26482\
        );

    \I__4251\ : InMux
    port map (
            O => \N__26498\,
            I => \N__26482\
        );

    \I__4250\ : InMux
    port map (
            O => \N__26497\,
            I => \N__26482\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__26494\,
            I => \nx.bit_ctr_29\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__26491\,
            I => \nx.bit_ctr_29\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__26482\,
            I => \nx.bit_ctr_29\
        );

    \I__4246\ : CascadeMux
    port map (
            O => \N__26475\,
            I => \nx.n11771_cascade_\
        );

    \I__4245\ : InMux
    port map (
            O => \N__26472\,
            I => \N__26469\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__26469\,
            I => \N__26466\
        );

    \I__4243\ : Odrv4
    port map (
            O => \N__26466\,
            I => \nx.n1470\
        );

    \I__4242\ : CascadeMux
    port map (
            O => \N__26463\,
            I => \N__26459\
        );

    \I__4241\ : CascadeMux
    port map (
            O => \N__26462\,
            I => \N__26456\
        );

    \I__4240\ : InMux
    port map (
            O => \N__26459\,
            I => \N__26452\
        );

    \I__4239\ : InMux
    port map (
            O => \N__26456\,
            I => \N__26449\
        );

    \I__4238\ : InMux
    port map (
            O => \N__26455\,
            I => \N__26446\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__26452\,
            I => \nx.n1403\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__26449\,
            I => \nx.n1403\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__26446\,
            I => \nx.n1403\
        );

    \I__4234\ : InMux
    port map (
            O => \N__26439\,
            I => \N__26434\
        );

    \I__4233\ : CascadeMux
    port map (
            O => \N__26438\,
            I => \N__26429\
        );

    \I__4232\ : InMux
    port map (
            O => \N__26437\,
            I => \N__26425\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__26434\,
            I => \N__26422\
        );

    \I__4230\ : InMux
    port map (
            O => \N__26433\,
            I => \N__26413\
        );

    \I__4229\ : InMux
    port map (
            O => \N__26432\,
            I => \N__26413\
        );

    \I__4228\ : InMux
    port map (
            O => \N__26429\,
            I => \N__26413\
        );

    \I__4227\ : InMux
    port map (
            O => \N__26428\,
            I => \N__26413\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__26425\,
            I => \nx.bit_ctr_30\
        );

    \I__4225\ : Odrv4
    port map (
            O => \N__26422\,
            I => \nx.bit_ctr_30\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__26413\,
            I => \nx.bit_ctr_30\
        );

    \I__4223\ : CascadeMux
    port map (
            O => \N__26406\,
            I => \N__26403\
        );

    \I__4222\ : InMux
    port map (
            O => \N__26403\,
            I => \N__26400\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__26400\,
            I => \N__26397\
        );

    \I__4220\ : Span4Mux_h
    port map (
            O => \N__26397\,
            I => \N__26394\
        );

    \I__4219\ : Odrv4
    port map (
            O => \N__26394\,
            I => \nx.n48_adj_704\
        );

    \I__4218\ : InMux
    port map (
            O => \N__26391\,
            I => \N__26386\
        );

    \I__4217\ : InMux
    port map (
            O => \N__26390\,
            I => \N__26381\
        );

    \I__4216\ : InMux
    port map (
            O => \N__26389\,
            I => \N__26381\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__26386\,
            I => \N__26378\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__26381\,
            I => \nx.n1008\
        );

    \I__4213\ : Odrv4
    port map (
            O => \N__26378\,
            I => \nx.n1008\
        );

    \I__4212\ : CascadeMux
    port map (
            O => \N__26373\,
            I => \nx.n7084_cascade_\
        );

    \I__4211\ : CascadeMux
    port map (
            O => \N__26370\,
            I => \nx.n838_cascade_\
        );

    \I__4210\ : CascadeMux
    port map (
            O => \N__26367\,
            I => \nx.n12595_cascade_\
        );

    \I__4209\ : CascadeMux
    port map (
            O => \N__26364\,
            I => \nx.n11617_cascade_\
        );

    \I__4208\ : InMux
    port map (
            O => \N__26361\,
            I => \N__26358\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__26358\,
            I => \nx.n1076\
        );

    \I__4206\ : CascadeMux
    port map (
            O => \N__26355\,
            I => \nx.n1037_cascade_\
        );

    \I__4205\ : CascadeMux
    port map (
            O => \N__26352\,
            I => \N__26348\
        );

    \I__4204\ : CascadeMux
    port map (
            O => \N__26351\,
            I => \N__26344\
        );

    \I__4203\ : InMux
    port map (
            O => \N__26348\,
            I => \N__26341\
        );

    \I__4202\ : InMux
    port map (
            O => \N__26347\,
            I => \N__26338\
        );

    \I__4201\ : InMux
    port map (
            O => \N__26344\,
            I => \N__26335\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__26341\,
            I => \N__26332\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__26338\,
            I => \N__26327\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__26335\,
            I => \N__26327\
        );

    \I__4197\ : Span4Mux_h
    port map (
            O => \N__26332\,
            I => \N__26324\
        );

    \I__4196\ : Span4Mux_h
    port map (
            O => \N__26327\,
            I => \N__26321\
        );

    \I__4195\ : Odrv4
    port map (
            O => \N__26324\,
            I => \nx.n1108\
        );

    \I__4194\ : Odrv4
    port map (
            O => \N__26321\,
            I => \nx.n1108\
        );

    \I__4193\ : CascadeMux
    port map (
            O => \N__26316\,
            I => \N__26312\
        );

    \I__4192\ : InMux
    port map (
            O => \N__26315\,
            I => \N__26309\
        );

    \I__4191\ : InMux
    port map (
            O => \N__26312\,
            I => \N__26306\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__26309\,
            I => \nx.n1007\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__26306\,
            I => \nx.n1007\
        );

    \I__4188\ : InMux
    port map (
            O => \N__26301\,
            I => \N__26298\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__26298\,
            I => \N__26295\
        );

    \I__4186\ : Odrv4
    port map (
            O => \N__26295\,
            I => \nx.n1074\
        );

    \I__4185\ : CascadeMux
    port map (
            O => \N__26292\,
            I => \N__26288\
        );

    \I__4184\ : InMux
    port map (
            O => \N__26291\,
            I => \N__26285\
        );

    \I__4183\ : InMux
    port map (
            O => \N__26288\,
            I => \N__26281\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__26285\,
            I => \N__26278\
        );

    \I__4181\ : InMux
    port map (
            O => \N__26284\,
            I => \N__26275\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__26281\,
            I => \N__26272\
        );

    \I__4179\ : Span4Mux_h
    port map (
            O => \N__26278\,
            I => \N__26269\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__26275\,
            I => \N__26266\
        );

    \I__4177\ : Span4Mux_h
    port map (
            O => \N__26272\,
            I => \N__26263\
        );

    \I__4176\ : Span4Mux_s2_v
    port map (
            O => \N__26269\,
            I => \N__26258\
        );

    \I__4175\ : Span4Mux_h
    port map (
            O => \N__26266\,
            I => \N__26258\
        );

    \I__4174\ : Odrv4
    port map (
            O => \N__26263\,
            I => \nx.n1106\
        );

    \I__4173\ : Odrv4
    port map (
            O => \N__26258\,
            I => \nx.n1106\
        );

    \I__4172\ : CascadeMux
    port map (
            O => \N__26253\,
            I => \N__26250\
        );

    \I__4171\ : InMux
    port map (
            O => \N__26250\,
            I => \N__26246\
        );

    \I__4170\ : InMux
    port map (
            O => \N__26249\,
            I => \N__26243\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__26246\,
            I => \N__26240\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__26243\,
            I => \nx.n1009\
        );

    \I__4167\ : Odrv4
    port map (
            O => \N__26240\,
            I => \nx.n1009\
        );

    \I__4166\ : CascadeMux
    port map (
            O => \N__26235\,
            I => \N__26232\
        );

    \I__4165\ : InMux
    port map (
            O => \N__26232\,
            I => \N__26227\
        );

    \I__4164\ : InMux
    port map (
            O => \N__26231\,
            I => \N__26224\
        );

    \I__4163\ : InMux
    port map (
            O => \N__26230\,
            I => \N__26220\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__26227\,
            I => \N__26216\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__26224\,
            I => \N__26213\
        );

    \I__4160\ : InMux
    port map (
            O => \N__26223\,
            I => \N__26210\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__26220\,
            I => \N__26207\
        );

    \I__4158\ : InMux
    port map (
            O => \N__26219\,
            I => \N__26204\
        );

    \I__4157\ : Span4Mux_v
    port map (
            O => \N__26216\,
            I => \N__26199\
        );

    \I__4156\ : Span4Mux_v
    port map (
            O => \N__26213\,
            I => \N__26199\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__26210\,
            I => \N__26196\
        );

    \I__4154\ : Span4Mux_v
    port map (
            O => \N__26207\,
            I => \N__26193\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__26204\,
            I => \nx.bit_ctr_25\
        );

    \I__4152\ : Odrv4
    port map (
            O => \N__26199\,
            I => \nx.bit_ctr_25\
        );

    \I__4151\ : Odrv4
    port map (
            O => \N__26196\,
            I => \nx.bit_ctr_25\
        );

    \I__4150\ : Odrv4
    port map (
            O => \N__26193\,
            I => \nx.bit_ctr_25\
        );

    \I__4149\ : CascadeMux
    port map (
            O => \N__26184\,
            I => \nx.n1009_cascade_\
        );

    \I__4148\ : InMux
    port map (
            O => \N__26181\,
            I => \N__26178\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__26178\,
            I => \nx.n7_adj_616\
        );

    \I__4146\ : InMux
    port map (
            O => \N__26175\,
            I => \N__26172\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__26172\,
            I => \N__26166\
        );

    \I__4144\ : InMux
    port map (
            O => \N__26171\,
            I => \N__26163\
        );

    \I__4143\ : InMux
    port map (
            O => \N__26170\,
            I => \N__26159\
        );

    \I__4142\ : InMux
    port map (
            O => \N__26169\,
            I => \N__26156\
        );

    \I__4141\ : Span4Mux_v
    port map (
            O => \N__26166\,
            I => \N__26153\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__26163\,
            I => \N__26150\
        );

    \I__4139\ : InMux
    port map (
            O => \N__26162\,
            I => \N__26147\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__26159\,
            I => \nx.bit_ctr_5\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__26156\,
            I => \nx.bit_ctr_5\
        );

    \I__4136\ : Odrv4
    port map (
            O => \N__26153\,
            I => \nx.bit_ctr_5\
        );

    \I__4135\ : Odrv12
    port map (
            O => \N__26150\,
            I => \nx.bit_ctr_5\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__26147\,
            I => \nx.bit_ctr_5\
        );

    \I__4133\ : InMux
    port map (
            O => \N__26136\,
            I => \N__26131\
        );

    \I__4132\ : InMux
    port map (
            O => \N__26135\,
            I => \N__26128\
        );

    \I__4131\ : InMux
    port map (
            O => \N__26134\,
            I => \N__26125\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__26131\,
            I => \N__26120\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__26128\,
            I => \N__26120\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__26125\,
            I => \N__26115\
        );

    \I__4127\ : Span4Mux_v
    port map (
            O => \N__26120\,
            I => \N__26112\
        );

    \I__4126\ : InMux
    port map (
            O => \N__26119\,
            I => \N__26109\
        );

    \I__4125\ : InMux
    port map (
            O => \N__26118\,
            I => \N__26106\
        );

    \I__4124\ : Span4Mux_v
    port map (
            O => \N__26115\,
            I => \N__26103\
        );

    \I__4123\ : Span4Mux_v
    port map (
            O => \N__26112\,
            I => \N__26100\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__26109\,
            I => \nx.bit_ctr_6\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__26106\,
            I => \nx.bit_ctr_6\
        );

    \I__4120\ : Odrv4
    port map (
            O => \N__26103\,
            I => \nx.bit_ctr_6\
        );

    \I__4119\ : Odrv4
    port map (
            O => \N__26100\,
            I => \nx.bit_ctr_6\
        );

    \I__4118\ : InMux
    port map (
            O => \N__26091\,
            I => \N__26088\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__26088\,
            I => \N__26085\
        );

    \I__4116\ : Odrv12
    port map (
            O => \N__26085\,
            I => \nx.n44_adj_708\
        );

    \I__4115\ : CascadeMux
    port map (
            O => \N__26082\,
            I => \N__26079\
        );

    \I__4114\ : InMux
    port map (
            O => \N__26079\,
            I => \N__26076\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__26076\,
            I => \N__26072\
        );

    \I__4112\ : InMux
    port map (
            O => \N__26075\,
            I => \N__26069\
        );

    \I__4111\ : Odrv4
    port map (
            O => \N__26072\,
            I => \nx.n1005\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__26069\,
            I => \nx.n1005\
        );

    \I__4109\ : InMux
    port map (
            O => \N__26064\,
            I => \N__26061\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__26061\,
            I => \N__26058\
        );

    \I__4107\ : Odrv4
    port map (
            O => \N__26058\,
            I => \nx.n1072\
        );

    \I__4106\ : CascadeMux
    port map (
            O => \N__26055\,
            I => \nx.n1005_cascade_\
        );

    \I__4105\ : InMux
    port map (
            O => \N__26052\,
            I => \N__26049\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__26049\,
            I => \N__26041\
        );

    \I__4103\ : InMux
    port map (
            O => \N__26048\,
            I => \N__26038\
        );

    \I__4102\ : InMux
    port map (
            O => \N__26047\,
            I => \N__26033\
        );

    \I__4101\ : InMux
    port map (
            O => \N__26046\,
            I => \N__26033\
        );

    \I__4100\ : InMux
    port map (
            O => \N__26045\,
            I => \N__26028\
        );

    \I__4099\ : InMux
    port map (
            O => \N__26044\,
            I => \N__26028\
        );

    \I__4098\ : Span4Mux_h
    port map (
            O => \N__26041\,
            I => \N__26025\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__26038\,
            I => \nx.n1037\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__26033\,
            I => \nx.n1037\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__26028\,
            I => \nx.n1037\
        );

    \I__4094\ : Odrv4
    port map (
            O => \N__26025\,
            I => \nx.n1037\
        );

    \I__4093\ : CascadeMux
    port map (
            O => \N__26016\,
            I => \N__26013\
        );

    \I__4092\ : InMux
    port map (
            O => \N__26013\,
            I => \N__26008\
        );

    \I__4091\ : InMux
    port map (
            O => \N__26012\,
            I => \N__26005\
        );

    \I__4090\ : InMux
    port map (
            O => \N__26011\,
            I => \N__26002\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__26008\,
            I => \N__25999\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__26005\,
            I => \N__25994\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__26002\,
            I => \N__25994\
        );

    \I__4086\ : Span4Mux_h
    port map (
            O => \N__25999\,
            I => \N__25991\
        );

    \I__4085\ : Span4Mux_h
    port map (
            O => \N__25994\,
            I => \N__25988\
        );

    \I__4084\ : Odrv4
    port map (
            O => \N__25991\,
            I => \nx.n1104\
        );

    \I__4083\ : Odrv4
    port map (
            O => \N__25988\,
            I => \nx.n1104\
        );

    \I__4082\ : InMux
    port map (
            O => \N__25983\,
            I => \nx.n10472\
        );

    \I__4081\ : InMux
    port map (
            O => \N__25980\,
            I => \nx.n10473\
        );

    \I__4080\ : CascadeMux
    port map (
            O => \N__25977\,
            I => \N__25973\
        );

    \I__4079\ : InMux
    port map (
            O => \N__25976\,
            I => \N__25970\
        );

    \I__4078\ : InMux
    port map (
            O => \N__25973\,
            I => \N__25967\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__25970\,
            I => \N__25964\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__25967\,
            I => \N__25959\
        );

    \I__4075\ : Span4Mux_s1_h
    port map (
            O => \N__25964\,
            I => \N__25959\
        );

    \I__4074\ : Span4Mux_v
    port map (
            O => \N__25959\,
            I => \N__25956\
        );

    \I__4073\ : Odrv4
    port map (
            O => \N__25956\,
            I => \nx.n1103\
        );

    \I__4072\ : InMux
    port map (
            O => \N__25953\,
            I => \N__25950\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__25950\,
            I => \N__25947\
        );

    \I__4070\ : Span4Mux_h
    port map (
            O => \N__25947\,
            I => \N__25944\
        );

    \I__4069\ : Odrv4
    port map (
            O => \N__25944\,
            I => \nx.n46_adj_705\
        );

    \I__4068\ : InMux
    port map (
            O => \N__25941\,
            I => \N__25938\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__25938\,
            I => \nx.n1075\
        );

    \I__4066\ : CascadeMux
    port map (
            O => \N__25935\,
            I => \N__25932\
        );

    \I__4065\ : InMux
    port map (
            O => \N__25932\,
            I => \N__25927\
        );

    \I__4064\ : InMux
    port map (
            O => \N__25931\,
            I => \N__25924\
        );

    \I__4063\ : CascadeMux
    port map (
            O => \N__25930\,
            I => \N__25921\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__25927\,
            I => \N__25916\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__25924\,
            I => \N__25916\
        );

    \I__4060\ : InMux
    port map (
            O => \N__25921\,
            I => \N__25913\
        );

    \I__4059\ : Span4Mux_s3_v
    port map (
            O => \N__25916\,
            I => \N__25908\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__25913\,
            I => \N__25908\
        );

    \I__4057\ : Span4Mux_h
    port map (
            O => \N__25908\,
            I => \N__25905\
        );

    \I__4056\ : Odrv4
    port map (
            O => \N__25905\,
            I => \nx.n1107\
        );

    \I__4055\ : InMux
    port map (
            O => \N__25902\,
            I => \N__25899\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__25899\,
            I => \nx.n1073\
        );

    \I__4053\ : CascadeMux
    port map (
            O => \N__25896\,
            I => \N__25891\
        );

    \I__4052\ : InMux
    port map (
            O => \N__25895\,
            I => \N__25888\
        );

    \I__4051\ : InMux
    port map (
            O => \N__25894\,
            I => \N__25885\
        );

    \I__4050\ : InMux
    port map (
            O => \N__25891\,
            I => \N__25882\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__25888\,
            I => \N__25875\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__25885\,
            I => \N__25875\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__25882\,
            I => \N__25875\
        );

    \I__4046\ : Span4Mux_v
    port map (
            O => \N__25875\,
            I => \N__25872\
        );

    \I__4045\ : Odrv4
    port map (
            O => \N__25872\,
            I => \nx.n1105\
        );

    \I__4044\ : CascadeMux
    port map (
            O => \N__25869\,
            I => \N__25865\
        );

    \I__4043\ : InMux
    port map (
            O => \N__25868\,
            I => \N__25862\
        );

    \I__4042\ : InMux
    port map (
            O => \N__25865\,
            I => \N__25859\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__25862\,
            I => \N__25854\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__25859\,
            I => \N__25854\
        );

    \I__4039\ : Span4Mux_v
    port map (
            O => \N__25854\,
            I => \N__25851\
        );

    \I__4038\ : Odrv4
    port map (
            O => \N__25851\,
            I => \nx.n2894\
        );

    \I__4037\ : CascadeMux
    port map (
            O => \N__25848\,
            I => \N__25845\
        );

    \I__4036\ : InMux
    port map (
            O => \N__25845\,
            I => \N__25842\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__25842\,
            I => \N__25838\
        );

    \I__4034\ : InMux
    port map (
            O => \N__25841\,
            I => \N__25835\
        );

    \I__4033\ : Span4Mux_h
    port map (
            O => \N__25838\,
            I => \N__25832\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__25835\,
            I => \nx.n2993\
        );

    \I__4031\ : Odrv4
    port map (
            O => \N__25832\,
            I => \nx.n2993\
        );

    \I__4030\ : InMux
    port map (
            O => \N__25827\,
            I => \N__25824\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__25824\,
            I => \N__25821\
        );

    \I__4028\ : Span4Mux_h
    port map (
            O => \N__25821\,
            I => \N__25818\
        );

    \I__4027\ : Odrv4
    port map (
            O => \N__25818\,
            I => \nx.n3060\
        );

    \I__4026\ : CascadeMux
    port map (
            O => \N__25815\,
            I => \nx.n2993_cascade_\
        );

    \I__4025\ : InMux
    port map (
            O => \N__25812\,
            I => \N__25809\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__25809\,
            I => \N__25805\
        );

    \I__4023\ : InMux
    port map (
            O => \N__25808\,
            I => \N__25802\
        );

    \I__4022\ : Span12Mux_s4_h
    port map (
            O => \N__25805\,
            I => \N__25799\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__25802\,
            I => \nx.n3092\
        );

    \I__4020\ : Odrv12
    port map (
            O => \N__25799\,
            I => \nx.n3092\
        );

    \I__4019\ : InMux
    port map (
            O => \N__25794\,
            I => \N__25790\
        );

    \I__4018\ : InMux
    port map (
            O => \N__25793\,
            I => \N__25787\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__25790\,
            I => \N__25784\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__25787\,
            I => \N__25780\
        );

    \I__4015\ : Span4Mux_v
    port map (
            O => \N__25784\,
            I => \N__25777\
        );

    \I__4014\ : InMux
    port map (
            O => \N__25783\,
            I => \N__25774\
        );

    \I__4013\ : Span4Mux_h
    port map (
            O => \N__25780\,
            I => \N__25771\
        );

    \I__4012\ : Odrv4
    port map (
            O => \N__25777\,
            I => \nx.n3091\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__25774\,
            I => \nx.n3091\
        );

    \I__4010\ : Odrv4
    port map (
            O => \N__25771\,
            I => \nx.n3091\
        );

    \I__4009\ : CascadeMux
    port map (
            O => \N__25764\,
            I => \nx.n3092_cascade_\
        );

    \I__4008\ : InMux
    port map (
            O => \N__25761\,
            I => \N__25758\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__25758\,
            I => \N__25755\
        );

    \I__4006\ : Span4Mux_h
    port map (
            O => \N__25755\,
            I => \N__25752\
        );

    \I__4005\ : Odrv4
    port map (
            O => \N__25752\,
            I => \nx.n46_adj_688\
        );

    \I__4004\ : InMux
    port map (
            O => \N__25749\,
            I => \N__25746\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__25746\,
            I => \N__25743\
        );

    \I__4002\ : Span4Mux_s1_h
    port map (
            O => \N__25743\,
            I => \N__25740\
        );

    \I__4001\ : Odrv4
    port map (
            O => \N__25740\,
            I => \nx.n50\
        );

    \I__4000\ : InMux
    port map (
            O => \N__25737\,
            I => \N__25734\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__25734\,
            I => \N__25730\
        );

    \I__3998\ : InMux
    port map (
            O => \N__25733\,
            I => \N__25726\
        );

    \I__3997\ : Span4Mux_h
    port map (
            O => \N__25730\,
            I => \N__25723\
        );

    \I__3996\ : InMux
    port map (
            O => \N__25729\,
            I => \N__25720\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__25726\,
            I => \nx.n3093\
        );

    \I__3994\ : Odrv4
    port map (
            O => \N__25723\,
            I => \nx.n3093\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__25720\,
            I => \nx.n3093\
        );

    \I__3992\ : InMux
    port map (
            O => \N__25713\,
            I => \N__25710\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__25710\,
            I => \nx.n36_adj_687\
        );

    \I__3990\ : InMux
    port map (
            O => \N__25707\,
            I => \N__25704\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__25704\,
            I => \N__25701\
        );

    \I__3988\ : Span12Mux_s6_v
    port map (
            O => \N__25701\,
            I => \N__25698\
        );

    \I__3987\ : Odrv12
    port map (
            O => \N__25698\,
            I => \nx.n1077\
        );

    \I__3986\ : InMux
    port map (
            O => \N__25695\,
            I => \bfn_5_26_0_\
        );

    \I__3985\ : InMux
    port map (
            O => \N__25692\,
            I => \nx.n10468\
        );

    \I__3984\ : InMux
    port map (
            O => \N__25689\,
            I => \nx.n10469\
        );

    \I__3983\ : InMux
    port map (
            O => \N__25686\,
            I => \nx.n10470\
        );

    \I__3982\ : InMux
    port map (
            O => \N__25683\,
            I => \nx.n10471\
        );

    \I__3981\ : InMux
    port map (
            O => \N__25680\,
            I => \N__25677\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__25677\,
            I => \nx.n2959\
        );

    \I__3979\ : InMux
    port map (
            O => \N__25674\,
            I => \nx.n10854\
        );

    \I__3978\ : CascadeMux
    port map (
            O => \N__25671\,
            I => \N__25668\
        );

    \I__3977\ : InMux
    port map (
            O => \N__25668\,
            I => \N__25665\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__25665\,
            I => \nx.n2958\
        );

    \I__3975\ : InMux
    port map (
            O => \N__25662\,
            I => \nx.n10855\
        );

    \I__3974\ : InMux
    port map (
            O => \N__25659\,
            I => \N__25656\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__25656\,
            I => \nx.n2957\
        );

    \I__3972\ : InMux
    port map (
            O => \N__25653\,
            I => \nx.n10856\
        );

    \I__3971\ : InMux
    port map (
            O => \N__25650\,
            I => \N__25647\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__25647\,
            I => \nx.n2956\
        );

    \I__3969\ : InMux
    port map (
            O => \N__25644\,
            I => \nx.n10857\
        );

    \I__3968\ : InMux
    port map (
            O => \N__25641\,
            I => \N__25638\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__25638\,
            I => \nx.n2955\
        );

    \I__3966\ : InMux
    port map (
            O => \N__25635\,
            I => \nx.n10858\
        );

    \I__3965\ : InMux
    port map (
            O => \N__25632\,
            I => \N__25629\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__25629\,
            I => \N__25626\
        );

    \I__3963\ : Odrv4
    port map (
            O => \N__25626\,
            I => \nx.n2954\
        );

    \I__3962\ : InMux
    port map (
            O => \N__25623\,
            I => \nx.n10859\
        );

    \I__3961\ : InMux
    port map (
            O => \N__25620\,
            I => \N__25617\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__25617\,
            I => \N__25614\
        );

    \I__3959\ : Odrv4
    port map (
            O => \N__25614\,
            I => \nx.n2953\
        );

    \I__3958\ : InMux
    port map (
            O => \N__25611\,
            I => \bfn_5_25_0_\
        );

    \I__3957\ : InMux
    port map (
            O => \N__25608\,
            I => \nx.n10861\
        );

    \I__3956\ : InMux
    port map (
            O => \N__25605\,
            I => \N__25602\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__25602\,
            I => \N__25598\
        );

    \I__3954\ : InMux
    port map (
            O => \N__25601\,
            I => \N__25595\
        );

    \I__3953\ : Span4Mux_v
    port map (
            O => \N__25598\,
            I => \N__25592\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__25595\,
            I => \N__25589\
        );

    \I__3951\ : Odrv4
    port map (
            O => \N__25592\,
            I => \nx.n2984\
        );

    \I__3950\ : Odrv4
    port map (
            O => \N__25589\,
            I => \nx.n2984\
        );

    \I__3949\ : InMux
    port map (
            O => \N__25584\,
            I => \N__25581\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__25581\,
            I => \nx.n2961\
        );

    \I__3947\ : CascadeMux
    port map (
            O => \N__25578\,
            I => \N__25575\
        );

    \I__3946\ : InMux
    port map (
            O => \N__25575\,
            I => \N__25572\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__25572\,
            I => \N__25569\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__25569\,
            I => \nx.n2967\
        );

    \I__3943\ : InMux
    port map (
            O => \N__25566\,
            I => \nx.n10846\
        );

    \I__3942\ : CascadeMux
    port map (
            O => \N__25563\,
            I => \N__25560\
        );

    \I__3941\ : InMux
    port map (
            O => \N__25560\,
            I => \N__25556\
        );

    \I__3940\ : InMux
    port map (
            O => \N__25559\,
            I => \N__25553\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__25556\,
            I => \nx.n2899\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__25553\,
            I => \nx.n2899\
        );

    \I__3937\ : InMux
    port map (
            O => \N__25548\,
            I => \N__25545\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__25545\,
            I => \nx.n2966\
        );

    \I__3935\ : InMux
    port map (
            O => \N__25542\,
            I => \nx.n10847\
        );

    \I__3934\ : CascadeMux
    port map (
            O => \N__25539\,
            I => \N__25535\
        );

    \I__3933\ : InMux
    port map (
            O => \N__25538\,
            I => \N__25532\
        );

    \I__3932\ : InMux
    port map (
            O => \N__25535\,
            I => \N__25529\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__25532\,
            I => \N__25526\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__25529\,
            I => \N__25523\
        );

    \I__3929\ : Odrv4
    port map (
            O => \N__25526\,
            I => \nx.n2898\
        );

    \I__3928\ : Odrv4
    port map (
            O => \N__25523\,
            I => \nx.n2898\
        );

    \I__3927\ : CascadeMux
    port map (
            O => \N__25518\,
            I => \N__25515\
        );

    \I__3926\ : InMux
    port map (
            O => \N__25515\,
            I => \N__25512\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__25512\,
            I => \nx.n2965\
        );

    \I__3924\ : InMux
    port map (
            O => \N__25509\,
            I => \nx.n10848\
        );

    \I__3923\ : CascadeMux
    port map (
            O => \N__25506\,
            I => \N__25502\
        );

    \I__3922\ : CascadeMux
    port map (
            O => \N__25505\,
            I => \N__25499\
        );

    \I__3921\ : InMux
    port map (
            O => \N__25502\,
            I => \N__25496\
        );

    \I__3920\ : InMux
    port map (
            O => \N__25499\,
            I => \N__25493\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__25496\,
            I => \N__25487\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__25493\,
            I => \N__25487\
        );

    \I__3917\ : InMux
    port map (
            O => \N__25492\,
            I => \N__25484\
        );

    \I__3916\ : Odrv4
    port map (
            O => \N__25487\,
            I => \nx.n2897\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__25484\,
            I => \nx.n2897\
        );

    \I__3914\ : InMux
    port map (
            O => \N__25479\,
            I => \N__25476\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__25476\,
            I => \nx.n2964\
        );

    \I__3912\ : InMux
    port map (
            O => \N__25473\,
            I => \nx.n10849\
        );

    \I__3911\ : CascadeMux
    port map (
            O => \N__25470\,
            I => \N__25466\
        );

    \I__3910\ : InMux
    port map (
            O => \N__25469\,
            I => \N__25463\
        );

    \I__3909\ : InMux
    port map (
            O => \N__25466\,
            I => \N__25460\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__25463\,
            I => \N__25457\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__25460\,
            I => \nx.n2896\
        );

    \I__3906\ : Odrv4
    port map (
            O => \N__25457\,
            I => \nx.n2896\
        );

    \I__3905\ : InMux
    port map (
            O => \N__25452\,
            I => \N__25449\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__25449\,
            I => \N__25446\
        );

    \I__3903\ : Odrv4
    port map (
            O => \N__25446\,
            I => \nx.n2963\
        );

    \I__3902\ : InMux
    port map (
            O => \N__25443\,
            I => \nx.n10850\
        );

    \I__3901\ : InMux
    port map (
            O => \N__25440\,
            I => \N__25437\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__25437\,
            I => \nx.n2962\
        );

    \I__3899\ : InMux
    port map (
            O => \N__25434\,
            I => \nx.n10851\
        );

    \I__3898\ : InMux
    port map (
            O => \N__25431\,
            I => \bfn_5_24_0_\
        );

    \I__3897\ : InMux
    port map (
            O => \N__25428\,
            I => \N__25425\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__25425\,
            I => \nx.n2960\
        );

    \I__3895\ : InMux
    port map (
            O => \N__25422\,
            I => \nx.n10853\
        );

    \I__3894\ : CascadeMux
    port map (
            O => \N__25419\,
            I => \N__25416\
        );

    \I__3893\ : InMux
    port map (
            O => \N__25416\,
            I => \N__25412\
        );

    \I__3892\ : InMux
    port map (
            O => \N__25415\,
            I => \N__25409\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__25412\,
            I => \N__25404\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__25409\,
            I => \N__25404\
        );

    \I__3889\ : Span4Mux_v
    port map (
            O => \N__25404\,
            I => \N__25401\
        );

    \I__3888\ : Odrv4
    port map (
            O => \N__25401\,
            I => \nx.n2908\
        );

    \I__3887\ : InMux
    port map (
            O => \N__25398\,
            I => \N__25395\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__25395\,
            I => \N__25392\
        );

    \I__3885\ : Span4Mux_h
    port map (
            O => \N__25392\,
            I => \N__25389\
        );

    \I__3884\ : Odrv4
    port map (
            O => \N__25389\,
            I => \nx.n2975\
        );

    \I__3883\ : InMux
    port map (
            O => \N__25386\,
            I => \nx.n10838\
        );

    \I__3882\ : CascadeMux
    port map (
            O => \N__25383\,
            I => \N__25379\
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__25382\,
            I => \N__25376\
        );

    \I__3880\ : InMux
    port map (
            O => \N__25379\,
            I => \N__25373\
        );

    \I__3879\ : InMux
    port map (
            O => \N__25376\,
            I => \N__25369\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__25373\,
            I => \N__25366\
        );

    \I__3877\ : InMux
    port map (
            O => \N__25372\,
            I => \N__25363\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__25369\,
            I => \nx.n2907\
        );

    \I__3875\ : Odrv4
    port map (
            O => \N__25366\,
            I => \nx.n2907\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__25363\,
            I => \nx.n2907\
        );

    \I__3873\ : InMux
    port map (
            O => \N__25356\,
            I => \N__25353\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__25353\,
            I => \nx.n2974\
        );

    \I__3871\ : InMux
    port map (
            O => \N__25350\,
            I => \nx.n10839\
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__25347\,
            I => \N__25343\
        );

    \I__3869\ : InMux
    port map (
            O => \N__25346\,
            I => \N__25339\
        );

    \I__3868\ : InMux
    port map (
            O => \N__25343\,
            I => \N__25336\
        );

    \I__3867\ : InMux
    port map (
            O => \N__25342\,
            I => \N__25333\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__25339\,
            I => \nx.n2906\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__25336\,
            I => \nx.n2906\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__25333\,
            I => \nx.n2906\
        );

    \I__3863\ : InMux
    port map (
            O => \N__25326\,
            I => \N__25323\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__25323\,
            I => \nx.n2973\
        );

    \I__3861\ : InMux
    port map (
            O => \N__25320\,
            I => \nx.n10840\
        );

    \I__3860\ : InMux
    port map (
            O => \N__25317\,
            I => \N__25314\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__25314\,
            I => \N__25311\
        );

    \I__3858\ : Odrv4
    port map (
            O => \N__25311\,
            I => \nx.n2972\
        );

    \I__3857\ : InMux
    port map (
            O => \N__25308\,
            I => \nx.n10841\
        );

    \I__3856\ : InMux
    port map (
            O => \N__25305\,
            I => \nx.n10842\
        );

    \I__3855\ : CascadeMux
    port map (
            O => \N__25302\,
            I => \N__25299\
        );

    \I__3854\ : InMux
    port map (
            O => \N__25299\,
            I => \N__25296\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__25296\,
            I => \N__25293\
        );

    \I__3852\ : Odrv4
    port map (
            O => \N__25293\,
            I => \nx.n2970\
        );

    \I__3851\ : InMux
    port map (
            O => \N__25290\,
            I => \nx.n10843\
        );

    \I__3850\ : CascadeMux
    port map (
            O => \N__25287\,
            I => \N__25284\
        );

    \I__3849\ : InMux
    port map (
            O => \N__25284\,
            I => \N__25281\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__25281\,
            I => \N__25278\
        );

    \I__3847\ : Span4Mux_s2_h
    port map (
            O => \N__25278\,
            I => \N__25275\
        );

    \I__3846\ : Odrv4
    port map (
            O => \N__25275\,
            I => \nx.n2969\
        );

    \I__3845\ : InMux
    port map (
            O => \N__25272\,
            I => \bfn_5_23_0_\
        );

    \I__3844\ : CascadeMux
    port map (
            O => \N__25269\,
            I => \N__25265\
        );

    \I__3843\ : InMux
    port map (
            O => \N__25268\,
            I => \N__25262\
        );

    \I__3842\ : InMux
    port map (
            O => \N__25265\,
            I => \N__25259\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__25262\,
            I => \N__25253\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__25259\,
            I => \N__25253\
        );

    \I__3839\ : InMux
    port map (
            O => \N__25258\,
            I => \N__25250\
        );

    \I__3838\ : Odrv4
    port map (
            O => \N__25253\,
            I => \nx.n2901\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__25250\,
            I => \nx.n2901\
        );

    \I__3836\ : InMux
    port map (
            O => \N__25245\,
            I => \N__25242\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__25242\,
            I => \nx.n2968\
        );

    \I__3834\ : InMux
    port map (
            O => \N__25239\,
            I => \nx.n10845\
        );

    \I__3833\ : CascadeMux
    port map (
            O => \N__25236\,
            I => \nx.n2896_cascade_\
        );

    \I__3832\ : CascadeMux
    port map (
            O => \N__25233\,
            I => \nx.n2898_cascade_\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__25230\,
            I => \nx.n42_adj_675_cascade_\
        );

    \I__3830\ : InMux
    port map (
            O => \N__25227\,
            I => \N__25224\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__25224\,
            I => \nx.n32_adj_674\
        );

    \I__3828\ : InMux
    port map (
            O => \N__25221\,
            I => \N__25218\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__25218\,
            I => \N__25215\
        );

    \I__3826\ : Odrv4
    port map (
            O => \N__25215\,
            I => \nx.n46\
        );

    \I__3825\ : InMux
    port map (
            O => \N__25212\,
            I => \N__25209\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__25209\,
            I => \N__25206\
        );

    \I__3823\ : Span4Mux_v
    port map (
            O => \N__25206\,
            I => \N__25203\
        );

    \I__3822\ : Odrv4
    port map (
            O => \N__25203\,
            I => \nx.n2977\
        );

    \I__3821\ : InMux
    port map (
            O => \N__25200\,
            I => \bfn_5_22_0_\
        );

    \I__3820\ : CascadeMux
    port map (
            O => \N__25197\,
            I => \N__25194\
        );

    \I__3819\ : InMux
    port map (
            O => \N__25194\,
            I => \N__25191\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__25191\,
            I => \N__25188\
        );

    \I__3817\ : Span4Mux_h
    port map (
            O => \N__25188\,
            I => \N__25185\
        );

    \I__3816\ : Odrv4
    port map (
            O => \N__25185\,
            I => \nx.n2976\
        );

    \I__3815\ : InMux
    port map (
            O => \N__25182\,
            I => \nx.n10837\
        );

    \I__3814\ : CascadeMux
    port map (
            O => \N__25179\,
            I => \N__25176\
        );

    \I__3813\ : InMux
    port map (
            O => \N__25176\,
            I => \N__25172\
        );

    \I__3812\ : InMux
    port map (
            O => \N__25175\,
            I => \N__25169\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__25172\,
            I => \N__25165\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__25169\,
            I => \N__25162\
        );

    \I__3809\ : InMux
    port map (
            O => \N__25168\,
            I => \N__25159\
        );

    \I__3808\ : Span4Mux_v
    port map (
            O => \N__25165\,
            I => \N__25156\
        );

    \I__3807\ : Odrv4
    port map (
            O => \N__25162\,
            I => timer_20
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__25159\,
            I => timer_20
        );

    \I__3805\ : Odrv4
    port map (
            O => \N__25156\,
            I => timer_20
        );

    \I__3804\ : InMux
    port map (
            O => \N__25149\,
            I => \N__25143\
        );

    \I__3803\ : InMux
    port map (
            O => \N__25148\,
            I => \N__25143\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__25143\,
            I => neo_pixel_transmitter_t0_20
        );

    \I__3801\ : CascadeMux
    port map (
            O => \N__25140\,
            I => \nx.n2809_cascade_\
        );

    \I__3800\ : CascadeMux
    port map (
            O => \N__25137\,
            I => \nx.n31_adj_613_cascade_\
        );

    \I__3799\ : InMux
    port map (
            O => \N__25134\,
            I => \N__25131\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__25131\,
            I => \nx.n39_adj_614\
        );

    \I__3797\ : InMux
    port map (
            O => \N__25128\,
            I => \N__25125\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__25125\,
            I => \N__25121\
        );

    \I__3795\ : InMux
    port map (
            O => \N__25124\,
            I => \N__25117\
        );

    \I__3794\ : Span4Mux_v
    port map (
            O => \N__25121\,
            I => \N__25114\
        );

    \I__3793\ : InMux
    port map (
            O => \N__25120\,
            I => \N__25111\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__25117\,
            I => \N__25108\
        );

    \I__3791\ : Odrv4
    port map (
            O => \N__25114\,
            I => timer_19
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__25111\,
            I => timer_19
        );

    \I__3789\ : Odrv12
    port map (
            O => \N__25108\,
            I => timer_19
        );

    \I__3788\ : InMux
    port map (
            O => \N__25101\,
            I => \N__25098\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__25098\,
            I => \N__25095\
        );

    \I__3786\ : Odrv4
    port map (
            O => \N__25095\,
            I => n13171
        );

    \I__3785\ : InMux
    port map (
            O => \N__25092\,
            I => \N__25089\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__25089\,
            I => n13170
        );

    \I__3783\ : InMux
    port map (
            O => \N__25086\,
            I => \N__25082\
        );

    \I__3782\ : InMux
    port map (
            O => \N__25085\,
            I => \N__25079\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__25082\,
            I => neo_pixel_transmitter_t0_9
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__25079\,
            I => neo_pixel_transmitter_t0_9
        );

    \I__3779\ : InMux
    port map (
            O => \N__25074\,
            I => \N__25071\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__25071\,
            I => \N__25068\
        );

    \I__3777\ : Span4Mux_v
    port map (
            O => \N__25068\,
            I => \N__25065\
        );

    \I__3776\ : Span4Mux_s2_h
    port map (
            O => \N__25065\,
            I => \N__25062\
        );

    \I__3775\ : Odrv4
    port map (
            O => \N__25062\,
            I => \nx.n24\
        );

    \I__3774\ : InMux
    port map (
            O => \N__25059\,
            I => \N__25055\
        );

    \I__3773\ : InMux
    port map (
            O => \N__25058\,
            I => \N__25052\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__25055\,
            I => neo_pixel_transmitter_t0_19
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__25052\,
            I => neo_pixel_transmitter_t0_19
        );

    \I__3770\ : CascadeMux
    port map (
            O => \N__25047\,
            I => \N__25044\
        );

    \I__3769\ : InMux
    port map (
            O => \N__25044\,
            I => \N__25041\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__25041\,
            I => \N__25038\
        );

    \I__3767\ : Span4Mux_h
    port map (
            O => \N__25038\,
            I => \N__25035\
        );

    \I__3766\ : Span4Mux_v
    port map (
            O => \N__25035\,
            I => \N__25032\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__25032\,
            I => \nx.n14\
        );

    \I__3764\ : InMux
    port map (
            O => \N__25029\,
            I => \N__25026\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__25026\,
            I => neopxl_color_prev_6
        );

    \I__3762\ : InMux
    port map (
            O => \N__25023\,
            I => \N__25020\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__25020\,
            I => \N__25017\
        );

    \I__3760\ : Odrv4
    port map (
            O => \N__25017\,
            I => neopxl_color_prev_15
        );

    \I__3759\ : InMux
    port map (
            O => \N__25014\,
            I => \N__25011\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__25011\,
            I => \N__25008\
        );

    \I__3757\ : Odrv12
    port map (
            O => \N__25008\,
            I => n11_adj_775
        );

    \I__3756\ : CascadeMux
    port map (
            O => \N__25005\,
            I => \N__25002\
        );

    \I__3755\ : InMux
    port map (
            O => \N__25002\,
            I => \N__24999\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__24999\,
            I => \N__24996\
        );

    \I__3753\ : Span4Mux_v
    port map (
            O => \N__24996\,
            I => \N__24993\
        );

    \I__3752\ : Odrv4
    port map (
            O => \N__24993\,
            I => neopxl_color_prev_13
        );

    \I__3751\ : InMux
    port map (
            O => \N__24990\,
            I => \N__24987\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__24987\,
            I => \N__24984\
        );

    \I__3749\ : Span4Mux_h
    port map (
            O => \N__24984\,
            I => \N__24981\
        );

    \I__3748\ : Span4Mux_v
    port map (
            O => \N__24981\,
            I => \N__24978\
        );

    \I__3747\ : Odrv4
    port map (
            O => \N__24978\,
            I => \nx.n13_adj_649\
        );

    \I__3746\ : InMux
    port map (
            O => \N__24975\,
            I => \N__24972\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__24972\,
            I => \N__24965\
        );

    \I__3744\ : InMux
    port map (
            O => \N__24971\,
            I => \N__24962\
        );

    \I__3743\ : InMux
    port map (
            O => \N__24970\,
            I => \N__24959\
        );

    \I__3742\ : InMux
    port map (
            O => \N__24969\,
            I => \N__24956\
        );

    \I__3741\ : InMux
    port map (
            O => \N__24968\,
            I => \N__24953\
        );

    \I__3740\ : Span4Mux_s1_v
    port map (
            O => \N__24965\,
            I => \N__24946\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__24962\,
            I => \N__24946\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__24959\,
            I => \N__24946\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__24956\,
            I => \nx.bit_ctr_21\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__24953\,
            I => \nx.bit_ctr_21\
        );

    \I__3735\ : Odrv4
    port map (
            O => \N__24946\,
            I => \nx.bit_ctr_21\
        );

    \I__3734\ : InMux
    port map (
            O => \N__24939\,
            I => \N__24936\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__24936\,
            I => \nx.n1477\
        );

    \I__3732\ : CascadeMux
    port map (
            O => \N__24933\,
            I => \nx.n1509_cascade_\
        );

    \I__3731\ : InMux
    port map (
            O => \N__24930\,
            I => \N__24927\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__24927\,
            I => \nx.n16_adj_629\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__24924\,
            I => \nx.n18_adj_630_cascade_\
        );

    \I__3728\ : InMux
    port map (
            O => \N__24921\,
            I => \N__24918\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__24918\,
            I => \nx.n13_adj_631\
        );

    \I__3726\ : InMux
    port map (
            O => \N__24915\,
            I => \N__24912\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__24912\,
            I => \N__24909\
        );

    \I__3724\ : Odrv4
    port map (
            O => \N__24909\,
            I => \nx.n1469\
        );

    \I__3723\ : CascadeMux
    port map (
            O => \N__24906\,
            I => \nx.n1433_cascade_\
        );

    \I__3722\ : CascadeMux
    port map (
            O => \N__24903\,
            I => \N__24899\
        );

    \I__3721\ : InMux
    port map (
            O => \N__24902\,
            I => \N__24895\
        );

    \I__3720\ : InMux
    port map (
            O => \N__24899\,
            I => \N__24890\
        );

    \I__3719\ : InMux
    port map (
            O => \N__24898\,
            I => \N__24890\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__24895\,
            I => \nx.n1402\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__24890\,
            I => \nx.n1402\
        );

    \I__3716\ : CascadeMux
    port map (
            O => \N__24885\,
            I => \nx.n1501_cascade_\
        );

    \I__3715\ : InMux
    port map (
            O => \N__24882\,
            I => \N__24879\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__24879\,
            I => \nx.n9672\
        );

    \I__3713\ : InMux
    port map (
            O => \N__24876\,
            I => \N__24873\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__24873\,
            I => \N__24869\
        );

    \I__3711\ : InMux
    port map (
            O => \N__24872\,
            I => \N__24865\
        );

    \I__3710\ : Span4Mux_h
    port map (
            O => \N__24869\,
            I => \N__24862\
        );

    \I__3709\ : InMux
    port map (
            O => \N__24868\,
            I => \N__24859\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__24865\,
            I => \N__24856\
        );

    \I__3707\ : Odrv4
    port map (
            O => \N__24862\,
            I => timer_22
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__24859\,
            I => timer_22
        );

    \I__3705\ : Odrv12
    port map (
            O => \N__24856\,
            I => timer_22
        );

    \I__3704\ : InMux
    port map (
            O => \N__24849\,
            I => \nx.n10421\
        );

    \I__3703\ : CEMux
    port map (
            O => \N__24846\,
            I => \N__24841\
        );

    \I__3702\ : CEMux
    port map (
            O => \N__24845\,
            I => \N__24837\
        );

    \I__3701\ : CEMux
    port map (
            O => \N__24844\,
            I => \N__24834\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__24841\,
            I => \N__24831\
        );

    \I__3699\ : CEMux
    port map (
            O => \N__24840\,
            I => \N__24828\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__24837\,
            I => \N__24825\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__24834\,
            I => \N__24822\
        );

    \I__3696\ : Span4Mux_h
    port map (
            O => \N__24831\,
            I => \N__24817\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__24828\,
            I => \N__24817\
        );

    \I__3694\ : Span4Mux_v
    port map (
            O => \N__24825\,
            I => \N__24814\
        );

    \I__3693\ : Span4Mux_h
    port map (
            O => \N__24822\,
            I => \N__24811\
        );

    \I__3692\ : Span4Mux_v
    port map (
            O => \N__24817\,
            I => \N__24808\
        );

    \I__3691\ : Span4Mux_v
    port map (
            O => \N__24814\,
            I => \N__24805\
        );

    \I__3690\ : Span4Mux_v
    port map (
            O => \N__24811\,
            I => \N__24802\
        );

    \I__3689\ : Span4Mux_h
    port map (
            O => \N__24808\,
            I => \N__24799\
        );

    \I__3688\ : Span4Mux_v
    port map (
            O => \N__24805\,
            I => \N__24796\
        );

    \I__3687\ : Span4Mux_v
    port map (
            O => \N__24802\,
            I => \N__24793\
        );

    \I__3686\ : Span4Mux_v
    port map (
            O => \N__24799\,
            I => \N__24790\
        );

    \I__3685\ : Odrv4
    port map (
            O => \N__24796\,
            I => \nx.n7230\
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__24793\,
            I => \nx.n7230\
        );

    \I__3683\ : Odrv4
    port map (
            O => \N__24790\,
            I => \nx.n7230\
        );

    \I__3682\ : SRMux
    port map (
            O => \N__24783\,
            I => \N__24780\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__24780\,
            I => \N__24775\
        );

    \I__3680\ : SRMux
    port map (
            O => \N__24779\,
            I => \N__24772\
        );

    \I__3679\ : SRMux
    port map (
            O => \N__24778\,
            I => \N__24769\
        );

    \I__3678\ : Span4Mux_v
    port map (
            O => \N__24775\,
            I => \N__24765\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__24772\,
            I => \N__24760\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__24769\,
            I => \N__24760\
        );

    \I__3675\ : SRMux
    port map (
            O => \N__24768\,
            I => \N__24757\
        );

    \I__3674\ : Span4Mux_h
    port map (
            O => \N__24765\,
            I => \N__24750\
        );

    \I__3673\ : Span4Mux_v
    port map (
            O => \N__24760\,
            I => \N__24750\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__24757\,
            I => \N__24750\
        );

    \I__3671\ : Span4Mux_h
    port map (
            O => \N__24750\,
            I => \N__24747\
        );

    \I__3670\ : Span4Mux_v
    port map (
            O => \N__24747\,
            I => \N__24744\
        );

    \I__3669\ : Span4Mux_v
    port map (
            O => \N__24744\,
            I => \N__24741\
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__24741\,
            I => \nx.n7411\
        );

    \I__3667\ : InMux
    port map (
            O => \N__24738\,
            I => \N__24735\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__24735\,
            I => \N__24730\
        );

    \I__3665\ : CascadeMux
    port map (
            O => \N__24734\,
            I => \N__24727\
        );

    \I__3664\ : InMux
    port map (
            O => \N__24733\,
            I => \N__24724\
        );

    \I__3663\ : Span4Mux_h
    port map (
            O => \N__24730\,
            I => \N__24721\
        );

    \I__3662\ : InMux
    port map (
            O => \N__24727\,
            I => \N__24718\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__24724\,
            I => \N__24715\
        );

    \I__3660\ : Odrv4
    port map (
            O => \N__24721\,
            I => \nx.n1308\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__24718\,
            I => \nx.n1308\
        );

    \I__3658\ : Odrv4
    port map (
            O => \N__24715\,
            I => \nx.n1308\
        );

    \I__3657\ : CascadeMux
    port map (
            O => \N__24708\,
            I => \N__24705\
        );

    \I__3656\ : InMux
    port map (
            O => \N__24705\,
            I => \N__24702\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__24702\,
            I => \N__24699\
        );

    \I__3654\ : Odrv4
    port map (
            O => \N__24699\,
            I => \nx.n1375\
        );

    \I__3653\ : InMux
    port map (
            O => \N__24696\,
            I => \N__24693\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__24693\,
            I => \N__24690\
        );

    \I__3651\ : Odrv4
    port map (
            O => \N__24690\,
            I => \nx.n1373\
        );

    \I__3650\ : InMux
    port map (
            O => \N__24687\,
            I => \N__24684\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__24684\,
            I => \N__24680\
        );

    \I__3648\ : CascadeMux
    port map (
            O => \N__24683\,
            I => \N__24677\
        );

    \I__3647\ : Span4Mux_s2_v
    port map (
            O => \N__24680\,
            I => \N__24674\
        );

    \I__3646\ : InMux
    port map (
            O => \N__24677\,
            I => \N__24671\
        );

    \I__3645\ : Odrv4
    port map (
            O => \N__24674\,
            I => \nx.n1306\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__24671\,
            I => \nx.n1306\
        );

    \I__3643\ : InMux
    port map (
            O => \N__24666\,
            I => \N__24663\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__24663\,
            I => \N__24660\
        );

    \I__3641\ : Odrv4
    port map (
            O => \N__24660\,
            I => \nx.n1371\
        );

    \I__3640\ : CascadeMux
    port map (
            O => \N__24657\,
            I => \N__24654\
        );

    \I__3639\ : InMux
    port map (
            O => \N__24654\,
            I => \N__24649\
        );

    \I__3638\ : InMux
    port map (
            O => \N__24653\,
            I => \N__24646\
        );

    \I__3637\ : InMux
    port map (
            O => \N__24652\,
            I => \N__24643\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__24649\,
            I => \nx.n1304\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__24646\,
            I => \nx.n1304\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__24643\,
            I => \nx.n1304\
        );

    \I__3633\ : InMux
    port map (
            O => \N__24636\,
            I => \N__24632\
        );

    \I__3632\ : InMux
    port map (
            O => \N__24635\,
            I => \N__24628\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__24632\,
            I => \N__24625\
        );

    \I__3630\ : CascadeMux
    port map (
            O => \N__24631\,
            I => \N__24622\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__24628\,
            I => \N__24619\
        );

    \I__3628\ : Span4Mux_h
    port map (
            O => \N__24625\,
            I => \N__24616\
        );

    \I__3627\ : InMux
    port map (
            O => \N__24622\,
            I => \N__24613\
        );

    \I__3626\ : Span4Mux_h
    port map (
            O => \N__24619\,
            I => \N__24610\
        );

    \I__3625\ : Odrv4
    port map (
            O => \N__24616\,
            I => \nx.n1305\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__24613\,
            I => \nx.n1305\
        );

    \I__3623\ : Odrv4
    port map (
            O => \N__24610\,
            I => \nx.n1305\
        );

    \I__3622\ : CascadeMux
    port map (
            O => \N__24603\,
            I => \N__24600\
        );

    \I__3621\ : InMux
    port map (
            O => \N__24600\,
            I => \N__24597\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__24597\,
            I => \N__24594\
        );

    \I__3619\ : Odrv4
    port map (
            O => \N__24594\,
            I => \nx.n1372\
        );

    \I__3618\ : CascadeMux
    port map (
            O => \N__24591\,
            I => \N__24582\
        );

    \I__3617\ : InMux
    port map (
            O => \N__24590\,
            I => \N__24577\
        );

    \I__3616\ : InMux
    port map (
            O => \N__24589\,
            I => \N__24572\
        );

    \I__3615\ : InMux
    port map (
            O => \N__24588\,
            I => \N__24572\
        );

    \I__3614\ : InMux
    port map (
            O => \N__24587\,
            I => \N__24567\
        );

    \I__3613\ : InMux
    port map (
            O => \N__24586\,
            I => \N__24567\
        );

    \I__3612\ : InMux
    port map (
            O => \N__24585\,
            I => \N__24558\
        );

    \I__3611\ : InMux
    port map (
            O => \N__24582\,
            I => \N__24558\
        );

    \I__3610\ : InMux
    port map (
            O => \N__24581\,
            I => \N__24558\
        );

    \I__3609\ : InMux
    port map (
            O => \N__24580\,
            I => \N__24558\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__24577\,
            I => \N__24553\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__24572\,
            I => \N__24553\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__24567\,
            I => \nx.n1334\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__24558\,
            I => \nx.n1334\
        );

    \I__3604\ : Odrv4
    port map (
            O => \N__24553\,
            I => \nx.n1334\
        );

    \I__3603\ : CascadeMux
    port map (
            O => \N__24546\,
            I => \nx.n1404_cascade_\
        );

    \I__3602\ : InMux
    port map (
            O => \N__24543\,
            I => \N__24538\
        );

    \I__3601\ : InMux
    port map (
            O => \N__24542\,
            I => \N__24535\
        );

    \I__3600\ : InMux
    port map (
            O => \N__24541\,
            I => \N__24530\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__24538\,
            I => \N__24527\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__24535\,
            I => \N__24524\
        );

    \I__3597\ : InMux
    port map (
            O => \N__24534\,
            I => \N__24521\
        );

    \I__3596\ : InMux
    port map (
            O => \N__24533\,
            I => \N__24518\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__24530\,
            I => \N__24513\
        );

    \I__3594\ : Span4Mux_s3_h
    port map (
            O => \N__24527\,
            I => \N__24513\
        );

    \I__3593\ : Span4Mux_s3_h
    port map (
            O => \N__24524\,
            I => \N__24510\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__24521\,
            I => \nx.bit_ctr_23\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__24518\,
            I => \nx.bit_ctr_23\
        );

    \I__3590\ : Odrv4
    port map (
            O => \N__24513\,
            I => \nx.bit_ctr_23\
        );

    \I__3589\ : Odrv4
    port map (
            O => \N__24510\,
            I => \nx.bit_ctr_23\
        );

    \I__3588\ : InMux
    port map (
            O => \N__24501\,
            I => \N__24498\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__24498\,
            I => \N__24495\
        );

    \I__3586\ : Span4Mux_h
    port map (
            O => \N__24495\,
            I => \N__24492\
        );

    \I__3585\ : Odrv4
    port map (
            O => \N__24492\,
            I => \nx.n47_adj_706\
        );

    \I__3584\ : CascadeMux
    port map (
            O => \N__24489\,
            I => \N__24485\
        );

    \I__3583\ : InMux
    port map (
            O => \N__24488\,
            I => \N__24482\
        );

    \I__3582\ : InMux
    port map (
            O => \N__24485\,
            I => \N__24479\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__24482\,
            I => \nx.n1404\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__24479\,
            I => \nx.n1404\
        );

    \I__3579\ : InMux
    port map (
            O => \N__24474\,
            I => \N__24471\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__24471\,
            I => \nx.n1471\
        );

    \I__3577\ : InMux
    port map (
            O => \N__24468\,
            I => \nx.n10412\
        );

    \I__3576\ : InMux
    port map (
            O => \N__24465\,
            I => \nx.n10413\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__24462\,
            I => \N__24457\
        );

    \I__3574\ : InMux
    port map (
            O => \N__24461\,
            I => \N__24451\
        );

    \I__3573\ : InMux
    port map (
            O => \N__24460\,
            I => \N__24451\
        );

    \I__3572\ : InMux
    port map (
            O => \N__24457\,
            I => \N__24448\
        );

    \I__3571\ : InMux
    port map (
            O => \N__24456\,
            I => \N__24445\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__24451\,
            I => \N__24441\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__24448\,
            I => \N__24436\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__24445\,
            I => \N__24436\
        );

    \I__3567\ : InMux
    port map (
            O => \N__24444\,
            I => \N__24433\
        );

    \I__3566\ : Span4Mux_s1_h
    port map (
            O => \N__24441\,
            I => \N__24428\
        );

    \I__3565\ : Span4Mux_v
    port map (
            O => \N__24436\,
            I => \N__24428\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__24433\,
            I => \nx.bit_ctr_24\
        );

    \I__3563\ : Odrv4
    port map (
            O => \N__24428\,
            I => \nx.bit_ctr_24\
        );

    \I__3562\ : InMux
    port map (
            O => \N__24423\,
            I => \bfn_4_30_0_\
        );

    \I__3561\ : InMux
    port map (
            O => \N__24420\,
            I => \nx.n10415\
        );

    \I__3560\ : InMux
    port map (
            O => \N__24417\,
            I => \nx.n10416\
        );

    \I__3559\ : InMux
    port map (
            O => \N__24414\,
            I => \nx.n10417\
        );

    \I__3558\ : InMux
    port map (
            O => \N__24411\,
            I => \nx.n10418\
        );

    \I__3557\ : InMux
    port map (
            O => \N__24408\,
            I => \nx.n10419\
        );

    \I__3556\ : InMux
    port map (
            O => \N__24405\,
            I => \nx.n10420\
        );

    \I__3555\ : InMux
    port map (
            O => \N__24402\,
            I => \nx.n10403\
        );

    \I__3554\ : InMux
    port map (
            O => \N__24399\,
            I => \nx.n10404\
        );

    \I__3553\ : InMux
    port map (
            O => \N__24396\,
            I => \nx.n10405\
        );

    \I__3552\ : InMux
    port map (
            O => \N__24393\,
            I => \bfn_4_29_0_\
        );

    \I__3551\ : InMux
    port map (
            O => \N__24390\,
            I => \nx.n10407\
        );

    \I__3550\ : InMux
    port map (
            O => \N__24387\,
            I => \nx.n10408\
        );

    \I__3549\ : InMux
    port map (
            O => \N__24384\,
            I => \nx.n10409\
        );

    \I__3548\ : InMux
    port map (
            O => \N__24381\,
            I => \nx.n10410\
        );

    \I__3547\ : InMux
    port map (
            O => \N__24378\,
            I => \nx.n10411\
        );

    \I__3546\ : InMux
    port map (
            O => \N__24375\,
            I => \N__24371\
        );

    \I__3545\ : InMux
    port map (
            O => \N__24374\,
            I => \N__24366\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__24371\,
            I => \N__24363\
        );

    \I__3543\ : InMux
    port map (
            O => \N__24370\,
            I => \N__24360\
        );

    \I__3542\ : InMux
    port map (
            O => \N__24369\,
            I => \N__24357\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__24366\,
            I => \N__24353\
        );

    \I__3540\ : Span4Mux_v
    port map (
            O => \N__24363\,
            I => \N__24350\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__24360\,
            I => \N__24345\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__24357\,
            I => \N__24345\
        );

    \I__3537\ : InMux
    port map (
            O => \N__24356\,
            I => \N__24342\
        );

    \I__3536\ : Span4Mux_v
    port map (
            O => \N__24353\,
            I => \N__24335\
        );

    \I__3535\ : Span4Mux_s1_h
    port map (
            O => \N__24350\,
            I => \N__24335\
        );

    \I__3534\ : Span4Mux_v
    port map (
            O => \N__24345\,
            I => \N__24335\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__24342\,
            I => \nx.bit_ctr_4\
        );

    \I__3532\ : Odrv4
    port map (
            O => \N__24335\,
            I => \nx.bit_ctr_4\
        );

    \I__3531\ : InMux
    port map (
            O => \N__24330\,
            I => \nx.n10394\
        );

    \I__3530\ : InMux
    port map (
            O => \N__24327\,
            I => \nx.n10395\
        );

    \I__3529\ : InMux
    port map (
            O => \N__24324\,
            I => \nx.n10396\
        );

    \I__3528\ : InMux
    port map (
            O => \N__24321\,
            I => \nx.n10397\
        );

    \I__3527\ : InMux
    port map (
            O => \N__24318\,
            I => \bfn_4_28_0_\
        );

    \I__3526\ : InMux
    port map (
            O => \N__24315\,
            I => \nx.n10399\
        );

    \I__3525\ : InMux
    port map (
            O => \N__24312\,
            I => \nx.n10400\
        );

    \I__3524\ : InMux
    port map (
            O => \N__24309\,
            I => \nx.n10401\
        );

    \I__3523\ : InMux
    port map (
            O => \N__24306\,
            I => \nx.n10402\
        );

    \I__3522\ : InMux
    port map (
            O => \N__24303\,
            I => \N__24300\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__24300\,
            I => \N__24297\
        );

    \I__3520\ : Span4Mux_h
    port map (
            O => \N__24297\,
            I => \N__24294\
        );

    \I__3519\ : Odrv4
    port map (
            O => \N__24294\,
            I => \nx.n3157\
        );

    \I__3518\ : CascadeMux
    port map (
            O => \N__24291\,
            I => \nx.n12361_cascade_\
        );

    \I__3517\ : CascadeMux
    port map (
            O => \N__24288\,
            I => \N__24285\
        );

    \I__3516\ : InMux
    port map (
            O => \N__24285\,
            I => \N__24282\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__24282\,
            I => \N__24278\
        );

    \I__3514\ : InMux
    port map (
            O => \N__24281\,
            I => \N__24274\
        );

    \I__3513\ : Span4Mux_v
    port map (
            O => \N__24278\,
            I => \N__24271\
        );

    \I__3512\ : InMux
    port map (
            O => \N__24277\,
            I => \N__24268\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__24274\,
            I => \nx.n3090\
        );

    \I__3510\ : Odrv4
    port map (
            O => \N__24271\,
            I => \nx.n3090\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__24268\,
            I => \nx.n3090\
        );

    \I__3508\ : InMux
    port map (
            O => \N__24261\,
            I => \N__24258\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__24258\,
            I => \N__24255\
        );

    \I__3506\ : Span4Mux_h
    port map (
            O => \N__24255\,
            I => \N__24252\
        );

    \I__3505\ : Odrv4
    port map (
            O => \N__24252\,
            I => \nx.n3156\
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__24249\,
            I => \nx.n12363_cascade_\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__24246\,
            I => \N__24243\
        );

    \I__3502\ : InMux
    port map (
            O => \N__24243\,
            I => \N__24231\
        );

    \I__3501\ : InMux
    port map (
            O => \N__24242\,
            I => \N__24218\
        );

    \I__3500\ : InMux
    port map (
            O => \N__24241\,
            I => \N__24218\
        );

    \I__3499\ : InMux
    port map (
            O => \N__24240\,
            I => \N__24218\
        );

    \I__3498\ : InMux
    port map (
            O => \N__24239\,
            I => \N__24218\
        );

    \I__3497\ : InMux
    port map (
            O => \N__24238\,
            I => \N__24218\
        );

    \I__3496\ : InMux
    port map (
            O => \N__24237\,
            I => \N__24218\
        );

    \I__3495\ : CascadeMux
    port map (
            O => \N__24236\,
            I => \N__24215\
        );

    \I__3494\ : CascadeMux
    port map (
            O => \N__24235\,
            I => \N__24210\
        );

    \I__3493\ : InMux
    port map (
            O => \N__24234\,
            I => \N__24204\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__24231\,
            I => \N__24201\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__24218\,
            I => \N__24198\
        );

    \I__3490\ : InMux
    port map (
            O => \N__24215\,
            I => \N__24195\
        );

    \I__3489\ : InMux
    port map (
            O => \N__24214\,
            I => \N__24190\
        );

    \I__3488\ : InMux
    port map (
            O => \N__24213\,
            I => \N__24190\
        );

    \I__3487\ : InMux
    port map (
            O => \N__24210\,
            I => \N__24185\
        );

    \I__3486\ : InMux
    port map (
            O => \N__24209\,
            I => \N__24185\
        );

    \I__3485\ : CascadeMux
    port map (
            O => \N__24208\,
            I => \N__24182\
        );

    \I__3484\ : CascadeMux
    port map (
            O => \N__24207\,
            I => \N__24178\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__24204\,
            I => \N__24164\
        );

    \I__3482\ : Span4Mux_v
    port map (
            O => \N__24201\,
            I => \N__24157\
        );

    \I__3481\ : Span4Mux_v
    port map (
            O => \N__24198\,
            I => \N__24157\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__24195\,
            I => \N__24157\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__24190\,
            I => \N__24152\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__24185\,
            I => \N__24152\
        );

    \I__3477\ : InMux
    port map (
            O => \N__24182\,
            I => \N__24137\
        );

    \I__3476\ : InMux
    port map (
            O => \N__24181\,
            I => \N__24137\
        );

    \I__3475\ : InMux
    port map (
            O => \N__24178\,
            I => \N__24137\
        );

    \I__3474\ : InMux
    port map (
            O => \N__24177\,
            I => \N__24137\
        );

    \I__3473\ : InMux
    port map (
            O => \N__24176\,
            I => \N__24137\
        );

    \I__3472\ : InMux
    port map (
            O => \N__24175\,
            I => \N__24137\
        );

    \I__3471\ : InMux
    port map (
            O => \N__24174\,
            I => \N__24137\
        );

    \I__3470\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24132\
        );

    \I__3469\ : InMux
    port map (
            O => \N__24172\,
            I => \N__24132\
        );

    \I__3468\ : InMux
    port map (
            O => \N__24171\,
            I => \N__24127\
        );

    \I__3467\ : InMux
    port map (
            O => \N__24170\,
            I => \N__24127\
        );

    \I__3466\ : InMux
    port map (
            O => \N__24169\,
            I => \N__24120\
        );

    \I__3465\ : InMux
    port map (
            O => \N__24168\,
            I => \N__24120\
        );

    \I__3464\ : InMux
    port map (
            O => \N__24167\,
            I => \N__24120\
        );

    \I__3463\ : Odrv4
    port map (
            O => \N__24164\,
            I => \nx.n3116\
        );

    \I__3462\ : Odrv4
    port map (
            O => \N__24157\,
            I => \nx.n3116\
        );

    \I__3461\ : Odrv4
    port map (
            O => \N__24152\,
            I => \nx.n3116\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__24137\,
            I => \nx.n3116\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__24132\,
            I => \nx.n3116\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__24127\,
            I => \nx.n3116\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__24120\,
            I => \nx.n3116\
        );

    \I__3456\ : InMux
    port map (
            O => \N__24105\,
            I => \N__24102\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__24102\,
            I => \N__24098\
        );

    \I__3454\ : InMux
    port map (
            O => \N__24101\,
            I => \N__24095\
        );

    \I__3453\ : Span4Mux_v
    port map (
            O => \N__24098\,
            I => \N__24092\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__24095\,
            I => \nx.n3088\
        );

    \I__3451\ : Odrv4
    port map (
            O => \N__24092\,
            I => \nx.n3088\
        );

    \I__3450\ : CascadeMux
    port map (
            O => \N__24087\,
            I => \nx.n12365_cascade_\
        );

    \I__3449\ : InMux
    port map (
            O => \N__24084\,
            I => \N__24081\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__24081\,
            I => \N__24078\
        );

    \I__3447\ : Span4Mux_h
    port map (
            O => \N__24078\,
            I => \N__24075\
        );

    \I__3446\ : Odrv4
    port map (
            O => \N__24075\,
            I => \nx.n3155\
        );

    \I__3445\ : InMux
    port map (
            O => \N__24072\,
            I => \N__24069\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__24069\,
            I => \N__24066\
        );

    \I__3443\ : Span4Mux_s1_h
    port map (
            O => \N__24066\,
            I => \N__24063\
        );

    \I__3442\ : Span4Mux_v
    port map (
            O => \N__24063\,
            I => \N__24060\
        );

    \I__3441\ : Odrv4
    port map (
            O => \N__24060\,
            I => \nx.n12367\
        );

    \I__3440\ : CascadeMux
    port map (
            O => \N__24057\,
            I => \N__24054\
        );

    \I__3439\ : InMux
    port map (
            O => \N__24054\,
            I => \N__24050\
        );

    \I__3438\ : InMux
    port map (
            O => \N__24053\,
            I => \N__24047\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__24050\,
            I => \N__24044\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__24047\,
            I => \N__24040\
        );

    \I__3435\ : Span4Mux_v
    port map (
            O => \N__24044\,
            I => \N__24037\
        );

    \I__3434\ : InMux
    port map (
            O => \N__24043\,
            I => \N__24034\
        );

    \I__3433\ : Odrv4
    port map (
            O => \N__24040\,
            I => \nx.n2990\
        );

    \I__3432\ : Odrv4
    port map (
            O => \N__24037\,
            I => \nx.n2990\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__24034\,
            I => \nx.n2990\
        );

    \I__3430\ : CascadeMux
    port map (
            O => \N__24027\,
            I => \N__24024\
        );

    \I__3429\ : InMux
    port map (
            O => \N__24024\,
            I => \N__24021\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__24021\,
            I => \N__24018\
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__24018\,
            I => \nx.n3057\
        );

    \I__3426\ : InMux
    port map (
            O => \N__24015\,
            I => \N__24011\
        );

    \I__3425\ : InMux
    port map (
            O => \N__24014\,
            I => \N__24008\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__24011\,
            I => \N__24005\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__24008\,
            I => \N__23999\
        );

    \I__3422\ : Span4Mux_s3_h
    port map (
            O => \N__24005\,
            I => \N__23999\
        );

    \I__3421\ : InMux
    port map (
            O => \N__24004\,
            I => \N__23996\
        );

    \I__3420\ : Odrv4
    port map (
            O => \N__23999\,
            I => \nx.n3089\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__23996\,
            I => \nx.n3089\
        );

    \I__3418\ : InMux
    port map (
            O => \N__23991\,
            I => \N__23986\
        );

    \I__3417\ : InMux
    port map (
            O => \N__23990\,
            I => \N__23983\
        );

    \I__3416\ : InMux
    port map (
            O => \N__23989\,
            I => \N__23980\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__23986\,
            I => \N__23976\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__23983\,
            I => \N__23971\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__23980\,
            I => \N__23971\
        );

    \I__3412\ : InMux
    port map (
            O => \N__23979\,
            I => \N__23968\
        );

    \I__3411\ : Span4Mux_v
    port map (
            O => \N__23976\,
            I => \N__23963\
        );

    \I__3410\ : Span4Mux_v
    port map (
            O => \N__23971\,
            I => \N__23963\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__23968\,
            I => \N__23960\
        );

    \I__3408\ : Span4Mux_v
    port map (
            O => \N__23963\,
            I => \N__23956\
        );

    \I__3407\ : Span12Mux_v
    port map (
            O => \N__23960\,
            I => \N__23953\
        );

    \I__3406\ : InMux
    port map (
            O => \N__23959\,
            I => \N__23950\
        );

    \I__3405\ : Odrv4
    port map (
            O => \N__23956\,
            I => \nx.bit_ctr_0\
        );

    \I__3404\ : Odrv12
    port map (
            O => \N__23953\,
            I => \nx.bit_ctr_0\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__23950\,
            I => \nx.bit_ctr_0\
        );

    \I__3402\ : InMux
    port map (
            O => \N__23943\,
            I => \bfn_4_27_0_\
        );

    \I__3401\ : CascadeMux
    port map (
            O => \N__23940\,
            I => \N__23937\
        );

    \I__3400\ : InMux
    port map (
            O => \N__23937\,
            I => \N__23934\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__23934\,
            I => \N__23931\
        );

    \I__3398\ : Span4Mux_s3_h
    port map (
            O => \N__23931\,
            I => \N__23928\
        );

    \I__3397\ : Span4Mux_v
    port map (
            O => \N__23928\,
            I => \N__23924\
        );

    \I__3396\ : InMux
    port map (
            O => \N__23927\,
            I => \N__23921\
        );

    \I__3395\ : Odrv4
    port map (
            O => \N__23924\,
            I => \nx.bit_ctr_1\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__23921\,
            I => \nx.bit_ctr_1\
        );

    \I__3393\ : InMux
    port map (
            O => \N__23916\,
            I => \nx.n10391\
        );

    \I__3392\ : InMux
    port map (
            O => \N__23913\,
            I => \N__23910\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__23910\,
            I => \N__23907\
        );

    \I__3390\ : Span4Mux_v
    port map (
            O => \N__23907\,
            I => \N__23904\
        );

    \I__3389\ : Span4Mux_v
    port map (
            O => \N__23904\,
            I => \N__23900\
        );

    \I__3388\ : InMux
    port map (
            O => \N__23903\,
            I => \N__23897\
        );

    \I__3387\ : Odrv4
    port map (
            O => \N__23900\,
            I => \nx.bit_ctr_2\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__23897\,
            I => \nx.bit_ctr_2\
        );

    \I__3385\ : InMux
    port map (
            O => \N__23892\,
            I => \nx.n10392\
        );

    \I__3384\ : InMux
    port map (
            O => \N__23889\,
            I => \N__23882\
        );

    \I__3383\ : InMux
    port map (
            O => \N__23888\,
            I => \N__23882\
        );

    \I__3382\ : InMux
    port map (
            O => \N__23887\,
            I => \N__23879\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__23882\,
            I => \N__23874\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__23879\,
            I => \N__23871\
        );

    \I__3379\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23868\
        );

    \I__3378\ : InMux
    port map (
            O => \N__23877\,
            I => \N__23865\
        );

    \I__3377\ : Span4Mux_v
    port map (
            O => \N__23874\,
            I => \N__23858\
        );

    \I__3376\ : Span4Mux_v
    port map (
            O => \N__23871\,
            I => \N__23858\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__23868\,
            I => \N__23858\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__23865\,
            I => \N__23853\
        );

    \I__3373\ : Span4Mux_v
    port map (
            O => \N__23858\,
            I => \N__23853\
        );

    \I__3372\ : Odrv4
    port map (
            O => \N__23853\,
            I => \nx.bit_ctr_3\
        );

    \I__3371\ : InMux
    port map (
            O => \N__23850\,
            I => \nx.n10393\
        );

    \I__3370\ : CascadeMux
    port map (
            O => \N__23847\,
            I => \N__23843\
        );

    \I__3369\ : CascadeMux
    port map (
            O => \N__23846\,
            I => \N__23840\
        );

    \I__3368\ : InMux
    port map (
            O => \N__23843\,
            I => \N__23837\
        );

    \I__3367\ : InMux
    port map (
            O => \N__23840\,
            I => \N__23834\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__23837\,
            I => \N__23829\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__23834\,
            I => \N__23829\
        );

    \I__3364\ : Span4Mux_v
    port map (
            O => \N__23829\,
            I => \N__23825\
        );

    \I__3363\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23822\
        );

    \I__3362\ : Odrv4
    port map (
            O => \N__23825\,
            I => \nx.n2992\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__23822\,
            I => \nx.n2992\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__23817\,
            I => \N__23814\
        );

    \I__3359\ : InMux
    port map (
            O => \N__23814\,
            I => \N__23810\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__23813\,
            I => \N__23807\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__23810\,
            I => \N__23804\
        );

    \I__3356\ : InMux
    port map (
            O => \N__23807\,
            I => \N__23800\
        );

    \I__3355\ : Span4Mux_v
    port map (
            O => \N__23804\,
            I => \N__23797\
        );

    \I__3354\ : InMux
    port map (
            O => \N__23803\,
            I => \N__23794\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__23800\,
            I => \nx.n2989\
        );

    \I__3352\ : Odrv4
    port map (
            O => \N__23797\,
            I => \nx.n2989\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__23794\,
            I => \nx.n2989\
        );

    \I__3350\ : InMux
    port map (
            O => \N__23787\,
            I => \N__23784\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__23784\,
            I => \N__23781\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__23781\,
            I => \nx.n3056\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__23778\,
            I => \N__23773\
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__23777\,
            I => \N__23770\
        );

    \I__3345\ : InMux
    port map (
            O => \N__23776\,
            I => \N__23767\
        );

    \I__3344\ : InMux
    port map (
            O => \N__23773\,
            I => \N__23764\
        );

    \I__3343\ : InMux
    port map (
            O => \N__23770\,
            I => \N__23761\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__23767\,
            I => \N__23758\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__23764\,
            I => \nx.n3104\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__23761\,
            I => \nx.n3104\
        );

    \I__3339\ : Odrv4
    port map (
            O => \N__23758\,
            I => \nx.n3104\
        );

    \I__3338\ : CascadeMux
    port map (
            O => \N__23751\,
            I => \nx.n3088_cascade_\
        );

    \I__3337\ : InMux
    port map (
            O => \N__23748\,
            I => \N__23745\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__23745\,
            I => \N__23742\
        );

    \I__3335\ : Odrv4
    port map (
            O => \N__23742\,
            I => \nx.n44_adj_690\
        );

    \I__3334\ : InMux
    port map (
            O => \N__23739\,
            I => \N__23736\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__23736\,
            I => \N__23733\
        );

    \I__3332\ : Odrv4
    port map (
            O => \N__23733\,
            I => \nx.n3061\
        );

    \I__3331\ : CascadeMux
    port map (
            O => \N__23730\,
            I => \N__23726\
        );

    \I__3330\ : InMux
    port map (
            O => \N__23729\,
            I => \N__23723\
        );

    \I__3329\ : InMux
    port map (
            O => \N__23726\,
            I => \N__23720\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__23723\,
            I => \N__23717\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__23720\,
            I => \N__23712\
        );

    \I__3326\ : Span4Mux_v
    port map (
            O => \N__23717\,
            I => \N__23712\
        );

    \I__3325\ : Odrv4
    port map (
            O => \N__23712\,
            I => \nx.n2994\
        );

    \I__3324\ : CascadeMux
    port map (
            O => \N__23709\,
            I => \N__23706\
        );

    \I__3323\ : InMux
    port map (
            O => \N__23706\,
            I => \N__23702\
        );

    \I__3322\ : InMux
    port map (
            O => \N__23705\,
            I => \N__23699\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__23702\,
            I => \N__23696\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__23699\,
            I => \N__23690\
        );

    \I__3319\ : Span4Mux_v
    port map (
            O => \N__23696\,
            I => \N__23690\
        );

    \I__3318\ : InMux
    port map (
            O => \N__23695\,
            I => \N__23687\
        );

    \I__3317\ : Odrv4
    port map (
            O => \N__23690\,
            I => \nx.n2991\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__23687\,
            I => \nx.n2991\
        );

    \I__3315\ : InMux
    port map (
            O => \N__23682\,
            I => \N__23679\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__23679\,
            I => \N__23676\
        );

    \I__3313\ : Odrv4
    port map (
            O => \N__23676\,
            I => \nx.n3058\
        );

    \I__3312\ : InMux
    port map (
            O => \N__23673\,
            I => \N__23670\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__23670\,
            I => \N__23667\
        );

    \I__3310\ : Span4Mux_h
    port map (
            O => \N__23667\,
            I => \N__23664\
        );

    \I__3309\ : Odrv4
    port map (
            O => \N__23664\,
            I => \nx.n3161\
        );

    \I__3308\ : InMux
    port map (
            O => \N__23661\,
            I => \N__23658\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__23658\,
            I => \N__23655\
        );

    \I__3306\ : Odrv4
    port map (
            O => \N__23655\,
            I => \nx.n12353\
        );

    \I__3305\ : CascadeMux
    port map (
            O => \N__23652\,
            I => \N__23649\
        );

    \I__3304\ : InMux
    port map (
            O => \N__23649\,
            I => \N__23646\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__23646\,
            I => \N__23643\
        );

    \I__3302\ : Span4Mux_h
    port map (
            O => \N__23643\,
            I => \N__23640\
        );

    \I__3301\ : Odrv4
    port map (
            O => \N__23640\,
            I => \nx.n3160\
        );

    \I__3300\ : InMux
    port map (
            O => \N__23637\,
            I => \N__23634\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__23634\,
            I => \nx.n12355\
        );

    \I__3298\ : CascadeMux
    port map (
            O => \N__23631\,
            I => \nx.n12357_cascade_\
        );

    \I__3297\ : InMux
    port map (
            O => \N__23628\,
            I => \N__23625\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__23625\,
            I => \N__23622\
        );

    \I__3295\ : Span4Mux_v
    port map (
            O => \N__23622\,
            I => \N__23619\
        );

    \I__3294\ : Odrv4
    port map (
            O => \N__23619\,
            I => \nx.n3159\
        );

    \I__3293\ : InMux
    port map (
            O => \N__23616\,
            I => \N__23613\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__23613\,
            I => \N__23610\
        );

    \I__3291\ : Span4Mux_v
    port map (
            O => \N__23610\,
            I => \N__23607\
        );

    \I__3290\ : Odrv4
    port map (
            O => \N__23607\,
            I => \nx.n3158\
        );

    \I__3289\ : CascadeMux
    port map (
            O => \N__23604\,
            I => \nx.n12359_cascade_\
        );

    \I__3288\ : CascadeMux
    port map (
            O => \N__23601\,
            I => \N__23596\
        );

    \I__3287\ : InMux
    port map (
            O => \N__23600\,
            I => \N__23591\
        );

    \I__3286\ : InMux
    port map (
            O => \N__23599\,
            I => \N__23591\
        );

    \I__3285\ : InMux
    port map (
            O => \N__23596\,
            I => \N__23588\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__23591\,
            I => \N__23585\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__23588\,
            I => \N__23582\
        );

    \I__3282\ : Odrv4
    port map (
            O => \N__23585\,
            I => \nx.n3004\
        );

    \I__3281\ : Odrv4
    port map (
            O => \N__23582\,
            I => \nx.n3004\
        );

    \I__3280\ : CascadeMux
    port map (
            O => \N__23577\,
            I => \N__23573\
        );

    \I__3279\ : InMux
    port map (
            O => \N__23576\,
            I => \N__23570\
        );

    \I__3278\ : InMux
    port map (
            O => \N__23573\,
            I => \N__23567\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__23570\,
            I => \N__23564\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__23567\,
            I => \N__23561\
        );

    \I__3275\ : Span4Mux_s3_h
    port map (
            O => \N__23564\,
            I => \N__23558\
        );

    \I__3274\ : Span4Mux_v
    port map (
            O => \N__23561\,
            I => \N__23555\
        );

    \I__3273\ : Odrv4
    port map (
            O => \N__23558\,
            I => \nx.n2988\
        );

    \I__3272\ : Odrv4
    port map (
            O => \N__23555\,
            I => \nx.n2988\
        );

    \I__3271\ : CascadeMux
    port map (
            O => \N__23550\,
            I => \nx.n2988_cascade_\
        );

    \I__3270\ : InMux
    port map (
            O => \N__23547\,
            I => \N__23544\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__23544\,
            I => \N__23541\
        );

    \I__3268\ : Odrv4
    port map (
            O => \N__23541\,
            I => \nx.n41_adj_686\
        );

    \I__3267\ : CascadeMux
    port map (
            O => \N__23538\,
            I => \nx.n2994_cascade_\
        );

    \I__3266\ : CascadeMux
    port map (
            O => \N__23535\,
            I => \N__23531\
        );

    \I__3265\ : CascadeMux
    port map (
            O => \N__23534\,
            I => \N__23528\
        );

    \I__3264\ : InMux
    port map (
            O => \N__23531\,
            I => \N__23525\
        );

    \I__3263\ : InMux
    port map (
            O => \N__23528\,
            I => \N__23522\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__23525\,
            I => \N__23518\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__23522\,
            I => \N__23515\
        );

    \I__3260\ : InMux
    port map (
            O => \N__23521\,
            I => \N__23512\
        );

    \I__3259\ : Span4Mux_v
    port map (
            O => \N__23518\,
            I => \N__23509\
        );

    \I__3258\ : Odrv4
    port map (
            O => \N__23515\,
            I => \nx.n3002\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__23512\,
            I => \nx.n3002\
        );

    \I__3256\ : Odrv4
    port map (
            O => \N__23509\,
            I => \nx.n3002\
        );

    \I__3255\ : InMux
    port map (
            O => \N__23502\,
            I => \N__23499\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__23499\,
            I => \N__23496\
        );

    \I__3253\ : Odrv4
    port map (
            O => \N__23496\,
            I => \nx.n42_adj_684\
        );

    \I__3252\ : InMux
    port map (
            O => \N__23493\,
            I => \N__23489\
        );

    \I__3251\ : InMux
    port map (
            O => \N__23492\,
            I => \N__23486\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__23489\,
            I => \N__23482\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__23486\,
            I => \N__23479\
        );

    \I__3248\ : CascadeMux
    port map (
            O => \N__23485\,
            I => \N__23476\
        );

    \I__3247\ : Span4Mux_s3_h
    port map (
            O => \N__23482\,
            I => \N__23471\
        );

    \I__3246\ : Span4Mux_h
    port map (
            O => \N__23479\,
            I => \N__23471\
        );

    \I__3245\ : InMux
    port map (
            O => \N__23476\,
            I => \N__23468\
        );

    \I__3244\ : Odrv4
    port map (
            O => \N__23471\,
            I => \nx.n3009\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__23468\,
            I => \nx.n3009\
        );

    \I__3242\ : CascadeMux
    port map (
            O => \N__23463\,
            I => \nx.n2985_cascade_\
        );

    \I__3241\ : CascadeMux
    port map (
            O => \N__23460\,
            I => \N__23457\
        );

    \I__3240\ : InMux
    port map (
            O => \N__23457\,
            I => \N__23453\
        );

    \I__3239\ : InMux
    port map (
            O => \N__23456\,
            I => \N__23450\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__23453\,
            I => \N__23447\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__23450\,
            I => \N__23444\
        );

    \I__3236\ : Span4Mux_s3_h
    port map (
            O => \N__23447\,
            I => \N__23440\
        );

    \I__3235\ : Sp12to4
    port map (
            O => \N__23444\,
            I => \N__23437\
        );

    \I__3234\ : InMux
    port map (
            O => \N__23443\,
            I => \N__23434\
        );

    \I__3233\ : Odrv4
    port map (
            O => \N__23440\,
            I => \nx.n2986\
        );

    \I__3232\ : Odrv12
    port map (
            O => \N__23437\,
            I => \nx.n2986\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__23434\,
            I => \nx.n2986\
        );

    \I__3230\ : InMux
    port map (
            O => \N__23427\,
            I => \N__23424\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__23424\,
            I => \N__23421\
        );

    \I__3228\ : Span4Mux_s3_h
    port map (
            O => \N__23421\,
            I => \N__23418\
        );

    \I__3227\ : Odrv4
    port map (
            O => \N__23418\,
            I => \nx.n40_adj_683\
        );

    \I__3226\ : CascadeMux
    port map (
            O => \N__23415\,
            I => \N__23412\
        );

    \I__3225\ : InMux
    port map (
            O => \N__23412\,
            I => \N__23409\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__23409\,
            I => \N__23406\
        );

    \I__3223\ : Odrv4
    port map (
            O => \N__23406\,
            I => \nx.n43_adj_677\
        );

    \I__3222\ : InMux
    port map (
            O => \N__23403\,
            I => \N__23400\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__23400\,
            I => \nx.n40_adj_678\
        );

    \I__3220\ : CascadeMux
    port map (
            O => \N__23397\,
            I => \nx.n47_cascade_\
        );

    \I__3219\ : CascadeMux
    port map (
            O => \N__23394\,
            I => \nx.n2918_cascade_\
        );

    \I__3218\ : CascadeMux
    port map (
            O => \N__23391\,
            I => \N__23387\
        );

    \I__3217\ : InMux
    port map (
            O => \N__23390\,
            I => \N__23383\
        );

    \I__3216\ : InMux
    port map (
            O => \N__23387\,
            I => \N__23380\
        );

    \I__3215\ : InMux
    port map (
            O => \N__23386\,
            I => \N__23377\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__23383\,
            I => \N__23372\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__23380\,
            I => \N__23372\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__23377\,
            I => \N__23369\
        );

    \I__3211\ : Span4Mux_v
    port map (
            O => \N__23372\,
            I => \N__23366\
        );

    \I__3210\ : Odrv4
    port map (
            O => \N__23369\,
            I => \nx.n3000\
        );

    \I__3209\ : Odrv4
    port map (
            O => \N__23366\,
            I => \nx.n3000\
        );

    \I__3208\ : InMux
    port map (
            O => \N__23361\,
            I => \N__23358\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__23358\,
            I => \nx.n38_adj_676\
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__23355\,
            I => \N__23351\
        );

    \I__3205\ : CascadeMux
    port map (
            O => \N__23354\,
            I => \N__23348\
        );

    \I__3204\ : InMux
    port map (
            O => \N__23351\,
            I => \N__23344\
        );

    \I__3203\ : InMux
    port map (
            O => \N__23348\,
            I => \N__23341\
        );

    \I__3202\ : InMux
    port map (
            O => \N__23347\,
            I => \N__23338\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__23344\,
            I => \N__23335\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__23341\,
            I => \N__23332\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__23338\,
            I => \N__23329\
        );

    \I__3198\ : Span12Mux_s3_h
    port map (
            O => \N__23335\,
            I => \N__23326\
        );

    \I__3197\ : Odrv4
    port map (
            O => \N__23332\,
            I => \nx.n2996\
        );

    \I__3196\ : Odrv4
    port map (
            O => \N__23329\,
            I => \nx.n2996\
        );

    \I__3195\ : Odrv12
    port map (
            O => \N__23326\,
            I => \nx.n2996\
        );

    \I__3194\ : InMux
    port map (
            O => \N__23319\,
            I => \N__23315\
        );

    \I__3193\ : CascadeMux
    port map (
            O => \N__23318\,
            I => \N__23312\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__23315\,
            I => \N__23308\
        );

    \I__3191\ : InMux
    port map (
            O => \N__23312\,
            I => \N__23305\
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__23311\,
            I => \N__23302\
        );

    \I__3189\ : Span4Mux_s3_h
    port map (
            O => \N__23308\,
            I => \N__23297\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__23305\,
            I => \N__23297\
        );

    \I__3187\ : InMux
    port map (
            O => \N__23302\,
            I => \N__23294\
        );

    \I__3186\ : Span4Mux_v
    port map (
            O => \N__23297\,
            I => \N__23291\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__23294\,
            I => \N__23288\
        );

    \I__3184\ : Odrv4
    port map (
            O => \N__23291\,
            I => \nx.n2997\
        );

    \I__3183\ : Odrv4
    port map (
            O => \N__23288\,
            I => \nx.n2997\
        );

    \I__3182\ : CascadeMux
    port map (
            O => \N__23283\,
            I => \N__23279\
        );

    \I__3181\ : CascadeMux
    port map (
            O => \N__23282\,
            I => \N__23276\
        );

    \I__3180\ : InMux
    port map (
            O => \N__23279\,
            I => \N__23273\
        );

    \I__3179\ : InMux
    port map (
            O => \N__23276\,
            I => \N__23270\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__23273\,
            I => \N__23267\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__23270\,
            I => \N__23264\
        );

    \I__3176\ : Span4Mux_h
    port map (
            O => \N__23267\,
            I => \N__23260\
        );

    \I__3175\ : Span4Mux_v
    port map (
            O => \N__23264\,
            I => \N__23257\
        );

    \I__3174\ : InMux
    port map (
            O => \N__23263\,
            I => \N__23254\
        );

    \I__3173\ : Odrv4
    port map (
            O => \N__23260\,
            I => \nx.n2987\
        );

    \I__3172\ : Odrv4
    port map (
            O => \N__23257\,
            I => \nx.n2987\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__23254\,
            I => \nx.n2987\
        );

    \I__3170\ : CascadeMux
    port map (
            O => \N__23247\,
            I => \N__23243\
        );

    \I__3169\ : InMux
    port map (
            O => \N__23246\,
            I => \N__23240\
        );

    \I__3168\ : InMux
    port map (
            O => \N__23243\,
            I => \N__23237\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__23240\,
            I => \N__23234\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__23237\,
            I => \N__23230\
        );

    \I__3165\ : Span12Mux_s3_h
    port map (
            O => \N__23234\,
            I => \N__23227\
        );

    \I__3164\ : InMux
    port map (
            O => \N__23233\,
            I => \N__23224\
        );

    \I__3163\ : Span4Mux_v
    port map (
            O => \N__23230\,
            I => \N__23221\
        );

    \I__3162\ : Odrv12
    port map (
            O => \N__23227\,
            I => \nx.n3005\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__23224\,
            I => \nx.n3005\
        );

    \I__3160\ : Odrv4
    port map (
            O => \N__23221\,
            I => \nx.n3005\
        );

    \I__3159\ : InMux
    port map (
            O => \N__23214\,
            I => \N__23210\
        );

    \I__3158\ : InMux
    port map (
            O => \N__23213\,
            I => \N__23207\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__23210\,
            I => \N__23202\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__23207\,
            I => \N__23202\
        );

    \I__3155\ : Odrv4
    port map (
            O => \N__23202\,
            I => neo_pixel_transmitter_t0_7
        );

    \I__3154\ : InMux
    port map (
            O => \N__23199\,
            I => \N__23196\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__23196\,
            I => \nx.n26\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__23193\,
            I => \N__23189\
        );

    \I__3151\ : InMux
    port map (
            O => \N__23192\,
            I => \N__23186\
        );

    \I__3150\ : InMux
    port map (
            O => \N__23189\,
            I => \N__23183\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__23186\,
            I => \N__23179\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__23183\,
            I => \N__23176\
        );

    \I__3147\ : InMux
    port map (
            O => \N__23182\,
            I => \N__23173\
        );

    \I__3146\ : Span4Mux_s3_h
    port map (
            O => \N__23179\,
            I => \N__23168\
        );

    \I__3145\ : Span4Mux_v
    port map (
            O => \N__23176\,
            I => \N__23168\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__23173\,
            I => \nx.n3006\
        );

    \I__3143\ : Odrv4
    port map (
            O => \N__23168\,
            I => \nx.n3006\
        );

    \I__3142\ : CascadeMux
    port map (
            O => \N__23163\,
            I => \nx.n2899_cascade_\
        );

    \I__3141\ : CascadeMux
    port map (
            O => \N__23160\,
            I => \N__23156\
        );

    \I__3140\ : InMux
    port map (
            O => \N__23159\,
            I => \N__23153\
        );

    \I__3139\ : InMux
    port map (
            O => \N__23156\,
            I => \N__23150\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__23153\,
            I => \N__23147\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__23150\,
            I => \N__23144\
        );

    \I__3136\ : Span4Mux_s3_h
    port map (
            O => \N__23147\,
            I => \N__23138\
        );

    \I__3135\ : Span4Mux_v
    port map (
            O => \N__23144\,
            I => \N__23138\
        );

    \I__3134\ : InMux
    port map (
            O => \N__23143\,
            I => \N__23135\
        );

    \I__3133\ : Odrv4
    port map (
            O => \N__23138\,
            I => \nx.n2998\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__23135\,
            I => \nx.n2998\
        );

    \I__3131\ : CascadeMux
    port map (
            O => \N__23130\,
            I => \nx.n2894_cascade_\
        );

    \I__3130\ : CascadeMux
    port map (
            O => \N__23127\,
            I => \N__23123\
        );

    \I__3129\ : CascadeMux
    port map (
            O => \N__23126\,
            I => \N__23120\
        );

    \I__3128\ : InMux
    port map (
            O => \N__23123\,
            I => \N__23117\
        );

    \I__3127\ : InMux
    port map (
            O => \N__23120\,
            I => \N__23114\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__23117\,
            I => \N__23111\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__23114\,
            I => \N__23108\
        );

    \I__3124\ : Span12Mux_s3_h
    port map (
            O => \N__23111\,
            I => \N__23105\
        );

    \I__3123\ : Span4Mux_v
    port map (
            O => \N__23108\,
            I => \N__23102\
        );

    \I__3122\ : Odrv12
    port map (
            O => \N__23105\,
            I => \nx.n2985\
        );

    \I__3121\ : Odrv4
    port map (
            O => \N__23102\,
            I => \nx.n2985\
        );

    \I__3120\ : CascadeMux
    port map (
            O => \N__23097\,
            I => \N__23094\
        );

    \I__3119\ : InMux
    port map (
            O => \N__23094\,
            I => \N__23091\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__23091\,
            I => \N__23088\
        );

    \I__3117\ : Span4Mux_v
    port map (
            O => \N__23088\,
            I => \N__23085\
        );

    \I__3116\ : Span4Mux_h
    port map (
            O => \N__23085\,
            I => \N__23082\
        );

    \I__3115\ : Odrv4
    port map (
            O => \N__23082\,
            I => \nx.n5\
        );

    \I__3114\ : CascadeMux
    port map (
            O => \N__23079\,
            I => \N__23076\
        );

    \I__3113\ : InMux
    port map (
            O => \N__23076\,
            I => \N__23070\
        );

    \I__3112\ : InMux
    port map (
            O => \N__23075\,
            I => \N__23070\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__23070\,
            I => neo_pixel_transmitter_t0_25
        );

    \I__3110\ : InMux
    port map (
            O => \N__23067\,
            I => \N__23064\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__23064\,
            I => \N__23061\
        );

    \I__3108\ : Span4Mux_v
    port map (
            O => \N__23061\,
            I => \N__23058\
        );

    \I__3107\ : Odrv4
    port map (
            O => \N__23058\,
            I => \nx.n8\
        );

    \I__3106\ : InMux
    port map (
            O => \N__23055\,
            I => \N__23049\
        );

    \I__3105\ : InMux
    port map (
            O => \N__23054\,
            I => \N__23049\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__23049\,
            I => neo_pixel_transmitter_t0_18
        );

    \I__3103\ : InMux
    port map (
            O => \N__23046\,
            I => \N__23043\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__23043\,
            I => \N__23040\
        );

    \I__3101\ : Span4Mux_v
    port map (
            O => \N__23040\,
            I => \N__23037\
        );

    \I__3100\ : Odrv4
    port map (
            O => \N__23037\,
            I => \nx.n15\
        );

    \I__3099\ : InMux
    port map (
            O => \N__23034\,
            I => \N__23031\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__23031\,
            I => \N__23026\
        );

    \I__3097\ : InMux
    port map (
            O => \N__23030\,
            I => \N__23023\
        );

    \I__3096\ : InMux
    port map (
            O => \N__23029\,
            I => \N__23020\
        );

    \I__3095\ : Span12Mux_s8_v
    port map (
            O => \N__23026\,
            I => \N__23017\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__23023\,
            I => timer_28
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__23020\,
            I => timer_28
        );

    \I__3092\ : Odrv12
    port map (
            O => \N__23017\,
            I => timer_28
        );

    \I__3091\ : CascadeMux
    port map (
            O => \N__23010\,
            I => \N__23007\
        );

    \I__3090\ : InMux
    port map (
            O => \N__23007\,
            I => \N__23001\
        );

    \I__3089\ : InMux
    port map (
            O => \N__23006\,
            I => \N__23001\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__23001\,
            I => neo_pixel_transmitter_t0_28
        );

    \I__3087\ : CascadeMux
    port map (
            O => \N__22998\,
            I => \nx.n2995_cascade_\
        );

    \I__3086\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22992\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__22992\,
            I => \nx.n44_adj_681\
        );

    \I__3084\ : CascadeMux
    port map (
            O => \N__22989\,
            I => \nx.n33_adj_682_cascade_\
        );

    \I__3083\ : InMux
    port map (
            O => \N__22986\,
            I => \N__22983\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__22983\,
            I => \N__22980\
        );

    \I__3081\ : Span4Mux_s3_h
    port map (
            O => \N__22980\,
            I => \N__22977\
        );

    \I__3080\ : Odrv4
    port map (
            O => \N__22977\,
            I => \nx.n48\
        );

    \I__3079\ : CascadeMux
    port map (
            O => \N__22974\,
            I => \N__22971\
        );

    \I__3078\ : InMux
    port map (
            O => \N__22971\,
            I => \N__22966\
        );

    \I__3077\ : InMux
    port map (
            O => \N__22970\,
            I => \N__22963\
        );

    \I__3076\ : InMux
    port map (
            O => \N__22969\,
            I => \N__22960\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__22966\,
            I => \N__22957\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__22963\,
            I => timer_21
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__22960\,
            I => timer_21
        );

    \I__3072\ : Odrv12
    port map (
            O => \N__22957\,
            I => timer_21
        );

    \I__3071\ : CascadeMux
    port map (
            O => \N__22950\,
            I => \N__22947\
        );

    \I__3070\ : InMux
    port map (
            O => \N__22947\,
            I => \N__22944\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__22944\,
            I => \N__22939\
        );

    \I__3068\ : InMux
    port map (
            O => \N__22943\,
            I => \N__22936\
        );

    \I__3067\ : InMux
    port map (
            O => \N__22942\,
            I => \N__22933\
        );

    \I__3066\ : Span4Mux_v
    port map (
            O => \N__22939\,
            I => \N__22930\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__22936\,
            I => timer_13
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__22933\,
            I => timer_13
        );

    \I__3063\ : Odrv4
    port map (
            O => \N__22930\,
            I => timer_13
        );

    \I__3062\ : InMux
    port map (
            O => \N__22923\,
            I => \N__22919\
        );

    \I__3061\ : InMux
    port map (
            O => \N__22922\,
            I => \N__22916\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__22919\,
            I => neo_pixel_transmitter_t0_11
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__22916\,
            I => neo_pixel_transmitter_t0_11
        );

    \I__3058\ : InMux
    port map (
            O => \N__22911\,
            I => \N__22908\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__22908\,
            I => \N__22905\
        );

    \I__3056\ : Span4Mux_h
    port map (
            O => \N__22905\,
            I => \N__22902\
        );

    \I__3055\ : Odrv4
    port map (
            O => \N__22902\,
            I => \nx.n22_adj_618\
        );

    \I__3054\ : InMux
    port map (
            O => \N__22899\,
            I => \N__22893\
        );

    \I__3053\ : InMux
    port map (
            O => \N__22898\,
            I => \N__22893\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__22893\,
            I => neo_pixel_transmitter_t0_13
        );

    \I__3051\ : InMux
    port map (
            O => \N__22890\,
            I => \N__22887\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__22887\,
            I => \N__22884\
        );

    \I__3049\ : Odrv4
    port map (
            O => \N__22884\,
            I => \nx.n20\
        );

    \I__3048\ : CascadeMux
    port map (
            O => \N__22881\,
            I => \N__22878\
        );

    \I__3047\ : InMux
    port map (
            O => \N__22878\,
            I => \N__22874\
        );

    \I__3046\ : InMux
    port map (
            O => \N__22877\,
            I => \N__22871\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__22874\,
            I => \N__22867\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__22871\,
            I => \N__22864\
        );

    \I__3043\ : InMux
    port map (
            O => \N__22870\,
            I => \N__22861\
        );

    \I__3042\ : Span4Mux_v
    port map (
            O => \N__22867\,
            I => \N__22858\
        );

    \I__3041\ : Odrv4
    port map (
            O => \N__22864\,
            I => timer_7
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__22861\,
            I => timer_7
        );

    \I__3039\ : Odrv4
    port map (
            O => \N__22858\,
            I => timer_7
        );

    \I__3038\ : InMux
    port map (
            O => \N__22851\,
            I => \N__22848\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__22848\,
            I => \N__22845\
        );

    \I__3036\ : Span4Mux_s3_h
    port map (
            O => \N__22845\,
            I => \N__22842\
        );

    \I__3035\ : Odrv4
    port map (
            O => \N__22842\,
            I => \nx.n13159\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__22839\,
            I => \N__22836\
        );

    \I__3033\ : InMux
    port map (
            O => \N__22836\,
            I => \N__22830\
        );

    \I__3032\ : InMux
    port map (
            O => \N__22835\,
            I => \N__22830\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__22830\,
            I => neo_pixel_transmitter_t0_21
        );

    \I__3030\ : InMux
    port map (
            O => \N__22827\,
            I => \N__22824\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__22824\,
            I => \N__22821\
        );

    \I__3028\ : Span4Mux_v
    port map (
            O => \N__22821\,
            I => \N__22818\
        );

    \I__3027\ : Odrv4
    port map (
            O => \N__22818\,
            I => \nx.n12\
        );

    \I__3026\ : CascadeMux
    port map (
            O => \N__22815\,
            I => \N__22812\
        );

    \I__3025\ : InMux
    port map (
            O => \N__22812\,
            I => \N__22809\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__22809\,
            I => \N__22804\
        );

    \I__3023\ : InMux
    port map (
            O => \N__22808\,
            I => \N__22801\
        );

    \I__3022\ : InMux
    port map (
            O => \N__22807\,
            I => \N__22798\
        );

    \I__3021\ : Span4Mux_v
    port map (
            O => \N__22804\,
            I => \N__22795\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__22801\,
            I => timer_25
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__22798\,
            I => timer_25
        );

    \I__3018\ : Odrv4
    port map (
            O => \N__22795\,
            I => timer_25
        );

    \I__3017\ : CascadeMux
    port map (
            O => \N__22788\,
            I => \N__22785\
        );

    \I__3016\ : InMux
    port map (
            O => \N__22785\,
            I => \N__22780\
        );

    \I__3015\ : InMux
    port map (
            O => \N__22784\,
            I => \N__22777\
        );

    \I__3014\ : InMux
    port map (
            O => \N__22783\,
            I => \N__22774\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__22780\,
            I => \N__22771\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__22777\,
            I => timer_18
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__22774\,
            I => timer_18
        );

    \I__3010\ : Odrv12
    port map (
            O => \N__22771\,
            I => timer_18
        );

    \I__3009\ : InMux
    port map (
            O => \N__22764\,
            I => \N__22761\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__22761\,
            I => \N__22758\
        );

    \I__3007\ : Span4Mux_v
    port map (
            O => \N__22758\,
            I => \N__22755\
        );

    \I__3006\ : Odrv4
    port map (
            O => \N__22755\,
            I => \nx.n31_adj_650\
        );

    \I__3005\ : CascadeMux
    port map (
            O => \N__22752\,
            I => \N__22749\
        );

    \I__3004\ : InMux
    port map (
            O => \N__22749\,
            I => \N__22746\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__22746\,
            I => \N__22743\
        );

    \I__3002\ : Span4Mux_v
    port map (
            O => \N__22743\,
            I => \N__22740\
        );

    \I__3001\ : Odrv4
    port map (
            O => \N__22740\,
            I => \nx.n16_adj_661\
        );

    \I__3000\ : InMux
    port map (
            O => \N__22737\,
            I => \N__22733\
        );

    \I__2999\ : InMux
    port map (
            O => \N__22736\,
            I => \N__22730\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__22733\,
            I => \N__22726\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__22730\,
            I => \N__22723\
        );

    \I__2996\ : InMux
    port map (
            O => \N__22729\,
            I => \N__22720\
        );

    \I__2995\ : Span4Mux_v
    port map (
            O => \N__22726\,
            I => \N__22717\
        );

    \I__2994\ : Odrv4
    port map (
            O => \N__22723\,
            I => timer_17
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__22720\,
            I => timer_17
        );

    \I__2992\ : Odrv4
    port map (
            O => \N__22717\,
            I => timer_17
        );

    \I__2991\ : CascadeMux
    port map (
            O => \N__22710\,
            I => \N__22707\
        );

    \I__2990\ : InMux
    port map (
            O => \N__22707\,
            I => \N__22701\
        );

    \I__2989\ : InMux
    port map (
            O => \N__22706\,
            I => \N__22701\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__22701\,
            I => neo_pixel_transmitter_t0_17
        );

    \I__2987\ : CascadeMux
    port map (
            O => \N__22698\,
            I => \N__22695\
        );

    \I__2986\ : InMux
    port map (
            O => \N__22695\,
            I => \N__22690\
        );

    \I__2985\ : InMux
    port map (
            O => \N__22694\,
            I => \N__22687\
        );

    \I__2984\ : InMux
    port map (
            O => \N__22693\,
            I => \N__22684\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__22690\,
            I => \N__22681\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__22687\,
            I => timer_2
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__22684\,
            I => timer_2
        );

    \I__2980\ : Odrv12
    port map (
            O => \N__22681\,
            I => timer_2
        );

    \I__2979\ : InMux
    port map (
            O => \N__22674\,
            I => \N__22670\
        );

    \I__2978\ : InMux
    port map (
            O => \N__22673\,
            I => \N__22667\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__22670\,
            I => neo_pixel_transmitter_t0_2
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__22667\,
            I => neo_pixel_transmitter_t0_2
        );

    \I__2975\ : InMux
    port map (
            O => \N__22662\,
            I => \N__22658\
        );

    \I__2974\ : InMux
    port map (
            O => \N__22661\,
            I => \N__22655\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__22658\,
            I => \N__22651\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__22655\,
            I => \N__22648\
        );

    \I__2971\ : InMux
    port map (
            O => \N__22654\,
            I => \N__22645\
        );

    \I__2970\ : Span4Mux_v
    port map (
            O => \N__22651\,
            I => \N__22642\
        );

    \I__2969\ : Odrv4
    port map (
            O => \N__22648\,
            I => timer_29
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__22645\,
            I => timer_29
        );

    \I__2967\ : Odrv4
    port map (
            O => \N__22642\,
            I => timer_29
        );

    \I__2966\ : CascadeMux
    port map (
            O => \N__22635\,
            I => \N__22632\
        );

    \I__2965\ : InMux
    port map (
            O => \N__22632\,
            I => \N__22627\
        );

    \I__2964\ : InMux
    port map (
            O => \N__22631\,
            I => \N__22624\
        );

    \I__2963\ : InMux
    port map (
            O => \N__22630\,
            I => \N__22621\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__22627\,
            I => \N__22618\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__22624\,
            I => timer_9
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__22621\,
            I => timer_9
        );

    \I__2959\ : Odrv12
    port map (
            O => \N__22618\,
            I => timer_9
        );

    \I__2958\ : InMux
    port map (
            O => \N__22611\,
            I => \N__22607\
        );

    \I__2957\ : InMux
    port map (
            O => \N__22610\,
            I => \N__22604\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__22607\,
            I => \N__22601\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__22604\,
            I => neo_pixel_transmitter_t0_10
        );

    \I__2954\ : Odrv4
    port map (
            O => \N__22601\,
            I => neo_pixel_transmitter_t0_10
        );

    \I__2953\ : InMux
    port map (
            O => \N__22596\,
            I => \N__22593\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__22593\,
            I => \N__22590\
        );

    \I__2951\ : Span4Mux_v
    port map (
            O => \N__22590\,
            I => \N__22587\
        );

    \I__2950\ : Odrv4
    port map (
            O => \N__22587\,
            I => \nx.n23_adj_617\
        );

    \I__2949\ : InMux
    port map (
            O => \N__22584\,
            I => \N__22578\
        );

    \I__2948\ : InMux
    port map (
            O => \N__22583\,
            I => \N__22578\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__22578\,
            I => neo_pixel_transmitter_t0_29
        );

    \I__2946\ : CascadeMux
    port map (
            O => \N__22575\,
            I => \N__22572\
        );

    \I__2945\ : InMux
    port map (
            O => \N__22572\,
            I => \N__22569\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__22569\,
            I => \N__22566\
        );

    \I__2943\ : Span4Mux_s3_h
    port map (
            O => \N__22566\,
            I => \N__22563\
        );

    \I__2942\ : Span4Mux_v
    port map (
            O => \N__22563\,
            I => \N__22560\
        );

    \I__2941\ : Odrv4
    port map (
            O => \N__22560\,
            I => \nx.n4\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__22557\,
            I => \N__22554\
        );

    \I__2939\ : InMux
    port map (
            O => \N__22554\,
            I => \N__22549\
        );

    \I__2938\ : InMux
    port map (
            O => \N__22553\,
            I => \N__22546\
        );

    \I__2937\ : InMux
    port map (
            O => \N__22552\,
            I => \N__22543\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__22549\,
            I => \N__22540\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__22546\,
            I => timer_11
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__22543\,
            I => timer_11
        );

    \I__2933\ : Odrv12
    port map (
            O => \N__22540\,
            I => timer_11
        );

    \I__2932\ : InMux
    port map (
            O => \N__22533\,
            I => \nx.n10588\
        );

    \I__2931\ : InMux
    port map (
            O => \N__22530\,
            I => \bfn_3_32_0_\
        );

    \I__2930\ : InMux
    port map (
            O => \N__22527\,
            I => \nx.n10590\
        );

    \I__2929\ : InMux
    port map (
            O => \N__22524\,
            I => \nx.n10591\
        );

    \I__2928\ : InMux
    port map (
            O => \N__22521\,
            I => \N__22518\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__22518\,
            I => \N__22513\
        );

    \I__2926\ : CascadeMux
    port map (
            O => \N__22517\,
            I => \N__22510\
        );

    \I__2925\ : CascadeMux
    port map (
            O => \N__22516\,
            I => \N__22507\
        );

    \I__2924\ : Span4Mux_s2_v
    port map (
            O => \N__22513\,
            I => \N__22504\
        );

    \I__2923\ : InMux
    port map (
            O => \N__22510\,
            I => \N__22501\
        );

    \I__2922\ : InMux
    port map (
            O => \N__22507\,
            I => \N__22498\
        );

    \I__2921\ : Odrv4
    port map (
            O => \N__22504\,
            I => \nx.n1303\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__22501\,
            I => \nx.n1303\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__22498\,
            I => \nx.n1303\
        );

    \I__2918\ : CascadeMux
    port map (
            O => \N__22491\,
            I => \N__22488\
        );

    \I__2917\ : InMux
    port map (
            O => \N__22488\,
            I => \N__22485\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__22485\,
            I => \nx.n1370\
        );

    \I__2915\ : InMux
    port map (
            O => \N__22482\,
            I => \N__22476\
        );

    \I__2914\ : InMux
    port map (
            O => \N__22481\,
            I => \N__22476\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__22476\,
            I => \nx.n1400\
        );

    \I__2912\ : CascadeMux
    port map (
            O => \N__22473\,
            I => \N__22470\
        );

    \I__2911\ : InMux
    port map (
            O => \N__22470\,
            I => \N__22467\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__22467\,
            I => \N__22464\
        );

    \I__2909\ : Span4Mux_v
    port map (
            O => \N__22464\,
            I => \N__22461\
        );

    \I__2908\ : Span4Mux_v
    port map (
            O => \N__22461\,
            I => \N__22458\
        );

    \I__2907\ : Odrv4
    port map (
            O => \N__22458\,
            I => \nx.n3\
        );

    \I__2906\ : InMux
    port map (
            O => \N__22455\,
            I => \N__22451\
        );

    \I__2905\ : InMux
    port map (
            O => \N__22454\,
            I => \N__22448\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__22451\,
            I => \N__22445\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__22448\,
            I => \N__22441\
        );

    \I__2902\ : Span4Mux_v
    port map (
            O => \N__22445\,
            I => \N__22438\
        );

    \I__2901\ : InMux
    port map (
            O => \N__22444\,
            I => \N__22435\
        );

    \I__2900\ : Span4Mux_v
    port map (
            O => \N__22441\,
            I => \N__22432\
        );

    \I__2899\ : Odrv4
    port map (
            O => \N__22438\,
            I => timer_30
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__22435\,
            I => timer_30
        );

    \I__2897\ : Odrv4
    port map (
            O => \N__22432\,
            I => timer_30
        );

    \I__2896\ : InMux
    port map (
            O => \N__22425\,
            I => \N__22419\
        );

    \I__2895\ : InMux
    port map (
            O => \N__22424\,
            I => \N__22419\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__22419\,
            I => neo_pixel_transmitter_t0_30
        );

    \I__2893\ : InMux
    port map (
            O => \N__22416\,
            I => \N__22413\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__22413\,
            I => \N__22410\
        );

    \I__2891\ : Span4Mux_h
    port map (
            O => \N__22410\,
            I => \N__22407\
        );

    \I__2890\ : Odrv4
    port map (
            O => \N__22407\,
            I => \nx.n1272\
        );

    \I__2889\ : CascadeMux
    port map (
            O => \N__22404\,
            I => \N__22400\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__22403\,
            I => \N__22397\
        );

    \I__2887\ : InMux
    port map (
            O => \N__22400\,
            I => \N__22393\
        );

    \I__2886\ : InMux
    port map (
            O => \N__22397\,
            I => \N__22390\
        );

    \I__2885\ : InMux
    port map (
            O => \N__22396\,
            I => \N__22387\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__22393\,
            I => \nx.n1205\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__22390\,
            I => \nx.n1205\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__22387\,
            I => \nx.n1205\
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__22380\,
            I => \N__22374\
        );

    \I__2880\ : CascadeMux
    port map (
            O => \N__22379\,
            I => \N__22371\
        );

    \I__2879\ : CascadeMux
    port map (
            O => \N__22378\,
            I => \N__22368\
        );

    \I__2878\ : InMux
    port map (
            O => \N__22377\,
            I => \N__22355\
        );

    \I__2877\ : InMux
    port map (
            O => \N__22374\,
            I => \N__22355\
        );

    \I__2876\ : InMux
    port map (
            O => \N__22371\,
            I => \N__22355\
        );

    \I__2875\ : InMux
    port map (
            O => \N__22368\,
            I => \N__22355\
        );

    \I__2874\ : InMux
    port map (
            O => \N__22367\,
            I => \N__22350\
        );

    \I__2873\ : InMux
    port map (
            O => \N__22366\,
            I => \N__22350\
        );

    \I__2872\ : InMux
    port map (
            O => \N__22365\,
            I => \N__22345\
        );

    \I__2871\ : InMux
    port map (
            O => \N__22364\,
            I => \N__22345\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__22355\,
            I => \N__22342\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__22350\,
            I => \nx.n1235\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__22345\,
            I => \nx.n1235\
        );

    \I__2867\ : Odrv4
    port map (
            O => \N__22342\,
            I => \nx.n1235\
        );

    \I__2866\ : InMux
    port map (
            O => \N__22335\,
            I => \N__22332\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__22332\,
            I => \nx.n1377\
        );

    \I__2864\ : InMux
    port map (
            O => \N__22329\,
            I => \bfn_3_31_0_\
        );

    \I__2863\ : InMux
    port map (
            O => \N__22326\,
            I => \nx.n10582\
        );

    \I__2862\ : InMux
    port map (
            O => \N__22323\,
            I => \nx.n10583\
        );

    \I__2861\ : InMux
    port map (
            O => \N__22320\,
            I => \nx.n10584\
        );

    \I__2860\ : InMux
    port map (
            O => \N__22317\,
            I => \nx.n10585\
        );

    \I__2859\ : InMux
    port map (
            O => \N__22314\,
            I => \nx.n10586\
        );

    \I__2858\ : InMux
    port map (
            O => \N__22311\,
            I => \nx.n10587\
        );

    \I__2857\ : InMux
    port map (
            O => \N__22308\,
            I => \N__22305\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__22305\,
            I => \N__22302\
        );

    \I__2855\ : Span4Mux_v
    port map (
            O => \N__22302\,
            I => \N__22299\
        );

    \I__2854\ : Odrv4
    port map (
            O => \N__22299\,
            I => \nx.n3053\
        );

    \I__2853\ : InMux
    port map (
            O => \N__22296\,
            I => \bfn_3_29_0_\
        );

    \I__2852\ : InMux
    port map (
            O => \N__22293\,
            I => \N__22290\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__22290\,
            I => \nx.n3052\
        );

    \I__2850\ : InMux
    port map (
            O => \N__22287\,
            I => \nx.n10886\
        );

    \I__2849\ : InMux
    port map (
            O => \N__22284\,
            I => \nx.n10887\
        );

    \I__2848\ : CascadeMux
    port map (
            O => \N__22281\,
            I => \N__22278\
        );

    \I__2847\ : InMux
    port map (
            O => \N__22278\,
            I => \N__22274\
        );

    \I__2846\ : InMux
    port map (
            O => \N__22277\,
            I => \N__22271\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__22274\,
            I => \N__22268\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__22271\,
            I => \N__22265\
        );

    \I__2843\ : Span4Mux_s2_h
    port map (
            O => \N__22268\,
            I => \N__22262\
        );

    \I__2842\ : Odrv4
    port map (
            O => \N__22265\,
            I => \nx.n3083\
        );

    \I__2841\ : Odrv4
    port map (
            O => \N__22262\,
            I => \nx.n3083\
        );

    \I__2840\ : InMux
    port map (
            O => \N__22257\,
            I => \N__22254\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__22254\,
            I => \nx.n45_adj_707\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__22251\,
            I => \nx.n11_adj_628_cascade_\
        );

    \I__2837\ : InMux
    port map (
            O => \N__22248\,
            I => \N__22245\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__22245\,
            I => \nx.n16_adj_627\
        );

    \I__2835\ : InMux
    port map (
            O => \N__22242\,
            I => \N__22237\
        );

    \I__2834\ : InMux
    port map (
            O => \N__22241\,
            I => \N__22234\
        );

    \I__2833\ : InMux
    port map (
            O => \N__22240\,
            I => \N__22231\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__22237\,
            I => \nx.n1307\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__22234\,
            I => \nx.n1307\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__22231\,
            I => \nx.n1307\
        );

    \I__2829\ : CascadeMux
    port map (
            O => \N__22224\,
            I => \nx.n1334_cascade_\
        );

    \I__2828\ : InMux
    port map (
            O => \N__22221\,
            I => \N__22218\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__22218\,
            I => \nx.n1374\
        );

    \I__2826\ : InMux
    port map (
            O => \N__22215\,
            I => \N__22212\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__22212\,
            I => \N__22209\
        );

    \I__2824\ : Span4Mux_v
    port map (
            O => \N__22209\,
            I => \N__22206\
        );

    \I__2823\ : Odrv4
    port map (
            O => \N__22206\,
            I => \nx.n1277\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__22203\,
            I => \N__22199\
        );

    \I__2821\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22196\
        );

    \I__2820\ : InMux
    port map (
            O => \N__22199\,
            I => \N__22193\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__22196\,
            I => \nx.n1309\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__22193\,
            I => \nx.n1309\
        );

    \I__2817\ : InMux
    port map (
            O => \N__22188\,
            I => \N__22185\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__22185\,
            I => \nx.n1376\
        );

    \I__2815\ : CascadeMux
    port map (
            O => \N__22182\,
            I => \nx.n1309_cascade_\
        );

    \I__2814\ : InMux
    port map (
            O => \N__22179\,
            I => \bfn_3_28_0_\
        );

    \I__2813\ : InMux
    port map (
            O => \N__22176\,
            I => \nx.n10878\
        );

    \I__2812\ : InMux
    port map (
            O => \N__22173\,
            I => \N__22170\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__22170\,
            I => \nx.n3059\
        );

    \I__2810\ : InMux
    port map (
            O => \N__22167\,
            I => \nx.n10879\
        );

    \I__2809\ : InMux
    port map (
            O => \N__22164\,
            I => \nx.n10880\
        );

    \I__2808\ : InMux
    port map (
            O => \N__22161\,
            I => \nx.n10881\
        );

    \I__2807\ : InMux
    port map (
            O => \N__22158\,
            I => \nx.n10882\
        );

    \I__2806\ : InMux
    port map (
            O => \N__22155\,
            I => \N__22152\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__22152\,
            I => \N__22149\
        );

    \I__2804\ : Span4Mux_v
    port map (
            O => \N__22149\,
            I => \N__22146\
        );

    \I__2803\ : Odrv4
    port map (
            O => \N__22146\,
            I => \nx.n3055\
        );

    \I__2802\ : InMux
    port map (
            O => \N__22143\,
            I => \nx.n10883\
        );

    \I__2801\ : InMux
    port map (
            O => \N__22140\,
            I => \N__22137\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__22137\,
            I => \N__22134\
        );

    \I__2799\ : Span4Mux_v
    port map (
            O => \N__22134\,
            I => \N__22131\
        );

    \I__2798\ : Odrv4
    port map (
            O => \N__22131\,
            I => \nx.n3054\
        );

    \I__2797\ : InMux
    port map (
            O => \N__22128\,
            I => \nx.n10884\
        );

    \I__2796\ : CascadeMux
    port map (
            O => \N__22125\,
            I => \N__22122\
        );

    \I__2795\ : InMux
    port map (
            O => \N__22122\,
            I => \N__22119\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__22119\,
            I => \N__22116\
        );

    \I__2793\ : Span4Mux_v
    port map (
            O => \N__22116\,
            I => \N__22113\
        );

    \I__2792\ : Odrv4
    port map (
            O => \N__22113\,
            I => \nx.n3070\
        );

    \I__2791\ : InMux
    port map (
            O => \N__22110\,
            I => \nx.n10868\
        );

    \I__2790\ : InMux
    port map (
            O => \N__22107\,
            I => \N__22104\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__22104\,
            I => \N__22101\
        );

    \I__2788\ : Span4Mux_s2_h
    port map (
            O => \N__22101\,
            I => \N__22098\
        );

    \I__2787\ : Odrv4
    port map (
            O => \N__22098\,
            I => \nx.n3069\
        );

    \I__2786\ : InMux
    port map (
            O => \N__22095\,
            I => \bfn_3_27_0_\
        );

    \I__2785\ : CascadeMux
    port map (
            O => \N__22092\,
            I => \N__22089\
        );

    \I__2784\ : InMux
    port map (
            O => \N__22089\,
            I => \N__22086\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__22086\,
            I => \N__22081\
        );

    \I__2782\ : InMux
    port map (
            O => \N__22085\,
            I => \N__22078\
        );

    \I__2781\ : InMux
    port map (
            O => \N__22084\,
            I => \N__22075\
        );

    \I__2780\ : Span4Mux_v
    port map (
            O => \N__22081\,
            I => \N__22072\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__22078\,
            I => \nx.n3001\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__22075\,
            I => \nx.n3001\
        );

    \I__2777\ : Odrv4
    port map (
            O => \N__22072\,
            I => \nx.n3001\
        );

    \I__2776\ : InMux
    port map (
            O => \N__22065\,
            I => \N__22062\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__22062\,
            I => \N__22059\
        );

    \I__2774\ : Span4Mux_s2_h
    port map (
            O => \N__22059\,
            I => \N__22056\
        );

    \I__2773\ : Odrv4
    port map (
            O => \N__22056\,
            I => \nx.n3068\
        );

    \I__2772\ : InMux
    port map (
            O => \N__22053\,
            I => \nx.n10870\
        );

    \I__2771\ : CascadeMux
    port map (
            O => \N__22050\,
            I => \N__22047\
        );

    \I__2770\ : InMux
    port map (
            O => \N__22047\,
            I => \N__22044\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__22044\,
            I => \nx.n3067\
        );

    \I__2768\ : InMux
    port map (
            O => \N__22041\,
            I => \nx.n10871\
        );

    \I__2767\ : CascadeMux
    port map (
            O => \N__22038\,
            I => \N__22035\
        );

    \I__2766\ : InMux
    port map (
            O => \N__22035\,
            I => \N__22032\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__22032\,
            I => \N__22027\
        );

    \I__2764\ : InMux
    port map (
            O => \N__22031\,
            I => \N__22024\
        );

    \I__2763\ : InMux
    port map (
            O => \N__22030\,
            I => \N__22021\
        );

    \I__2762\ : Span4Mux_v
    port map (
            O => \N__22027\,
            I => \N__22018\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__22024\,
            I => \nx.n2999\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__22021\,
            I => \nx.n2999\
        );

    \I__2759\ : Odrv4
    port map (
            O => \N__22018\,
            I => \nx.n2999\
        );

    \I__2758\ : CascadeMux
    port map (
            O => \N__22011\,
            I => \N__22008\
        );

    \I__2757\ : InMux
    port map (
            O => \N__22008\,
            I => \N__22005\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__22005\,
            I => \N__22002\
        );

    \I__2755\ : Odrv4
    port map (
            O => \N__22002\,
            I => \nx.n3066\
        );

    \I__2754\ : InMux
    port map (
            O => \N__21999\,
            I => \nx.n10872\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__21996\,
            I => \N__21993\
        );

    \I__2752\ : InMux
    port map (
            O => \N__21993\,
            I => \N__21990\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__21990\,
            I => \N__21987\
        );

    \I__2750\ : Odrv4
    port map (
            O => \N__21987\,
            I => \nx.n3065\
        );

    \I__2749\ : InMux
    port map (
            O => \N__21984\,
            I => \nx.n10873\
        );

    \I__2748\ : CascadeMux
    port map (
            O => \N__21981\,
            I => \N__21978\
        );

    \I__2747\ : InMux
    port map (
            O => \N__21978\,
            I => \N__21975\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__21975\,
            I => \N__21972\
        );

    \I__2745\ : Span4Mux_s3_h
    port map (
            O => \N__21972\,
            I => \N__21969\
        );

    \I__2744\ : Odrv4
    port map (
            O => \N__21969\,
            I => \nx.n3064\
        );

    \I__2743\ : InMux
    port map (
            O => \N__21966\,
            I => \nx.n10874\
        );

    \I__2742\ : InMux
    port map (
            O => \N__21963\,
            I => \N__21960\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__21960\,
            I => \N__21957\
        );

    \I__2740\ : Span4Mux_s1_h
    port map (
            O => \N__21957\,
            I => \N__21954\
        );

    \I__2739\ : Span4Mux_v
    port map (
            O => \N__21954\,
            I => \N__21951\
        );

    \I__2738\ : Odrv4
    port map (
            O => \N__21951\,
            I => \nx.n3063\
        );

    \I__2737\ : InMux
    port map (
            O => \N__21948\,
            I => \nx.n10875\
        );

    \I__2736\ : InMux
    port map (
            O => \N__21945\,
            I => \nx.n10876\
        );

    \I__2735\ : InMux
    port map (
            O => \N__21942\,
            I => \N__21936\
        );

    \I__2734\ : InMux
    port map (
            O => \N__21941\,
            I => \N__21936\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__21936\,
            I => neo_pixel_transmitter_t0_27
        );

    \I__2732\ : InMux
    port map (
            O => \N__21933\,
            I => \N__21930\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__21930\,
            I => \nx.n6\
        );

    \I__2730\ : InMux
    port map (
            O => \N__21927\,
            I => \N__21924\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__21924\,
            I => \N__21921\
        );

    \I__2728\ : Odrv4
    port map (
            O => \N__21921\,
            I => \nx.n3077\
        );

    \I__2727\ : InMux
    port map (
            O => \N__21918\,
            I => \bfn_3_26_0_\
        );

    \I__2726\ : InMux
    port map (
            O => \N__21915\,
            I => \N__21912\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__21912\,
            I => \nx.n3076\
        );

    \I__2724\ : InMux
    port map (
            O => \N__21909\,
            I => \nx.n10862\
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__21906\,
            I => \N__21902\
        );

    \I__2722\ : InMux
    port map (
            O => \N__21905\,
            I => \N__21899\
        );

    \I__2721\ : InMux
    port map (
            O => \N__21902\,
            I => \N__21896\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__21899\,
            I => \N__21891\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__21896\,
            I => \N__21891\
        );

    \I__2718\ : Odrv4
    port map (
            O => \N__21891\,
            I => \nx.n3008\
        );

    \I__2717\ : CascadeMux
    port map (
            O => \N__21888\,
            I => \N__21885\
        );

    \I__2716\ : InMux
    port map (
            O => \N__21885\,
            I => \N__21882\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__21882\,
            I => \nx.n3075\
        );

    \I__2714\ : InMux
    port map (
            O => \N__21879\,
            I => \nx.n10863\
        );

    \I__2713\ : CascadeMux
    port map (
            O => \N__21876\,
            I => \N__21873\
        );

    \I__2712\ : InMux
    port map (
            O => \N__21873\,
            I => \N__21870\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__21870\,
            I => \N__21866\
        );

    \I__2710\ : InMux
    port map (
            O => \N__21869\,
            I => \N__21863\
        );

    \I__2709\ : Span4Mux_h
    port map (
            O => \N__21866\,
            I => \N__21860\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__21863\,
            I => \nx.n3007\
        );

    \I__2707\ : Odrv4
    port map (
            O => \N__21860\,
            I => \nx.n3007\
        );

    \I__2706\ : InMux
    port map (
            O => \N__21855\,
            I => \N__21852\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__21852\,
            I => \N__21849\
        );

    \I__2704\ : Span4Mux_s2_h
    port map (
            O => \N__21849\,
            I => \N__21846\
        );

    \I__2703\ : Odrv4
    port map (
            O => \N__21846\,
            I => \nx.n3074\
        );

    \I__2702\ : InMux
    port map (
            O => \N__21843\,
            I => \nx.n10864\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__21840\,
            I => \N__21837\
        );

    \I__2700\ : InMux
    port map (
            O => \N__21837\,
            I => \N__21834\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__21834\,
            I => \N__21831\
        );

    \I__2698\ : Span4Mux_s2_h
    port map (
            O => \N__21831\,
            I => \N__21828\
        );

    \I__2697\ : Odrv4
    port map (
            O => \N__21828\,
            I => \nx.n3073\
        );

    \I__2696\ : InMux
    port map (
            O => \N__21825\,
            I => \nx.n10865\
        );

    \I__2695\ : InMux
    port map (
            O => \N__21822\,
            I => \N__21819\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__21819\,
            I => \nx.n3072\
        );

    \I__2693\ : InMux
    port map (
            O => \N__21816\,
            I => \nx.n10866\
        );

    \I__2692\ : InMux
    port map (
            O => \N__21813\,
            I => \N__21810\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__21810\,
            I => \N__21807\
        );

    \I__2690\ : Odrv4
    port map (
            O => \N__21807\,
            I => \nx.n3071\
        );

    \I__2689\ : InMux
    port map (
            O => \N__21804\,
            I => \nx.n10867\
        );

    \I__2688\ : InMux
    port map (
            O => \N__21801\,
            I => \N__21798\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__21798\,
            I => \nx.n12973\
        );

    \I__2686\ : InMux
    port map (
            O => \N__21795\,
            I => \bfn_3_25_0_\
        );

    \I__2685\ : InMux
    port map (
            O => \N__21792\,
            I => \N__21789\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__21789\,
            I => \nx.n12975\
        );

    \I__2683\ : InMux
    port map (
            O => \N__21786\,
            I => \nx.n10449\
        );

    \I__2682\ : InMux
    port map (
            O => \N__21783\,
            I => \N__21780\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__21780\,
            I => \nx.n12977\
        );

    \I__2680\ : InMux
    port map (
            O => \N__21777\,
            I => \nx.n10450\
        );

    \I__2679\ : InMux
    port map (
            O => \N__21774\,
            I => \N__21771\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__21771\,
            I => \nx.n12979\
        );

    \I__2677\ : InMux
    port map (
            O => \N__21768\,
            I => \nx.n10451\
        );

    \I__2676\ : InMux
    port map (
            O => \N__21765\,
            I => \N__21761\
        );

    \I__2675\ : InMux
    port map (
            O => \N__21764\,
            I => \N__21758\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__21761\,
            I => \N__21754\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__21758\,
            I => \N__21751\
        );

    \I__2672\ : InMux
    port map (
            O => \N__21757\,
            I => \N__21748\
        );

    \I__2671\ : Span4Mux_v
    port map (
            O => \N__21754\,
            I => \N__21743\
        );

    \I__2670\ : Span4Mux_v
    port map (
            O => \N__21751\,
            I => \N__21743\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__21748\,
            I => timer_31
        );

    \I__2668\ : Odrv4
    port map (
            O => \N__21743\,
            I => timer_31
        );

    \I__2667\ : InMux
    port map (
            O => \N__21738\,
            I => \N__21735\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__21735\,
            I => \N__21732\
        );

    \I__2665\ : Span4Mux_v
    port map (
            O => \N__21732\,
            I => \N__21729\
        );

    \I__2664\ : Span4Mux_v
    port map (
            O => \N__21729\,
            I => \N__21726\
        );

    \I__2663\ : Odrv4
    port map (
            O => \N__21726\,
            I => \nx.n2\
        );

    \I__2662\ : CascadeMux
    port map (
            O => \N__21723\,
            I => \N__21720\
        );

    \I__2661\ : InMux
    port map (
            O => \N__21720\,
            I => \N__21717\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__21717\,
            I => \nx.n12981\
        );

    \I__2659\ : InMux
    port map (
            O => \N__21714\,
            I => \nx.n10452\
        );

    \I__2658\ : InMux
    port map (
            O => \N__21711\,
            I => \N__21706\
        );

    \I__2657\ : InMux
    port map (
            O => \N__21710\,
            I => \N__21703\
        );

    \I__2656\ : InMux
    port map (
            O => \N__21709\,
            I => \N__21700\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__21706\,
            I => \N__21697\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__21703\,
            I => \N__21692\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__21700\,
            I => \N__21692\
        );

    \I__2652\ : Span4Mux_s3_h
    port map (
            O => \N__21697\,
            I => \N__21689\
        );

    \I__2651\ : Span4Mux_s3_h
    port map (
            O => \N__21692\,
            I => \N__21686\
        );

    \I__2650\ : Span4Mux_v
    port map (
            O => \N__21689\,
            I => \N__21683\
        );

    \I__2649\ : Span4Mux_v
    port map (
            O => \N__21686\,
            I => \N__21680\
        );

    \I__2648\ : Odrv4
    port map (
            O => \N__21683\,
            I => \nx.n7181\
        );

    \I__2647\ : Odrv4
    port map (
            O => \N__21680\,
            I => \nx.n7181\
        );

    \I__2646\ : CascadeMux
    port map (
            O => \N__21675\,
            I => \N__21671\
        );

    \I__2645\ : InMux
    port map (
            O => \N__21674\,
            I => \N__21667\
        );

    \I__2644\ : InMux
    port map (
            O => \N__21671\,
            I => \N__21664\
        );

    \I__2643\ : InMux
    port map (
            O => \N__21670\,
            I => \N__21661\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__21667\,
            I => \N__21656\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__21664\,
            I => \N__21656\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__21661\,
            I => timer_27
        );

    \I__2639\ : Odrv12
    port map (
            O => \N__21656\,
            I => timer_27
        );

    \I__2638\ : InMux
    port map (
            O => \N__21651\,
            I => \N__21648\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__21648\,
            I => \nx.n12961\
        );

    \I__2636\ : InMux
    port map (
            O => \N__21645\,
            I => \bfn_3_24_0_\
        );

    \I__2635\ : InMux
    port map (
            O => \N__21642\,
            I => \N__21639\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__21639\,
            I => \nx.n12963\
        );

    \I__2633\ : InMux
    port map (
            O => \N__21636\,
            I => \nx.n10443\
        );

    \I__2632\ : InMux
    port map (
            O => \N__21633\,
            I => \N__21630\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__21630\,
            I => \nx.n12965\
        );

    \I__2630\ : InMux
    port map (
            O => \N__21627\,
            I => \N__21624\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__21624\,
            I => \N__21621\
        );

    \I__2628\ : Span4Mux_v
    port map (
            O => \N__21621\,
            I => \N__21618\
        );

    \I__2627\ : Span4Mux_v
    port map (
            O => \N__21618\,
            I => \N__21615\
        );

    \I__2626\ : Odrv4
    port map (
            O => \N__21615\,
            I => \nx.n10\
        );

    \I__2625\ : CascadeMux
    port map (
            O => \N__21612\,
            I => \N__21608\
        );

    \I__2624\ : InMux
    port map (
            O => \N__21611\,
            I => \N__21605\
        );

    \I__2623\ : InMux
    port map (
            O => \N__21608\,
            I => \N__21602\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__21605\,
            I => \N__21599\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__21602\,
            I => \N__21595\
        );

    \I__2620\ : Span4Mux_s2_h
    port map (
            O => \N__21599\,
            I => \N__21592\
        );

    \I__2619\ : InMux
    port map (
            O => \N__21598\,
            I => \N__21589\
        );

    \I__2618\ : Span4Mux_v
    port map (
            O => \N__21595\,
            I => \N__21586\
        );

    \I__2617\ : Odrv4
    port map (
            O => \N__21592\,
            I => timer_23
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__21589\,
            I => timer_23
        );

    \I__2615\ : Odrv4
    port map (
            O => \N__21586\,
            I => timer_23
        );

    \I__2614\ : InMux
    port map (
            O => \N__21579\,
            I => \nx.n10444\
        );

    \I__2613\ : InMux
    port map (
            O => \N__21576\,
            I => \N__21573\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__21573\,
            I => \N__21570\
        );

    \I__2611\ : Odrv4
    port map (
            O => \N__21570\,
            I => \nx.n12967\
        );

    \I__2610\ : InMux
    port map (
            O => \N__21567\,
            I => \N__21564\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__21564\,
            I => \N__21561\
        );

    \I__2608\ : Span4Mux_v
    port map (
            O => \N__21561\,
            I => \N__21558\
        );

    \I__2607\ : Odrv4
    port map (
            O => \N__21558\,
            I => \nx.n9\
        );

    \I__2606\ : InMux
    port map (
            O => \N__21555\,
            I => \N__21551\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__21554\,
            I => \N__21548\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__21551\,
            I => \N__21544\
        );

    \I__2603\ : InMux
    port map (
            O => \N__21548\,
            I => \N__21541\
        );

    \I__2602\ : InMux
    port map (
            O => \N__21547\,
            I => \N__21538\
        );

    \I__2601\ : Sp12to4
    port map (
            O => \N__21544\,
            I => \N__21533\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__21541\,
            I => \N__21533\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__21538\,
            I => timer_24
        );

    \I__2598\ : Odrv12
    port map (
            O => \N__21533\,
            I => timer_24
        );

    \I__2597\ : InMux
    port map (
            O => \N__21528\,
            I => \nx.n10445\
        );

    \I__2596\ : InMux
    port map (
            O => \N__21525\,
            I => \N__21522\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__21522\,
            I => \N__21519\
        );

    \I__2594\ : Odrv4
    port map (
            O => \N__21519\,
            I => \nx.n12969\
        );

    \I__2593\ : InMux
    port map (
            O => \N__21516\,
            I => \nx.n10446\
        );

    \I__2592\ : InMux
    port map (
            O => \N__21513\,
            I => \N__21510\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__21510\,
            I => \nx.n12971\
        );

    \I__2590\ : InMux
    port map (
            O => \N__21507\,
            I => \N__21504\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__21504\,
            I => \N__21501\
        );

    \I__2588\ : Span4Mux_v
    port map (
            O => \N__21501\,
            I => \N__21498\
        );

    \I__2587\ : Span4Mux_h
    port map (
            O => \N__21498\,
            I => \N__21495\
        );

    \I__2586\ : Odrv4
    port map (
            O => \N__21495\,
            I => \nx.n7_adj_597\
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__21492\,
            I => \N__21488\
        );

    \I__2584\ : InMux
    port map (
            O => \N__21491\,
            I => \N__21485\
        );

    \I__2583\ : InMux
    port map (
            O => \N__21488\,
            I => \N__21482\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__21485\,
            I => \N__21476\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__21482\,
            I => \N__21476\
        );

    \I__2580\ : InMux
    port map (
            O => \N__21481\,
            I => \N__21473\
        );

    \I__2579\ : Span4Mux_v
    port map (
            O => \N__21476\,
            I => \N__21470\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__21473\,
            I => timer_26
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__21470\,
            I => timer_26
        );

    \I__2576\ : InMux
    port map (
            O => \N__21465\,
            I => \nx.n10447\
        );

    \I__2575\ : InMux
    port map (
            O => \N__21462\,
            I => \N__21459\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__21459\,
            I => \nx.n12947\
        );

    \I__2573\ : InMux
    port map (
            O => \N__21456\,
            I => \N__21453\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__21453\,
            I => \N__21450\
        );

    \I__2571\ : Odrv4
    port map (
            O => \N__21450\,
            I => \nx.n19_adj_622\
        );

    \I__2570\ : CascadeMux
    port map (
            O => \N__21447\,
            I => \N__21444\
        );

    \I__2569\ : InMux
    port map (
            O => \N__21444\,
            I => \N__21441\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__21441\,
            I => \N__21436\
        );

    \I__2567\ : InMux
    port map (
            O => \N__21440\,
            I => \N__21433\
        );

    \I__2566\ : InMux
    port map (
            O => \N__21439\,
            I => \N__21430\
        );

    \I__2565\ : Span4Mux_v
    port map (
            O => \N__21436\,
            I => \N__21427\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__21433\,
            I => timer_14
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__21430\,
            I => timer_14
        );

    \I__2562\ : Odrv4
    port map (
            O => \N__21427\,
            I => timer_14
        );

    \I__2561\ : InMux
    port map (
            O => \N__21420\,
            I => \nx.n10435\
        );

    \I__2560\ : InMux
    port map (
            O => \N__21417\,
            I => \N__21414\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__21414\,
            I => \nx.n12949\
        );

    \I__2558\ : InMux
    port map (
            O => \N__21411\,
            I => \N__21408\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__21408\,
            I => \N__21405\
        );

    \I__2556\ : Span4Mux_v
    port map (
            O => \N__21405\,
            I => \N__21402\
        );

    \I__2555\ : Odrv4
    port map (
            O => \N__21402\,
            I => \nx.n18_adj_623\
        );

    \I__2554\ : InMux
    port map (
            O => \N__21399\,
            I => \N__21395\
        );

    \I__2553\ : CascadeMux
    port map (
            O => \N__21398\,
            I => \N__21392\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__21395\,
            I => \N__21389\
        );

    \I__2551\ : InMux
    port map (
            O => \N__21392\,
            I => \N__21385\
        );

    \I__2550\ : Span4Mux_v
    port map (
            O => \N__21389\,
            I => \N__21382\
        );

    \I__2549\ : InMux
    port map (
            O => \N__21388\,
            I => \N__21379\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__21385\,
            I => \N__21376\
        );

    \I__2547\ : Odrv4
    port map (
            O => \N__21382\,
            I => timer_15
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__21379\,
            I => timer_15
        );

    \I__2545\ : Odrv12
    port map (
            O => \N__21376\,
            I => timer_15
        );

    \I__2544\ : InMux
    port map (
            O => \N__21369\,
            I => \bfn_3_23_0_\
        );

    \I__2543\ : InMux
    port map (
            O => \N__21366\,
            I => \N__21363\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__21363\,
            I => \nx.n12951\
        );

    \I__2541\ : InMux
    port map (
            O => \N__21360\,
            I => \N__21357\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__21357\,
            I => \nx.n17\
        );

    \I__2539\ : InMux
    port map (
            O => \N__21354\,
            I => \N__21351\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__21351\,
            I => \N__21347\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__21350\,
            I => \N__21344\
        );

    \I__2536\ : Span4Mux_v
    port map (
            O => \N__21347\,
            I => \N__21341\
        );

    \I__2535\ : InMux
    port map (
            O => \N__21344\,
            I => \N__21338\
        );

    \I__2534\ : Span4Mux_v
    port map (
            O => \N__21341\,
            I => \N__21332\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__21338\,
            I => \N__21332\
        );

    \I__2532\ : InMux
    port map (
            O => \N__21337\,
            I => \N__21329\
        );

    \I__2531\ : Span4Mux_v
    port map (
            O => \N__21332\,
            I => \N__21326\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__21329\,
            I => timer_16
        );

    \I__2529\ : Odrv4
    port map (
            O => \N__21326\,
            I => timer_16
        );

    \I__2528\ : InMux
    port map (
            O => \N__21321\,
            I => \nx.n10437\
        );

    \I__2527\ : InMux
    port map (
            O => \N__21318\,
            I => \N__21315\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__21315\,
            I => \nx.n12953\
        );

    \I__2525\ : InMux
    port map (
            O => \N__21312\,
            I => \nx.n10438\
        );

    \I__2524\ : InMux
    port map (
            O => \N__21309\,
            I => \N__21306\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__21306\,
            I => \nx.n12955\
        );

    \I__2522\ : InMux
    port map (
            O => \N__21303\,
            I => \nx.n10439\
        );

    \I__2521\ : InMux
    port map (
            O => \N__21300\,
            I => \N__21297\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__21297\,
            I => \nx.n12957\
        );

    \I__2519\ : InMux
    port map (
            O => \N__21294\,
            I => \nx.n10440\
        );

    \I__2518\ : InMux
    port map (
            O => \N__21291\,
            I => \N__21288\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__21288\,
            I => \nx.n12959\
        );

    \I__2516\ : InMux
    port map (
            O => \N__21285\,
            I => \nx.n10441\
        );

    \I__2515\ : InMux
    port map (
            O => \N__21282\,
            I => \N__21278\
        );

    \I__2514\ : InMux
    port map (
            O => \N__21281\,
            I => \N__21274\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__21278\,
            I => \N__21271\
        );

    \I__2512\ : InMux
    port map (
            O => \N__21277\,
            I => \N__21268\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__21274\,
            I => \N__21265\
        );

    \I__2510\ : Odrv4
    port map (
            O => \N__21271\,
            I => timer_6
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__21268\,
            I => timer_6
        );

    \I__2508\ : Odrv12
    port map (
            O => \N__21265\,
            I => timer_6
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__21258\,
            I => \N__21255\
        );

    \I__2506\ : InMux
    port map (
            O => \N__21255\,
            I => \N__21252\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__21252\,
            I => \N__21249\
        );

    \I__2504\ : Odrv4
    port map (
            O => \N__21249\,
            I => \nx.n27\
        );

    \I__2503\ : InMux
    port map (
            O => \N__21246\,
            I => \N__21240\
        );

    \I__2502\ : InMux
    port map (
            O => \N__21245\,
            I => \N__21240\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__21240\,
            I => \N__21237\
        );

    \I__2500\ : Span4Mux_s2_h
    port map (
            O => \N__21237\,
            I => \N__21234\
        );

    \I__2499\ : Odrv4
    port map (
            O => \N__21234\,
            I => \nx.one_wire_N_528_6\
        );

    \I__2498\ : InMux
    port map (
            O => \N__21231\,
            I => \nx.n10427\
        );

    \I__2497\ : InMux
    port map (
            O => \N__21228\,
            I => \N__21224\
        );

    \I__2496\ : InMux
    port map (
            O => \N__21227\,
            I => \N__21221\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__21224\,
            I => \N__21218\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__21221\,
            I => \N__21213\
        );

    \I__2493\ : Span4Mux_s2_h
    port map (
            O => \N__21218\,
            I => \N__21213\
        );

    \I__2492\ : Odrv4
    port map (
            O => \N__21213\,
            I => \nx.one_wire_N_528_7\
        );

    \I__2491\ : InMux
    port map (
            O => \N__21210\,
            I => \nx.n10428\
        );

    \I__2490\ : InMux
    port map (
            O => \N__21207\,
            I => \N__21204\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__21204\,
            I => \N__21201\
        );

    \I__2488\ : Odrv4
    port map (
            O => \N__21201\,
            I => \nx.n25\
        );

    \I__2487\ : InMux
    port map (
            O => \N__21198\,
            I => \N__21194\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__21197\,
            I => \N__21191\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__21194\,
            I => \N__21188\
        );

    \I__2484\ : InMux
    port map (
            O => \N__21191\,
            I => \N__21184\
        );

    \I__2483\ : Span4Mux_v
    port map (
            O => \N__21188\,
            I => \N__21181\
        );

    \I__2482\ : InMux
    port map (
            O => \N__21187\,
            I => \N__21178\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__21184\,
            I => \N__21175\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__21181\,
            I => timer_8
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__21178\,
            I => timer_8
        );

    \I__2478\ : Odrv12
    port map (
            O => \N__21175\,
            I => timer_8
        );

    \I__2477\ : InMux
    port map (
            O => \N__21168\,
            I => \N__21163\
        );

    \I__2476\ : InMux
    port map (
            O => \N__21167\,
            I => \N__21160\
        );

    \I__2475\ : InMux
    port map (
            O => \N__21166\,
            I => \N__21157\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__21163\,
            I => \N__21152\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__21160\,
            I => \N__21152\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__21157\,
            I => \N__21149\
        );

    \I__2471\ : Span4Mux_v
    port map (
            O => \N__21152\,
            I => \N__21146\
        );

    \I__2470\ : Span4Mux_s3_h
    port map (
            O => \N__21149\,
            I => \N__21143\
        );

    \I__2469\ : Odrv4
    port map (
            O => \N__21146\,
            I => \nx.one_wire_N_528_8\
        );

    \I__2468\ : Odrv4
    port map (
            O => \N__21143\,
            I => \nx.one_wire_N_528_8\
        );

    \I__2467\ : InMux
    port map (
            O => \N__21138\,
            I => \bfn_3_22_0_\
        );

    \I__2466\ : CascadeMux
    port map (
            O => \N__21135\,
            I => \N__21131\
        );

    \I__2465\ : CascadeMux
    port map (
            O => \N__21134\,
            I => \N__21127\
        );

    \I__2464\ : InMux
    port map (
            O => \N__21131\,
            I => \N__21124\
        );

    \I__2463\ : InMux
    port map (
            O => \N__21130\,
            I => \N__21121\
        );

    \I__2462\ : InMux
    port map (
            O => \N__21127\,
            I => \N__21118\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__21124\,
            I => \N__21115\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__21121\,
            I => \N__21110\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__21118\,
            I => \N__21110\
        );

    \I__2458\ : Span4Mux_s2_h
    port map (
            O => \N__21115\,
            I => \N__21107\
        );

    \I__2457\ : Span4Mux_s2_h
    port map (
            O => \N__21110\,
            I => \N__21104\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__21107\,
            I => \nx.one_wire_N_528_9\
        );

    \I__2455\ : Odrv4
    port map (
            O => \N__21104\,
            I => \nx.one_wire_N_528_9\
        );

    \I__2454\ : InMux
    port map (
            O => \N__21099\,
            I => \nx.n10430\
        );

    \I__2453\ : InMux
    port map (
            O => \N__21096\,
            I => \N__21092\
        );

    \I__2452\ : CascadeMux
    port map (
            O => \N__21095\,
            I => \N__21089\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__21092\,
            I => \N__21086\
        );

    \I__2450\ : InMux
    port map (
            O => \N__21089\,
            I => \N__21083\
        );

    \I__2449\ : Span4Mux_v
    port map (
            O => \N__21086\,
            I => \N__21077\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__21083\,
            I => \N__21077\
        );

    \I__2447\ : InMux
    port map (
            O => \N__21082\,
            I => \N__21074\
        );

    \I__2446\ : Span4Mux_v
    port map (
            O => \N__21077\,
            I => \N__21071\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__21074\,
            I => timer_10
        );

    \I__2444\ : Odrv4
    port map (
            O => \N__21071\,
            I => timer_10
        );

    \I__2443\ : InMux
    port map (
            O => \N__21066\,
            I => \N__21061\
        );

    \I__2442\ : InMux
    port map (
            O => \N__21065\,
            I => \N__21058\
        );

    \I__2441\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21055\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__21061\,
            I => \N__21052\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__21058\,
            I => \N__21049\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__21055\,
            I => \N__21046\
        );

    \I__2437\ : Span12Mux_s2_h
    port map (
            O => \N__21052\,
            I => \N__21043\
        );

    \I__2436\ : Span4Mux_v
    port map (
            O => \N__21049\,
            I => \N__21038\
        );

    \I__2435\ : Span4Mux_s2_h
    port map (
            O => \N__21046\,
            I => \N__21038\
        );

    \I__2434\ : Odrv12
    port map (
            O => \N__21043\,
            I => \nx.one_wire_N_528_10\
        );

    \I__2433\ : Odrv4
    port map (
            O => \N__21038\,
            I => \nx.one_wire_N_528_10\
        );

    \I__2432\ : InMux
    port map (
            O => \N__21033\,
            I => \nx.n10431\
        );

    \I__2431\ : InMux
    port map (
            O => \N__21030\,
            I => \nx.n10432\
        );

    \I__2430\ : InMux
    port map (
            O => \N__21027\,
            I => \N__21024\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__21024\,
            I => \nx.one_wire_N_528_11\
        );

    \I__2428\ : InMux
    port map (
            O => \N__21021\,
            I => \N__21017\
        );

    \I__2427\ : InMux
    port map (
            O => \N__21020\,
            I => \N__21013\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__21017\,
            I => \N__21010\
        );

    \I__2425\ : InMux
    port map (
            O => \N__21016\,
            I => \N__21007\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__21013\,
            I => \N__21004\
        );

    \I__2423\ : Odrv4
    port map (
            O => \N__21010\,
            I => timer_12
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__21007\,
            I => timer_12
        );

    \I__2421\ : Odrv12
    port map (
            O => \N__21004\,
            I => timer_12
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__20997\,
            I => \N__20994\
        );

    \I__2419\ : InMux
    port map (
            O => \N__20994\,
            I => \N__20991\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__20991\,
            I => \N__20988\
        );

    \I__2417\ : Span4Mux_v
    port map (
            O => \N__20988\,
            I => \N__20985\
        );

    \I__2416\ : Span4Mux_s2_h
    port map (
            O => \N__20985\,
            I => \N__20982\
        );

    \I__2415\ : Odrv4
    port map (
            O => \N__20982\,
            I => \nx.n21_adj_620\
        );

    \I__2414\ : InMux
    port map (
            O => \N__20979\,
            I => \nx.n10433\
        );

    \I__2413\ : InMux
    port map (
            O => \N__20976\,
            I => \N__20973\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__20973\,
            I => \nx.n12945\
        );

    \I__2411\ : InMux
    port map (
            O => \N__20970\,
            I => \nx.n10434\
        );

    \I__2410\ : InMux
    port map (
            O => \N__20967\,
            I => \nx.n10508\
        );

    \I__2409\ : InMux
    port map (
            O => \N__20964\,
            I => \nx.n10509\
        );

    \I__2408\ : InMux
    port map (
            O => \N__20961\,
            I => \N__20958\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__20958\,
            I => \N__20955\
        );

    \I__2406\ : Odrv12
    port map (
            O => \N__20955\,
            I => \nx.n32_adj_651\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__20952\,
            I => \N__20948\
        );

    \I__2404\ : InMux
    port map (
            O => \N__20951\,
            I => \N__20944\
        );

    \I__2403\ : InMux
    port map (
            O => \N__20948\,
            I => \N__20941\
        );

    \I__2402\ : InMux
    port map (
            O => \N__20947\,
            I => \N__20938\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__20944\,
            I => \N__20933\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__20941\,
            I => \N__20933\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__20938\,
            I => timer_1
        );

    \I__2398\ : Odrv12
    port map (
            O => \N__20933\,
            I => timer_1
        );

    \I__2397\ : InMux
    port map (
            O => \N__20928\,
            I => \N__20925\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__20925\,
            I => \N__20921\
        );

    \I__2395\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20918\
        );

    \I__2394\ : Span4Mux_s2_h
    port map (
            O => \N__20921\,
            I => \N__20915\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__20918\,
            I => \nx.n11533\
        );

    \I__2392\ : Odrv4
    port map (
            O => \N__20915\,
            I => \nx.n11533\
        );

    \I__2391\ : InMux
    port map (
            O => \N__20910\,
            I => \nx.n10422\
        );

    \I__2390\ : InMux
    port map (
            O => \N__20907\,
            I => \N__20902\
        );

    \I__2389\ : InMux
    port map (
            O => \N__20906\,
            I => \N__20899\
        );

    \I__2388\ : InMux
    port map (
            O => \N__20905\,
            I => \N__20896\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__20902\,
            I => \N__20893\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__20899\,
            I => \nx.one_wire_N_528_2\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__20896\,
            I => \nx.one_wire_N_528_2\
        );

    \I__2384\ : Odrv4
    port map (
            O => \N__20893\,
            I => \nx.one_wire_N_528_2\
        );

    \I__2383\ : InMux
    port map (
            O => \N__20886\,
            I => \nx.n10423\
        );

    \I__2382\ : InMux
    port map (
            O => \N__20883\,
            I => \N__20880\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__20880\,
            I => \nx.n30_adj_598\
        );

    \I__2380\ : CascadeMux
    port map (
            O => \N__20877\,
            I => \N__20873\
        );

    \I__2379\ : InMux
    port map (
            O => \N__20876\,
            I => \N__20870\
        );

    \I__2378\ : InMux
    port map (
            O => \N__20873\,
            I => \N__20866\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__20870\,
            I => \N__20863\
        );

    \I__2376\ : InMux
    port map (
            O => \N__20869\,
            I => \N__20860\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__20866\,
            I => \N__20857\
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__20863\,
            I => timer_3
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__20860\,
            I => timer_3
        );

    \I__2372\ : Odrv12
    port map (
            O => \N__20857\,
            I => timer_3
        );

    \I__2371\ : InMux
    port map (
            O => \N__20850\,
            I => \N__20845\
        );

    \I__2370\ : InMux
    port map (
            O => \N__20849\,
            I => \N__20842\
        );

    \I__2369\ : InMux
    port map (
            O => \N__20848\,
            I => \N__20839\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__20845\,
            I => \N__20836\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__20842\,
            I => \nx.one_wire_N_528_3\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__20839\,
            I => \nx.one_wire_N_528_3\
        );

    \I__2365\ : Odrv4
    port map (
            O => \N__20836\,
            I => \nx.one_wire_N_528_3\
        );

    \I__2364\ : InMux
    port map (
            O => \N__20829\,
            I => \nx.n10424\
        );

    \I__2363\ : InMux
    port map (
            O => \N__20826\,
            I => \N__20823\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__20823\,
            I => \N__20820\
        );

    \I__2361\ : Odrv12
    port map (
            O => \N__20820\,
            I => \nx.n29\
        );

    \I__2360\ : InMux
    port map (
            O => \N__20817\,
            I => \N__20813\
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__20816\,
            I => \N__20810\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__20813\,
            I => \N__20807\
        );

    \I__2357\ : InMux
    port map (
            O => \N__20810\,
            I => \N__20804\
        );

    \I__2356\ : Span4Mux_v
    port map (
            O => \N__20807\,
            I => \N__20798\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__20804\,
            I => \N__20798\
        );

    \I__2354\ : InMux
    port map (
            O => \N__20803\,
            I => \N__20795\
        );

    \I__2353\ : Span4Mux_v
    port map (
            O => \N__20798\,
            I => \N__20792\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__20795\,
            I => timer_4
        );

    \I__2351\ : Odrv4
    port map (
            O => \N__20792\,
            I => timer_4
        );

    \I__2350\ : InMux
    port map (
            O => \N__20787\,
            I => \N__20781\
        );

    \I__2349\ : InMux
    port map (
            O => \N__20786\,
            I => \N__20781\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__20781\,
            I => \N__20778\
        );

    \I__2347\ : Odrv4
    port map (
            O => \N__20778\,
            I => \nx.one_wire_N_528_4\
        );

    \I__2346\ : InMux
    port map (
            O => \N__20775\,
            I => \nx.n10425\
        );

    \I__2345\ : InMux
    port map (
            O => \N__20772\,
            I => \N__20768\
        );

    \I__2344\ : InMux
    port map (
            O => \N__20771\,
            I => \N__20765\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__20768\,
            I => \N__20762\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__20765\,
            I => \N__20758\
        );

    \I__2341\ : Span12Mux_s2_h
    port map (
            O => \N__20762\,
            I => \N__20755\
        );

    \I__2340\ : InMux
    port map (
            O => \N__20761\,
            I => \N__20752\
        );

    \I__2339\ : Span4Mux_v
    port map (
            O => \N__20758\,
            I => \N__20749\
        );

    \I__2338\ : Odrv12
    port map (
            O => \N__20755\,
            I => timer_5
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__20752\,
            I => timer_5
        );

    \I__2336\ : Odrv4
    port map (
            O => \N__20749\,
            I => timer_5
        );

    \I__2335\ : CascadeMux
    port map (
            O => \N__20742\,
            I => \N__20739\
        );

    \I__2334\ : InMux
    port map (
            O => \N__20739\,
            I => \N__20736\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__20736\,
            I => \nx.n28\
        );

    \I__2332\ : InMux
    port map (
            O => \N__20733\,
            I => \N__20730\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__20730\,
            I => \N__20726\
        );

    \I__2330\ : InMux
    port map (
            O => \N__20729\,
            I => \N__20723\
        );

    \I__2329\ : Span12Mux_v
    port map (
            O => \N__20726\,
            I => \N__20720\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__20723\,
            I => \N__20717\
        );

    \I__2327\ : Odrv12
    port map (
            O => \N__20720\,
            I => \nx.one_wire_N_528_5\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__20717\,
            I => \nx.one_wire_N_528_5\
        );

    \I__2325\ : InMux
    port map (
            O => \N__20712\,
            I => \nx.n10426\
        );

    \I__2324\ : InMux
    port map (
            O => \N__20709\,
            I => \nx.n10499\
        );

    \I__2323\ : InMux
    port map (
            O => \N__20706\,
            I => \nx.n10500\
        );

    \I__2322\ : InMux
    port map (
            O => \N__20703\,
            I => \nx.n10501\
        );

    \I__2321\ : InMux
    port map (
            O => \N__20700\,
            I => \bfn_3_20_0_\
        );

    \I__2320\ : InMux
    port map (
            O => \N__20697\,
            I => \nx.n10503\
        );

    \I__2319\ : InMux
    port map (
            O => \N__20694\,
            I => \nx.n10504\
        );

    \I__2318\ : InMux
    port map (
            O => \N__20691\,
            I => \nx.n10505\
        );

    \I__2317\ : InMux
    port map (
            O => \N__20688\,
            I => \nx.n10506\
        );

    \I__2316\ : InMux
    port map (
            O => \N__20685\,
            I => \nx.n10507\
        );

    \I__2315\ : InMux
    port map (
            O => \N__20682\,
            I => \nx.n10490\
        );

    \I__2314\ : InMux
    port map (
            O => \N__20679\,
            I => \nx.n10491\
        );

    \I__2313\ : InMux
    port map (
            O => \N__20676\,
            I => \nx.n10492\
        );

    \I__2312\ : InMux
    port map (
            O => \N__20673\,
            I => \nx.n10493\
        );

    \I__2311\ : InMux
    port map (
            O => \N__20670\,
            I => \bfn_3_19_0_\
        );

    \I__2310\ : InMux
    port map (
            O => \N__20667\,
            I => \nx.n10495\
        );

    \I__2309\ : InMux
    port map (
            O => \N__20664\,
            I => \nx.n10496\
        );

    \I__2308\ : InMux
    port map (
            O => \N__20661\,
            I => \nx.n10497\
        );

    \I__2307\ : InMux
    port map (
            O => \N__20658\,
            I => \nx.n10498\
        );

    \I__2306\ : InMux
    port map (
            O => \N__20655\,
            I => \nx.n10480\
        );

    \I__2305\ : InMux
    port map (
            O => \N__20652\,
            I => \nx.n10481\
        );

    \I__2304\ : InMux
    port map (
            O => \N__20649\,
            I => \nx.n10482\
        );

    \I__2303\ : InMux
    port map (
            O => \N__20646\,
            I => \nx.n10483\
        );

    \I__2302\ : InMux
    port map (
            O => \N__20643\,
            I => \nx.n10484\
        );

    \I__2301\ : InMux
    port map (
            O => \N__20640\,
            I => \nx.n10485\
        );

    \I__2300\ : InMux
    port map (
            O => \N__20637\,
            I => \bfn_3_18_0_\
        );

    \I__2299\ : InMux
    port map (
            O => \N__20634\,
            I => \nx.n10487\
        );

    \I__2298\ : InMux
    port map (
            O => \N__20631\,
            I => \nx.n10488\
        );

    \I__2297\ : InMux
    port map (
            O => \N__20628\,
            I => \nx.n10489\
        );

    \I__2296\ : CascadeMux
    port map (
            O => \N__20625\,
            I => \N__20621\
        );

    \I__2295\ : InMux
    port map (
            O => \N__20624\,
            I => \N__20616\
        );

    \I__2294\ : InMux
    port map (
            O => \N__20621\,
            I => \N__20616\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__20616\,
            I => \nx.n1302\
        );

    \I__2292\ : CascadeMux
    port map (
            O => \N__20613\,
            I => \N__20610\
        );

    \I__2291\ : InMux
    port map (
            O => \N__20610\,
            I => \N__20607\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__20607\,
            I => \nx.n1369\
        );

    \I__2289\ : InMux
    port map (
            O => \N__20604\,
            I => \N__20598\
        );

    \I__2288\ : InMux
    port map (
            O => \N__20603\,
            I => \N__20598\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__20598\,
            I => neo_pixel_transmitter_t0_1
        );

    \I__2286\ : InMux
    port map (
            O => \N__20595\,
            I => \N__20591\
        );

    \I__2285\ : InMux
    port map (
            O => \N__20594\,
            I => \N__20588\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__20591\,
            I => neo_pixel_transmitter_t0_31
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__20588\,
            I => neo_pixel_transmitter_t0_31
        );

    \I__2282\ : InMux
    port map (
            O => \N__20583\,
            I => \N__20579\
        );

    \I__2281\ : InMux
    port map (
            O => \N__20582\,
            I => \N__20576\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__20579\,
            I => neo_pixel_transmitter_t0_4
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__20576\,
            I => neo_pixel_transmitter_t0_4
        );

    \I__2278\ : InMux
    port map (
            O => \N__20571\,
            I => \bfn_3_17_0_\
        );

    \I__2277\ : InMux
    port map (
            O => \N__20568\,
            I => \nx.n10479\
        );

    \I__2276\ : InMux
    port map (
            O => \N__20565\,
            I => \nx.n10573\
        );

    \I__2275\ : InMux
    port map (
            O => \N__20562\,
            I => \nx.n10574\
        );

    \I__2274\ : InMux
    port map (
            O => \N__20559\,
            I => \nx.n10575\
        );

    \I__2273\ : InMux
    port map (
            O => \N__20556\,
            I => \nx.n10576\
        );

    \I__2272\ : InMux
    port map (
            O => \N__20553\,
            I => \nx.n10577\
        );

    \I__2271\ : InMux
    port map (
            O => \N__20550\,
            I => \nx.n10578\
        );

    \I__2270\ : InMux
    port map (
            O => \N__20547\,
            I => \nx.n10579\
        );

    \I__2269\ : InMux
    port map (
            O => \N__20544\,
            I => \bfn_2_32_0_\
        );

    \I__2268\ : CascadeMux
    port map (
            O => \N__20541\,
            I => \N__20538\
        );

    \I__2267\ : InMux
    port map (
            O => \N__20538\,
            I => \N__20534\
        );

    \I__2266\ : InMux
    port map (
            O => \N__20537\,
            I => \N__20531\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__20534\,
            I => \nx.n1301\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__20531\,
            I => \nx.n1301\
        );

    \I__2263\ : InMux
    port map (
            O => \N__20526\,
            I => \nx.n10581\
        );

    \I__2262\ : InMux
    port map (
            O => \N__20523\,
            I => \N__20520\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__20520\,
            I => \nx.n1172\
        );

    \I__2260\ : CascadeMux
    port map (
            O => \N__20517\,
            I => \N__20514\
        );

    \I__2259\ : InMux
    port map (
            O => \N__20514\,
            I => \N__20510\
        );

    \I__2258\ : InMux
    port map (
            O => \N__20513\,
            I => \N__20507\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__20510\,
            I => \nx.n1204\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__20507\,
            I => \nx.n1204\
        );

    \I__2255\ : InMux
    port map (
            O => \N__20502\,
            I => \N__20499\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__20499\,
            I => \nx.n1271\
        );

    \I__2253\ : CascadeMux
    port map (
            O => \N__20496\,
            I => \nx.n1204_cascade_\
        );

    \I__2252\ : InMux
    port map (
            O => \N__20493\,
            I => \N__20490\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__20490\,
            I => \nx.n11_adj_624\
        );

    \I__2250\ : CascadeMux
    port map (
            O => \N__20487\,
            I => \N__20484\
        );

    \I__2249\ : InMux
    port map (
            O => \N__20484\,
            I => \N__20481\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__20481\,
            I => \nx.n13\
        );

    \I__2247\ : InMux
    port map (
            O => \N__20478\,
            I => \N__20474\
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__20477\,
            I => \N__20471\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__20474\,
            I => \N__20468\
        );

    \I__2244\ : InMux
    port map (
            O => \N__20471\,
            I => \N__20465\
        );

    \I__2243\ : Span4Mux_h
    port map (
            O => \N__20468\,
            I => \N__20462\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__20465\,
            I => \nx.n1206\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__20462\,
            I => \nx.n1206\
        );

    \I__2240\ : InMux
    port map (
            O => \N__20457\,
            I => \N__20454\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__20454\,
            I => \nx.n1275\
        );

    \I__2238\ : CascadeMux
    port map (
            O => \N__20451\,
            I => \nx.n1235_cascade_\
        );

    \I__2237\ : CascadeMux
    port map (
            O => \N__20448\,
            I => \N__20444\
        );

    \I__2236\ : InMux
    port map (
            O => \N__20447\,
            I => \N__20441\
        );

    \I__2235\ : InMux
    port map (
            O => \N__20444\,
            I => \N__20438\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__20441\,
            I => \nx.n1208\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__20438\,
            I => \nx.n1208\
        );

    \I__2232\ : InMux
    port map (
            O => \N__20433\,
            I => \N__20430\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__20430\,
            I => \nx.n1175\
        );

    \I__2230\ : InMux
    port map (
            O => \N__20427\,
            I => \N__20420\
        );

    \I__2229\ : CascadeMux
    port map (
            O => \N__20426\,
            I => \N__20416\
        );

    \I__2228\ : CascadeMux
    port map (
            O => \N__20425\,
            I => \N__20413\
        );

    \I__2227\ : InMux
    port map (
            O => \N__20424\,
            I => \N__20407\
        );

    \I__2226\ : InMux
    port map (
            O => \N__20423\,
            I => \N__20407\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__20420\,
            I => \N__20404\
        );

    \I__2224\ : InMux
    port map (
            O => \N__20419\,
            I => \N__20401\
        );

    \I__2223\ : InMux
    port map (
            O => \N__20416\,
            I => \N__20394\
        );

    \I__2222\ : InMux
    port map (
            O => \N__20413\,
            I => \N__20394\
        );

    \I__2221\ : InMux
    port map (
            O => \N__20412\,
            I => \N__20394\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__20407\,
            I => \nx.n1136\
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__20404\,
            I => \nx.n1136\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__20401\,
            I => \nx.n1136\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__20394\,
            I => \nx.n1136\
        );

    \I__2216\ : CascadeMux
    port map (
            O => \N__20385\,
            I => \N__20382\
        );

    \I__2215\ : InMux
    port map (
            O => \N__20382\,
            I => \N__20378\
        );

    \I__2214\ : InMux
    port map (
            O => \N__20381\,
            I => \N__20375\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__20378\,
            I => \nx.n1207\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__20375\,
            I => \nx.n1207\
        );

    \I__2211\ : InMux
    port map (
            O => \N__20370\,
            I => \N__20367\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__20367\,
            I => \nx.n1274\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__20364\,
            I => \nx.n1207_cascade_\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__20361\,
            I => \nx.n1306_cascade_\
        );

    \I__2207\ : InMux
    port map (
            O => \N__20358\,
            I => \N__20355\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__20355\,
            I => \N__20352\
        );

    \I__2205\ : Odrv4
    port map (
            O => \N__20352\,
            I => \nx.n10_adj_626\
        );

    \I__2204\ : InMux
    port map (
            O => \N__20349\,
            I => \bfn_2_31_0_\
        );

    \I__2203\ : InMux
    port map (
            O => \N__20346\,
            I => \N__20343\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__20343\,
            I => \nx.n1177\
        );

    \I__2201\ : InMux
    port map (
            O => \N__20340\,
            I => \bfn_2_29_0_\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__20337\,
            I => \N__20332\
        );

    \I__2199\ : InMux
    port map (
            O => \N__20336\,
            I => \N__20327\
        );

    \I__2198\ : InMux
    port map (
            O => \N__20335\,
            I => \N__20327\
        );

    \I__2197\ : InMux
    port map (
            O => \N__20332\,
            I => \N__20324\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__20327\,
            I => \nx.n1109\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__20324\,
            I => \nx.n1109\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__20319\,
            I => \N__20316\
        );

    \I__2193\ : InMux
    port map (
            O => \N__20316\,
            I => \N__20313\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__20313\,
            I => \N__20310\
        );

    \I__2191\ : Odrv4
    port map (
            O => \N__20310\,
            I => \nx.n1176\
        );

    \I__2190\ : InMux
    port map (
            O => \N__20307\,
            I => \nx.n10461\
        );

    \I__2189\ : InMux
    port map (
            O => \N__20304\,
            I => \nx.n10462\
        );

    \I__2188\ : InMux
    port map (
            O => \N__20301\,
            I => \N__20298\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__20298\,
            I => \N__20295\
        );

    \I__2186\ : Odrv4
    port map (
            O => \N__20295\,
            I => \nx.n1174\
        );

    \I__2185\ : InMux
    port map (
            O => \N__20292\,
            I => \nx.n10463\
        );

    \I__2184\ : InMux
    port map (
            O => \N__20289\,
            I => \nx.n10464\
        );

    \I__2183\ : InMux
    port map (
            O => \N__20286\,
            I => \nx.n10465\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__20283\,
            I => \N__20280\
        );

    \I__2181\ : InMux
    port map (
            O => \N__20280\,
            I => \N__20277\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__20277\,
            I => \nx.n1171\
        );

    \I__2179\ : InMux
    port map (
            O => \N__20274\,
            I => \nx.n10466\
        );

    \I__2178\ : InMux
    port map (
            O => \N__20271\,
            I => \nx.n10467\
        );

    \I__2177\ : InMux
    port map (
            O => \N__20268\,
            I => \N__20265\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__20265\,
            I => \N__20262\
        );

    \I__2175\ : Span4Mux_s1_v
    port map (
            O => \N__20262\,
            I => \N__20258\
        );

    \I__2174\ : InMux
    port map (
            O => \N__20261\,
            I => \N__20255\
        );

    \I__2173\ : Odrv4
    port map (
            O => \N__20258\,
            I => \nx.n1202\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__20255\,
            I => \nx.n1202\
        );

    \I__2171\ : CascadeMux
    port map (
            O => \N__20250\,
            I => \N__20247\
        );

    \I__2170\ : InMux
    port map (
            O => \N__20247\,
            I => \N__20244\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__20244\,
            I => \nx.n1173\
        );

    \I__2168\ : InMux
    port map (
            O => \N__20241\,
            I => \N__20238\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__20238\,
            I => \N__20235\
        );

    \I__2166\ : Odrv4
    port map (
            O => \N__20235\,
            I => \nx.n3151\
        );

    \I__2165\ : InMux
    port map (
            O => \N__20232\,
            I => \N__20229\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__20229\,
            I => \N__20226\
        );

    \I__2163\ : Odrv12
    port map (
            O => \N__20226\,
            I => \nx.n61\
        );

    \I__2162\ : CascadeMux
    port map (
            O => \N__20223\,
            I => \N__20218\
        );

    \I__2161\ : InMux
    port map (
            O => \N__20222\,
            I => \N__20215\
        );

    \I__2160\ : InMux
    port map (
            O => \N__20221\,
            I => \N__20212\
        );

    \I__2159\ : InMux
    port map (
            O => \N__20218\,
            I => \N__20209\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__20215\,
            I => \N__20204\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__20212\,
            I => \N__20204\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__20209\,
            I => \nx.n3099\
        );

    \I__2155\ : Odrv4
    port map (
            O => \N__20204\,
            I => \nx.n3099\
        );

    \I__2154\ : InMux
    port map (
            O => \N__20199\,
            I => \N__20196\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__20196\,
            I => \N__20193\
        );

    \I__2152\ : Span4Mux_v
    port map (
            O => \N__20193\,
            I => \N__20190\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__20190\,
            I => neopxl_color_prev_7
        );

    \I__2150\ : InMux
    port map (
            O => \N__20187\,
            I => \N__20184\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__20184\,
            I => \nx.n54\
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__20181\,
            I => \nx.n43_adj_709_cascade_\
        );

    \I__2147\ : InMux
    port map (
            O => \N__20178\,
            I => \N__20175\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__20175\,
            I => \nx.n49_adj_710\
        );

    \I__2145\ : InMux
    port map (
            O => \N__20172\,
            I => \N__20168\
        );

    \I__2144\ : InMux
    port map (
            O => \N__20171\,
            I => \N__20165\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__20168\,
            I => \N__20158\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__20165\,
            I => \N__20158\
        );

    \I__2141\ : InMux
    port map (
            O => \N__20164\,
            I => \N__20153\
        );

    \I__2140\ : InMux
    port map (
            O => \N__20163\,
            I => \N__20153\
        );

    \I__2139\ : Span4Mux_v
    port map (
            O => \N__20158\,
            I => \N__20148\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__20153\,
            I => \N__20148\
        );

    \I__2137\ : Span4Mux_v
    port map (
            O => \N__20148\,
            I => \N__20145\
        );

    \I__2136\ : Odrv4
    port map (
            O => \N__20145\,
            I => \state_3_N_377_1\
        );

    \I__2135\ : InMux
    port map (
            O => \N__20142\,
            I => \N__20139\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__20139\,
            I => \N__20134\
        );

    \I__2133\ : InMux
    port map (
            O => \N__20138\,
            I => \N__20131\
        );

    \I__2132\ : InMux
    port map (
            O => \N__20137\,
            I => \N__20128\
        );

    \I__2131\ : Span4Mux_s1_h
    port map (
            O => \N__20134\,
            I => \N__20125\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__20131\,
            I => \nx.n3084\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__20128\,
            I => \nx.n3084\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__20125\,
            I => \nx.n3084\
        );

    \I__2127\ : InMux
    port map (
            O => \N__20118\,
            I => \N__20115\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__20115\,
            I => \nx.n3174\
        );

    \I__2125\ : InMux
    port map (
            O => \N__20112\,
            I => \N__20109\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__20109\,
            I => \nx.n23_adj_700\
        );

    \I__2123\ : CascadeMux
    port map (
            O => \N__20106\,
            I => \N__20103\
        );

    \I__2122\ : InMux
    port map (
            O => \N__20103\,
            I => \N__20098\
        );

    \I__2121\ : InMux
    port map (
            O => \N__20102\,
            I => \N__20095\
        );

    \I__2120\ : InMux
    port map (
            O => \N__20101\,
            I => \N__20092\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__20098\,
            I => \nx.n3107\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__20095\,
            I => \nx.n3107\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__20092\,
            I => \nx.n3107\
        );

    \I__2116\ : InMux
    port map (
            O => \N__20085\,
            I => \N__20082\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__20082\,
            I => \nx.n3162\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__20079\,
            I => \nx.n12327_cascade_\
        );

    \I__2113\ : InMux
    port map (
            O => \N__20076\,
            I => \N__20072\
        );

    \I__2112\ : CascadeMux
    port map (
            O => \N__20075\,
            I => \N__20069\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__20072\,
            I => \N__20066\
        );

    \I__2110\ : InMux
    port map (
            O => \N__20069\,
            I => \N__20063\
        );

    \I__2109\ : Span4Mux_v
    port map (
            O => \N__20066\,
            I => \N__20059\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__20063\,
            I => \N__20056\
        );

    \I__2107\ : InMux
    port map (
            O => \N__20062\,
            I => \N__20053\
        );

    \I__2106\ : Odrv4
    port map (
            O => \N__20059\,
            I => \nx.n3095\
        );

    \I__2105\ : Odrv12
    port map (
            O => \N__20056\,
            I => \nx.n3095\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__20053\,
            I => \nx.n3095\
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__20046\,
            I => \N__20043\
        );

    \I__2102\ : InMux
    port map (
            O => \N__20043\,
            I => \N__20040\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__20040\,
            I => \nx.n3166\
        );

    \I__2100\ : InMux
    port map (
            O => \N__20037\,
            I => \N__20034\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__20034\,
            I => \nx.n3177\
        );

    \I__2098\ : InMux
    port map (
            O => \N__20031\,
            I => \N__20028\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__20028\,
            I => \N__20024\
        );

    \I__2096\ : InMux
    port map (
            O => \N__20027\,
            I => \N__20021\
        );

    \I__2095\ : Odrv12
    port map (
            O => \N__20024\,
            I => \nx.n3209\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__20021\,
            I => \nx.n3209\
        );

    \I__2093\ : InMux
    port map (
            O => \N__20016\,
            I => \N__20013\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__20013\,
            I => \nx.n3171\
        );

    \I__2091\ : InMux
    port map (
            O => \N__20010\,
            I => \N__20007\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__20007\,
            I => \nx.n3175\
        );

    \I__2089\ : InMux
    port map (
            O => \N__20004\,
            I => \N__19999\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__20003\,
            I => \N__19996\
        );

    \I__2087\ : InMux
    port map (
            O => \N__20002\,
            I => \N__19993\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__19999\,
            I => \N__19990\
        );

    \I__2085\ : InMux
    port map (
            O => \N__19996\,
            I => \N__19987\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__19993\,
            I => \nx.n3108\
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__19990\,
            I => \nx.n3108\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__19987\,
            I => \nx.n3108\
        );

    \I__2081\ : InMux
    port map (
            O => \N__19980\,
            I => \N__19977\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__19977\,
            I => \nx.n3165\
        );

    \I__2079\ : InMux
    port map (
            O => \N__19974\,
            I => \N__19970\
        );

    \I__2078\ : InMux
    port map (
            O => \N__19973\,
            I => \N__19967\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__19970\,
            I => \N__19961\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__19967\,
            I => \N__19961\
        );

    \I__2075\ : InMux
    port map (
            O => \N__19966\,
            I => \N__19958\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__19961\,
            I => \nx.n3098\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__19958\,
            I => \nx.n3098\
        );

    \I__2072\ : CascadeMux
    port map (
            O => \N__19953\,
            I => \nx.n13_adj_696_cascade_\
        );

    \I__2071\ : InMux
    port map (
            O => \N__19950\,
            I => \N__19947\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__19947\,
            I => \nx.n31_adj_702\
        );

    \I__2069\ : InMux
    port map (
            O => \N__19944\,
            I => \N__19941\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__19941\,
            I => \nx.n21_adj_701\
        );

    \I__2067\ : CascadeMux
    port map (
            O => \N__19938\,
            I => \nx.n12325_cascade_\
        );

    \I__2066\ : InMux
    port map (
            O => \N__19935\,
            I => \N__19932\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__19932\,
            I => \nx.n12339\
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__19929\,
            I => \N__19926\
        );

    \I__2063\ : InMux
    port map (
            O => \N__19926\,
            I => \N__19923\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__19923\,
            I => \nx.n12347\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__19920\,
            I => \N__19917\
        );

    \I__2060\ : InMux
    port map (
            O => \N__19917\,
            I => \N__19912\
        );

    \I__2059\ : InMux
    port map (
            O => \N__19916\,
            I => \N__19907\
        );

    \I__2058\ : InMux
    port map (
            O => \N__19915\,
            I => \N__19907\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__19912\,
            I => \N__19904\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__19907\,
            I => \nx.n3103\
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__19904\,
            I => \nx.n3103\
        );

    \I__2054\ : InMux
    port map (
            O => \N__19899\,
            I => \N__19895\
        );

    \I__2053\ : InMux
    port map (
            O => \N__19898\,
            I => \N__19892\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__19895\,
            I => \N__19889\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__19892\,
            I => \N__19886\
        );

    \I__2050\ : Odrv4
    port map (
            O => \N__19889\,
            I => \nx.n3097\
        );

    \I__2049\ : Odrv4
    port map (
            O => \N__19886\,
            I => \nx.n3097\
        );

    \I__2048\ : InMux
    port map (
            O => \N__19881\,
            I => \N__19878\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__19878\,
            I => \N__19875\
        );

    \I__2046\ : Odrv4
    port map (
            O => \N__19875\,
            I => \nx.n3164\
        );

    \I__2045\ : CascadeMux
    port map (
            O => \N__19872\,
            I => \nx.n3097_cascade_\
        );

    \I__2044\ : InMux
    port map (
            O => \N__19869\,
            I => \N__19866\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__19866\,
            I => \N__19863\
        );

    \I__2042\ : Odrv4
    port map (
            O => \N__19863\,
            I => \nx.n3168\
        );

    \I__2041\ : CascadeMux
    port map (
            O => \N__19860\,
            I => \nx.n35_adj_699_cascade_\
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__19857\,
            I => \N__19854\
        );

    \I__2039\ : InMux
    port map (
            O => \N__19854\,
            I => \N__19851\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__19851\,
            I => \N__19847\
        );

    \I__2037\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19843\
        );

    \I__2036\ : Span4Mux_v
    port map (
            O => \N__19847\,
            I => \N__19840\
        );

    \I__2035\ : InMux
    port map (
            O => \N__19846\,
            I => \N__19837\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__19843\,
            I => \nx.n3101\
        );

    \I__2033\ : Odrv4
    port map (
            O => \N__19840\,
            I => \nx.n3101\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__19837\,
            I => \nx.n3101\
        );

    \I__2031\ : InMux
    port map (
            O => \N__19830\,
            I => \N__19827\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__19827\,
            I => \nx.n12337\
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__19824\,
            I => \N__19819\
        );

    \I__2028\ : InMux
    port map (
            O => \N__19823\,
            I => \N__19816\
        );

    \I__2027\ : InMux
    port map (
            O => \N__19822\,
            I => \N__19813\
        );

    \I__2026\ : InMux
    port map (
            O => \N__19819\,
            I => \N__19810\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__19816\,
            I => \nx.n3109\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__19813\,
            I => \nx.n3109\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__19810\,
            I => \nx.n3109\
        );

    \I__2022\ : InMux
    port map (
            O => \N__19803\,
            I => \N__19800\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__19800\,
            I => \nx.n12349\
        );

    \I__2020\ : CascadeMux
    port map (
            O => \N__19797\,
            I => \N__19794\
        );

    \I__2019\ : InMux
    port map (
            O => \N__19794\,
            I => \N__19790\
        );

    \I__2018\ : InMux
    port map (
            O => \N__19793\,
            I => \N__19787\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__19790\,
            I => \N__19784\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__19787\,
            I => \N__19779\
        );

    \I__2015\ : Span4Mux_v
    port map (
            O => \N__19784\,
            I => \N__19779\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__19779\,
            I => \nx.n3096\
        );

    \I__2013\ : CascadeMux
    port map (
            O => \N__19776\,
            I => \nx.n3096_cascade_\
        );

    \I__2012\ : InMux
    port map (
            O => \N__19773\,
            I => \N__19770\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__19770\,
            I => \N__19767\
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__19767\,
            I => \nx.n47_adj_694\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__19764\,
            I => \N__19761\
        );

    \I__2008\ : InMux
    port map (
            O => \N__19761\,
            I => \N__19758\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__19758\,
            I => \nx.n45\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__19755\,
            I => \nx.n49_cascade_\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__19752\,
            I => \nx.n3017_cascade_\
        );

    \I__2004\ : InMux
    port map (
            O => \N__19749\,
            I => \N__19745\
        );

    \I__2003\ : InMux
    port map (
            O => \N__19748\,
            I => \N__19742\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__19745\,
            I => \N__19739\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__19742\,
            I => \N__19736\
        );

    \I__2000\ : Span4Mux_v
    port map (
            O => \N__19739\,
            I => \N__19733\
        );

    \I__1999\ : Odrv4
    port map (
            O => \N__19736\,
            I => \nx.n3086\
        );

    \I__1998\ : Odrv4
    port map (
            O => \N__19733\,
            I => \nx.n3086\
        );

    \I__1997\ : InMux
    port map (
            O => \N__19728\,
            I => \N__19724\
        );

    \I__1996\ : InMux
    port map (
            O => \N__19727\,
            I => \N__19721\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__19724\,
            I => \N__19718\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__19721\,
            I => \N__19714\
        );

    \I__1993\ : Span4Mux_v
    port map (
            O => \N__19718\,
            I => \N__19711\
        );

    \I__1992\ : InMux
    port map (
            O => \N__19717\,
            I => \N__19708\
        );

    \I__1991\ : Odrv4
    port map (
            O => \N__19714\,
            I => \nx.n3087\
        );

    \I__1990\ : Odrv4
    port map (
            O => \N__19711\,
            I => \nx.n3087\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__19708\,
            I => \nx.n3087\
        );

    \I__1988\ : CascadeMux
    port map (
            O => \N__19701\,
            I => \nx.n3086_cascade_\
        );

    \I__1987\ : InMux
    port map (
            O => \N__19698\,
            I => \N__19695\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__19695\,
            I => \N__19691\
        );

    \I__1985\ : InMux
    port map (
            O => \N__19694\,
            I => \N__19687\
        );

    \I__1984\ : Span4Mux_v
    port map (
            O => \N__19691\,
            I => \N__19684\
        );

    \I__1983\ : InMux
    port map (
            O => \N__19690\,
            I => \N__19681\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__19687\,
            I => \nx.n3085\
        );

    \I__1981\ : Odrv4
    port map (
            O => \N__19684\,
            I => \nx.n3085\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__19681\,
            I => \nx.n3085\
        );

    \I__1979\ : InMux
    port map (
            O => \N__19674\,
            I => \N__19671\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__19671\,
            I => \nx.n42_adj_689\
        );

    \I__1977\ : CascadeMux
    port map (
            O => \N__19668\,
            I => \N__19665\
        );

    \I__1976\ : InMux
    port map (
            O => \N__19665\,
            I => \N__19662\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__19662\,
            I => \nx.color_bit_N_571_4\
        );

    \I__1974\ : InMux
    port map (
            O => \N__19659\,
            I => \N__19656\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__19656\,
            I => \nx.n13158\
        );

    \I__1972\ : InMux
    port map (
            O => \N__19653\,
            I => \N__19650\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__19650\,
            I => \nx.n59\
        );

    \I__1970\ : CascadeMux
    port map (
            O => \N__19647\,
            I => \N__19644\
        );

    \I__1969\ : InMux
    port map (
            O => \N__19644\,
            I => \N__19641\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__19641\,
            I => \nx.n12371\
        );

    \I__1967\ : InMux
    port map (
            O => \N__19638\,
            I => \N__19635\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__19635\,
            I => \N__19632\
        );

    \I__1965\ : Span4Mux_v
    port map (
            O => \N__19632\,
            I => \N__19629\
        );

    \I__1964\ : Odrv4
    port map (
            O => \N__19629\,
            I => \nx.n13042\
        );

    \I__1963\ : InMux
    port map (
            O => \N__19626\,
            I => \N__19623\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__19623\,
            I => \nx.n10947\
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__19620\,
            I => \nx.n10947_cascade_\
        );

    \I__1960\ : InMux
    port map (
            O => \N__19617\,
            I => \N__19611\
        );

    \I__1959\ : InMux
    port map (
            O => \N__19616\,
            I => \N__19611\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__19611\,
            I => \nx.n10975\
        );

    \I__1957\ : CascadeMux
    port map (
            O => \N__19608\,
            I => \nx.n3008_cascade_\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__19605\,
            I => \N__19600\
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__19604\,
            I => \N__19597\
        );

    \I__1954\ : InMux
    port map (
            O => \N__19603\,
            I => \N__19587\
        );

    \I__1953\ : InMux
    port map (
            O => \N__19600\,
            I => \N__19587\
        );

    \I__1952\ : InMux
    port map (
            O => \N__19597\,
            I => \N__19587\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__19596\,
            I => \N__19583\
        );

    \I__1950\ : InMux
    port map (
            O => \N__19595\,
            I => \N__19575\
        );

    \I__1949\ : InMux
    port map (
            O => \N__19594\,
            I => \N__19575\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__19587\,
            I => \N__19571\
        );

    \I__1947\ : InMux
    port map (
            O => \N__19586\,
            I => \N__19566\
        );

    \I__1946\ : InMux
    port map (
            O => \N__19583\,
            I => \N__19566\
        );

    \I__1945\ : InMux
    port map (
            O => \N__19582\,
            I => \N__19561\
        );

    \I__1944\ : InMux
    port map (
            O => \N__19581\,
            I => \N__19556\
        );

    \I__1943\ : InMux
    port map (
            O => \N__19580\,
            I => \N__19556\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__19575\,
            I => \N__19553\
        );

    \I__1941\ : InMux
    port map (
            O => \N__19574\,
            I => \N__19550\
        );

    \I__1940\ : Span4Mux_v
    port map (
            O => \N__19571\,
            I => \N__19545\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__19566\,
            I => \N__19545\
        );

    \I__1938\ : InMux
    port map (
            O => \N__19565\,
            I => \N__19540\
        );

    \I__1937\ : InMux
    port map (
            O => \N__19564\,
            I => \N__19540\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__19561\,
            I => state_0_adj_727
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__19556\,
            I => state_0_adj_727
        );

    \I__1934\ : Odrv4
    port map (
            O => \N__19553\,
            I => state_0_adj_727
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__19550\,
            I => state_0_adj_727
        );

    \I__1932\ : Odrv4
    port map (
            O => \N__19545\,
            I => state_0_adj_727
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__19540\,
            I => state_0_adj_727
        );

    \I__1930\ : InMux
    port map (
            O => \N__19527\,
            I => \N__19524\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__19524\,
            I => \N__19520\
        );

    \I__1928\ : InMux
    port map (
            O => \N__19523\,
            I => \N__19517\
        );

    \I__1927\ : Span4Mux_v
    port map (
            O => \N__19520\,
            I => \N__19505\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__19517\,
            I => \N__19505\
        );

    \I__1925\ : CascadeMux
    port map (
            O => \N__19516\,
            I => \N__19501\
        );

    \I__1924\ : CascadeMux
    port map (
            O => \N__19515\,
            I => \N__19497\
        );

    \I__1923\ : InMux
    port map (
            O => \N__19514\,
            I => \N__19492\
        );

    \I__1922\ : InMux
    port map (
            O => \N__19513\,
            I => \N__19489\
        );

    \I__1921\ : InMux
    port map (
            O => \N__19512\,
            I => \N__19484\
        );

    \I__1920\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19484\
        );

    \I__1919\ : InMux
    port map (
            O => \N__19510\,
            I => \N__19481\
        );

    \I__1918\ : Span4Mux_v
    port map (
            O => \N__19505\,
            I => \N__19476\
        );

    \I__1917\ : InMux
    port map (
            O => \N__19504\,
            I => \N__19473\
        );

    \I__1916\ : InMux
    port map (
            O => \N__19501\,
            I => \N__19470\
        );

    \I__1915\ : InMux
    port map (
            O => \N__19500\,
            I => \N__19461\
        );

    \I__1914\ : InMux
    port map (
            O => \N__19497\,
            I => \N__19461\
        );

    \I__1913\ : InMux
    port map (
            O => \N__19496\,
            I => \N__19461\
        );

    \I__1912\ : InMux
    port map (
            O => \N__19495\,
            I => \N__19461\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__19492\,
            I => \N__19452\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__19489\,
            I => \N__19452\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__19484\,
            I => \N__19452\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__19481\,
            I => \N__19452\
        );

    \I__1907\ : InMux
    port map (
            O => \N__19480\,
            I => \N__19449\
        );

    \I__1906\ : InMux
    port map (
            O => \N__19479\,
            I => \N__19446\
        );

    \I__1905\ : Odrv4
    port map (
            O => \N__19476\,
            I => state_1_adj_726
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__19473\,
            I => state_1_adj_726
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__19470\,
            I => state_1_adj_726
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__19461\,
            I => state_1_adj_726
        );

    \I__1901\ : Odrv4
    port map (
            O => \N__19452\,
            I => state_1_adj_726
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__19449\,
            I => state_1_adj_726
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__19446\,
            I => state_1_adj_726
        );

    \I__1898\ : CEMux
    port map (
            O => \N__19431\,
            I => \N__19427\
        );

    \I__1897\ : InMux
    port map (
            O => \N__19430\,
            I => \N__19424\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__19427\,
            I => n7239
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__19424\,
            I => n7239
        );

    \I__1894\ : SRMux
    port map (
            O => \N__19419\,
            I => \N__19416\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__19416\,
            I => \N__19413\
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__19413\,
            I => \nx.n7392\
        );

    \I__1891\ : InMux
    port map (
            O => \N__19410\,
            I => \N__19407\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__19407\,
            I => \nx.n13155\
        );

    \I__1889\ : CascadeMux
    port map (
            O => \N__19404\,
            I => \nx.n13456_cascade_\
        );

    \I__1888\ : InMux
    port map (
            O => \N__19401\,
            I => \N__19398\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__19398\,
            I => \nx.n13156\
        );

    \I__1886\ : InMux
    port map (
            O => \N__19395\,
            I => \N__19392\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__19392\,
            I => \nx.n13459\
        );

    \I__1884\ : InMux
    port map (
            O => \N__19389\,
            I => \N__19382\
        );

    \I__1883\ : InMux
    port map (
            O => \N__19388\,
            I => \N__19382\
        );

    \I__1882\ : InMux
    port map (
            O => \N__19387\,
            I => \N__19379\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__19382\,
            I => \N__19374\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__19379\,
            I => \N__19371\
        );

    \I__1879\ : InMux
    port map (
            O => \N__19378\,
            I => \N__19366\
        );

    \I__1878\ : InMux
    port map (
            O => \N__19377\,
            I => \N__19366\
        );

    \I__1877\ : Span4Mux_v
    port map (
            O => \N__19374\,
            I => \N__19363\
        );

    \I__1876\ : Span4Mux_s1_h
    port map (
            O => \N__19371\,
            I => \N__19358\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__19366\,
            I => \N__19358\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__19363\,
            I => \nx.n4_adj_642\
        );

    \I__1873\ : Odrv4
    port map (
            O => \N__19358\,
            I => \nx.n4_adj_642\
        );

    \I__1872\ : InMux
    port map (
            O => \N__19353\,
            I => \N__19349\
        );

    \I__1871\ : InMux
    port map (
            O => \N__19352\,
            I => \N__19346\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__19349\,
            I => neo_pixel_transmitter_t0_26
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__19346\,
            I => neo_pixel_transmitter_t0_26
        );

    \I__1868\ : InMux
    port map (
            O => \N__19341\,
            I => \N__19337\
        );

    \I__1867\ : InMux
    port map (
            O => \N__19340\,
            I => \N__19334\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__19337\,
            I => neo_pixel_transmitter_t0_16
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__19334\,
            I => neo_pixel_transmitter_t0_16
        );

    \I__1864\ : InMux
    port map (
            O => \N__19329\,
            I => \N__19326\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__19326\,
            I => neopxl_color_prev_5
        );

    \I__1862\ : InMux
    port map (
            O => \N__19323\,
            I => \N__19320\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__19320\,
            I => \N__19317\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__19317\,
            I => n10_adj_776
        );

    \I__1859\ : InMux
    port map (
            O => \N__19314\,
            I => \N__19308\
        );

    \I__1858\ : InMux
    port map (
            O => \N__19313\,
            I => \N__19308\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__19308\,
            I => neo_pixel_transmitter_t0_3
        );

    \I__1856\ : InMux
    port map (
            O => \N__19305\,
            I => \N__19302\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__19302\,
            I => n12_adj_774
        );

    \I__1854\ : InMux
    port map (
            O => \N__19299\,
            I => \N__19295\
        );

    \I__1853\ : InMux
    port map (
            O => \N__19298\,
            I => \N__19292\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__19295\,
            I => neo_pixel_transmitter_t0_12
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__19292\,
            I => neo_pixel_transmitter_t0_12
        );

    \I__1850\ : CascadeMux
    port map (
            O => \N__19287\,
            I => \N__19283\
        );

    \I__1849\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19278\
        );

    \I__1848\ : InMux
    port map (
            O => \N__19283\,
            I => \N__19273\
        );

    \I__1847\ : InMux
    port map (
            O => \N__19282\,
            I => \N__19273\
        );

    \I__1846\ : InMux
    port map (
            O => \N__19281\,
            I => \N__19268\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__19278\,
            I => \N__19257\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__19273\,
            I => \N__19257\
        );

    \I__1843\ : InMux
    port map (
            O => \N__19272\,
            I => \N__19254\
        );

    \I__1842\ : InMux
    port map (
            O => \N__19271\,
            I => \N__19251\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__19268\,
            I => \N__19248\
        );

    \I__1840\ : InMux
    port map (
            O => \N__19267\,
            I => \N__19243\
        );

    \I__1839\ : InMux
    port map (
            O => \N__19266\,
            I => \N__19243\
        );

    \I__1838\ : InMux
    port map (
            O => \N__19265\,
            I => \N__19240\
        );

    \I__1837\ : InMux
    port map (
            O => \N__19264\,
            I => \N__19237\
        );

    \I__1836\ : InMux
    port map (
            O => \N__19263\,
            I => \N__19232\
        );

    \I__1835\ : InMux
    port map (
            O => \N__19262\,
            I => \N__19232\
        );

    \I__1834\ : Sp12to4
    port map (
            O => \N__19257\,
            I => \N__19227\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__19254\,
            I => \N__19227\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__19251\,
            I => \nx.neo_pixel_transmitter_done\
        );

    \I__1831\ : Odrv4
    port map (
            O => \N__19248\,
            I => \nx.neo_pixel_transmitter_done\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__19243\,
            I => \nx.neo_pixel_transmitter_done\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__19240\,
            I => \nx.neo_pixel_transmitter_done\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__19237\,
            I => \nx.neo_pixel_transmitter_done\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__19232\,
            I => \nx.neo_pixel_transmitter_done\
        );

    \I__1826\ : Odrv12
    port map (
            O => \N__19227\,
            I => \nx.neo_pixel_transmitter_done\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__19212\,
            I => \nx.n11487_cascade_\
        );

    \I__1824\ : InMux
    port map (
            O => \N__19209\,
            I => \N__19206\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__19206\,
            I => \nx.n103\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__19203\,
            I => \N__19200\
        );

    \I__1821\ : InMux
    port map (
            O => \N__19200\,
            I => \N__19197\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__19197\,
            I => \N__19194\
        );

    \I__1819\ : Span4Mux_v
    port map (
            O => \N__19194\,
            I => \N__19191\
        );

    \I__1818\ : Odrv4
    port map (
            O => \N__19191\,
            I => n9_adj_777
        );

    \I__1817\ : InMux
    port map (
            O => \N__19188\,
            I => \N__19185\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__19185\,
            I => neopxl_color_prev_4
        );

    \I__1815\ : InMux
    port map (
            O => \N__19182\,
            I => \N__19178\
        );

    \I__1814\ : CascadeMux
    port map (
            O => \N__19181\,
            I => \N__19175\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__19178\,
            I => \N__19170\
        );

    \I__1812\ : InMux
    port map (
            O => \N__19175\,
            I => \N__19165\
        );

    \I__1811\ : InMux
    port map (
            O => \N__19174\,
            I => \N__19165\
        );

    \I__1810\ : InMux
    port map (
            O => \N__19173\,
            I => \N__19162\
        );

    \I__1809\ : Odrv4
    port map (
            O => \N__19170\,
            I => \nx.n10918\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__19165\,
            I => \nx.n10918\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__19162\,
            I => \nx.n10918\
        );

    \I__1806\ : InMux
    port map (
            O => \N__19155\,
            I => \N__19151\
        );

    \I__1805\ : InMux
    port map (
            O => \N__19154\,
            I => \N__19146\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__19151\,
            I => \N__19139\
        );

    \I__1803\ : InMux
    port map (
            O => \N__19150\,
            I => \N__19134\
        );

    \I__1802\ : InMux
    port map (
            O => \N__19149\,
            I => \N__19134\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__19146\,
            I => \N__19131\
        );

    \I__1800\ : InMux
    port map (
            O => \N__19145\,
            I => \N__19126\
        );

    \I__1799\ : InMux
    port map (
            O => \N__19144\,
            I => \N__19126\
        );

    \I__1798\ : InMux
    port map (
            O => \N__19143\,
            I => \N__19123\
        );

    \I__1797\ : InMux
    port map (
            O => \N__19142\,
            I => \N__19119\
        );

    \I__1796\ : Span4Mux_h
    port map (
            O => \N__19139\,
            I => \N__19108\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__19134\,
            I => \N__19108\
        );

    \I__1794\ : Span4Mux_v
    port map (
            O => \N__19131\,
            I => \N__19108\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__19126\,
            I => \N__19108\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__19123\,
            I => \N__19108\
        );

    \I__1791\ : InMux
    port map (
            O => \N__19122\,
            I => \N__19105\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__19119\,
            I => \N__19102\
        );

    \I__1789\ : Span4Mux_v
    port map (
            O => \N__19108\,
            I => \N__19099\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__19105\,
            I => \nx.start\
        );

    \I__1787\ : Odrv12
    port map (
            O => \N__19102\,
            I => \nx.start\
        );

    \I__1786\ : Odrv4
    port map (
            O => \N__19099\,
            I => \nx.start\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__19092\,
            I => \nx.n18_adj_711_cascade_\
        );

    \I__1784\ : InMux
    port map (
            O => \N__19089\,
            I => \N__19086\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__19086\,
            I => \nx.n20_adj_712\
        );

    \I__1782\ : InMux
    port map (
            O => \N__19083\,
            I => \N__19077\
        );

    \I__1781\ : InMux
    port map (
            O => \N__19082\,
            I => \N__19077\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__19077\,
            I => neo_pixel_transmitter_t0_6
        );

    \I__1779\ : InMux
    port map (
            O => \N__19074\,
            I => \N__19068\
        );

    \I__1778\ : InMux
    port map (
            O => \N__19073\,
            I => \N__19068\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__19068\,
            I => neo_pixel_transmitter_t0_14
        );

    \I__1776\ : InMux
    port map (
            O => \N__19065\,
            I => \N__19061\
        );

    \I__1775\ : InMux
    port map (
            O => \N__19064\,
            I => \N__19058\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__19061\,
            I => \N__19055\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__19058\,
            I => neo_pixel_transmitter_t0_5
        );

    \I__1772\ : Odrv4
    port map (
            O => \N__19055\,
            I => neo_pixel_transmitter_t0_5
        );

    \I__1771\ : InMux
    port map (
            O => \N__19050\,
            I => \N__19044\
        );

    \I__1770\ : InMux
    port map (
            O => \N__19049\,
            I => \N__19044\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__19044\,
            I => neo_pixel_transmitter_t0_23
        );

    \I__1768\ : CascadeMux
    port map (
            O => \N__19041\,
            I => \N__19038\
        );

    \I__1767\ : InMux
    port map (
            O => \N__19038\,
            I => \N__19032\
        );

    \I__1766\ : InMux
    port map (
            O => \N__19037\,
            I => \N__19032\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__19032\,
            I => neo_pixel_transmitter_t0_24
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__19029\,
            I => \nx.n7_adj_713_cascade_\
        );

    \I__1763\ : CEMux
    port map (
            O => \N__19026\,
            I => \N__19023\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__19023\,
            I => \nx.n13491\
        );

    \I__1761\ : CascadeMux
    port map (
            O => \N__19020\,
            I => \nx.n12933_cascade_\
        );

    \I__1760\ : InMux
    port map (
            O => \N__19017\,
            I => \N__19014\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__19014\,
            I => \nx.n12939\
        );

    \I__1758\ : InMux
    port map (
            O => \N__19011\,
            I => \nx.n10459\
        );

    \I__1757\ : InMux
    port map (
            O => \N__19008\,
            I => \bfn_1_32_0_\
        );

    \I__1756\ : InMux
    port map (
            O => \N__19005\,
            I => \N__19001\
        );

    \I__1755\ : CascadeMux
    port map (
            O => \N__19004\,
            I => \N__18998\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__19001\,
            I => \N__18995\
        );

    \I__1753\ : InMux
    port map (
            O => \N__18998\,
            I => \N__18992\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__18995\,
            I => \nx.n1203\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__18992\,
            I => \nx.n1203\
        );

    \I__1750\ : InMux
    port map (
            O => \N__18987\,
            I => \N__18984\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__18984\,
            I => \nx.n1270\
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__18981\,
            I => \nx.n1302_cascade_\
        );

    \I__1747\ : InMux
    port map (
            O => \N__18978\,
            I => \N__18975\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__18975\,
            I => \nx.n1276\
        );

    \I__1745\ : InMux
    port map (
            O => \N__18972\,
            I => \N__18968\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__18971\,
            I => \N__18964\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__18968\,
            I => \N__18961\
        );

    \I__1742\ : InMux
    port map (
            O => \N__18967\,
            I => \N__18958\
        );

    \I__1741\ : InMux
    port map (
            O => \N__18964\,
            I => \N__18955\
        );

    \I__1740\ : Odrv4
    port map (
            O => \N__18961\,
            I => \nx.n1209\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__18958\,
            I => \nx.n1209\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__18955\,
            I => \nx.n1209\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__18948\,
            I => \nx.n1206_cascade_\
        );

    \I__1736\ : InMux
    port map (
            O => \N__18945\,
            I => \N__18942\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__18942\,
            I => \nx.n1273\
        );

    \I__1734\ : CEMux
    port map (
            O => \N__18939\,
            I => \N__18936\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__18936\,
            I => \N__18933\
        );

    \I__1732\ : Span4Mux_v
    port map (
            O => \N__18933\,
            I => \N__18930\
        );

    \I__1731\ : Span4Mux_s1_h
    port map (
            O => \N__18930\,
            I => \N__18927\
        );

    \I__1730\ : Odrv4
    port map (
            O => \N__18927\,
            I => \nx.n7\
        );

    \I__1729\ : CascadeMux
    port map (
            O => \N__18924\,
            I => \nx.n1203_cascade_\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__18921\,
            I => \nx.n1208_cascade_\
        );

    \I__1727\ : InMux
    port map (
            O => \N__18918\,
            I => \bfn_1_31_0_\
        );

    \I__1726\ : InMux
    port map (
            O => \N__18915\,
            I => \nx.n10453\
        );

    \I__1725\ : InMux
    port map (
            O => \N__18912\,
            I => \nx.n10454\
        );

    \I__1724\ : InMux
    port map (
            O => \N__18909\,
            I => \nx.n10455\
        );

    \I__1723\ : InMux
    port map (
            O => \N__18906\,
            I => \nx.n10456\
        );

    \I__1722\ : InMux
    port map (
            O => \N__18903\,
            I => \nx.n10457\
        );

    \I__1721\ : InMux
    port map (
            O => \N__18900\,
            I => \nx.n10458\
        );

    \I__1720\ : InMux
    port map (
            O => \N__18897\,
            I => \N__18894\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__18894\,
            I => \N__18891\
        );

    \I__1718\ : Odrv12
    port map (
            O => \N__18891\,
            I => \nx.n3152\
        );

    \I__1717\ : InMux
    port map (
            O => \N__18888\,
            I => \nx.n10912\
        );

    \I__1716\ : InMux
    port map (
            O => \N__18885\,
            I => \nx.n10913\
        );

    \I__1715\ : InMux
    port map (
            O => \N__18882\,
            I => \nx.n10914\
        );

    \I__1714\ : CascadeMux
    port map (
            O => \N__18879\,
            I => \nx.n10_adj_619_cascade_\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__18876\,
            I => \nx.n12_adj_621_cascade_\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__18873\,
            I => \nx.n1136_cascade_\
        );

    \I__1711\ : InMux
    port map (
            O => \N__18870\,
            I => \bfn_1_28_0_\
        );

    \I__1710\ : InMux
    port map (
            O => \N__18867\,
            I => \nx.n10904\
        );

    \I__1709\ : InMux
    port map (
            O => \N__18864\,
            I => \nx.n10905\
        );

    \I__1708\ : InMux
    port map (
            O => \N__18861\,
            I => \nx.n10906\
        );

    \I__1707\ : InMux
    port map (
            O => \N__18858\,
            I => \nx.n10907\
        );

    \I__1706\ : InMux
    port map (
            O => \N__18855\,
            I => \nx.n10908\
        );

    \I__1705\ : InMux
    port map (
            O => \N__18852\,
            I => \nx.n10909\
        );

    \I__1704\ : CascadeMux
    port map (
            O => \N__18849\,
            I => \N__18846\
        );

    \I__1703\ : InMux
    port map (
            O => \N__18846\,
            I => \N__18843\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__18843\,
            I => \N__18840\
        );

    \I__1701\ : Span4Mux_v
    port map (
            O => \N__18840\,
            I => \N__18837\
        );

    \I__1700\ : Odrv4
    port map (
            O => \N__18837\,
            I => \nx.n3154\
        );

    \I__1699\ : InMux
    port map (
            O => \N__18834\,
            I => \nx.n10910\
        );

    \I__1698\ : InMux
    port map (
            O => \N__18831\,
            I => \N__18828\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__18828\,
            I => \N__18825\
        );

    \I__1696\ : Span4Mux_v
    port map (
            O => \N__18825\,
            I => \N__18822\
        );

    \I__1695\ : Odrv4
    port map (
            O => \N__18822\,
            I => \nx.n3153\
        );

    \I__1694\ : InMux
    port map (
            O => \N__18819\,
            I => \bfn_1_29_0_\
        );

    \I__1693\ : CascadeMux
    port map (
            O => \N__18816\,
            I => \N__18812\
        );

    \I__1692\ : InMux
    port map (
            O => \N__18815\,
            I => \N__18808\
        );

    \I__1691\ : InMux
    port map (
            O => \N__18812\,
            I => \N__18805\
        );

    \I__1690\ : InMux
    port map (
            O => \N__18811\,
            I => \N__18802\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__18808\,
            I => \N__18797\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__18805\,
            I => \N__18797\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__18802\,
            I => \nx.n3102\
        );

    \I__1686\ : Odrv4
    port map (
            O => \N__18797\,
            I => \nx.n3102\
        );

    \I__1685\ : InMux
    port map (
            O => \N__18792\,
            I => \N__18789\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__18789\,
            I => \N__18786\
        );

    \I__1683\ : Odrv4
    port map (
            O => \N__18786\,
            I => \nx.n3169\
        );

    \I__1682\ : InMux
    port map (
            O => \N__18783\,
            I => \bfn_1_27_0_\
        );

    \I__1681\ : InMux
    port map (
            O => \N__18780\,
            I => \nx.n10896\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__18777\,
            I => \N__18774\
        );

    \I__1679\ : InMux
    port map (
            O => \N__18774\,
            I => \N__18771\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__18771\,
            I => \N__18767\
        );

    \I__1677\ : InMux
    port map (
            O => \N__18770\,
            I => \N__18764\
        );

    \I__1676\ : Odrv4
    port map (
            O => \N__18767\,
            I => \nx.n3100\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__18764\,
            I => \nx.n3100\
        );

    \I__1674\ : InMux
    port map (
            O => \N__18759\,
            I => \N__18756\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__18756\,
            I => \N__18753\
        );

    \I__1672\ : Odrv4
    port map (
            O => \N__18753\,
            I => \nx.n3167\
        );

    \I__1671\ : InMux
    port map (
            O => \N__18750\,
            I => \nx.n10897\
        );

    \I__1670\ : InMux
    port map (
            O => \N__18747\,
            I => \nx.n10898\
        );

    \I__1669\ : InMux
    port map (
            O => \N__18744\,
            I => \nx.n10899\
        );

    \I__1668\ : InMux
    port map (
            O => \N__18741\,
            I => \nx.n10900\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__18738\,
            I => \N__18735\
        );

    \I__1666\ : InMux
    port map (
            O => \N__18735\,
            I => \N__18732\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__18732\,
            I => \N__18729\
        );

    \I__1664\ : Odrv4
    port map (
            O => \N__18729\,
            I => \nx.n3163\
        );

    \I__1663\ : InMux
    port map (
            O => \N__18726\,
            I => \nx.n10901\
        );

    \I__1662\ : InMux
    port map (
            O => \N__18723\,
            I => \nx.n10902\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__18720\,
            I => \nx.n3116_cascade_\
        );

    \I__1660\ : InMux
    port map (
            O => \N__18717\,
            I => \bfn_1_26_0_\
        );

    \I__1659\ : InMux
    port map (
            O => \N__18714\,
            I => \N__18711\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__18711\,
            I => \N__18708\
        );

    \I__1657\ : Span4Mux_h
    port map (
            O => \N__18708\,
            I => \N__18705\
        );

    \I__1656\ : Odrv4
    port map (
            O => \N__18705\,
            I => \nx.n3176\
        );

    \I__1655\ : InMux
    port map (
            O => \N__18702\,
            I => \nx.n10888\
        );

    \I__1654\ : InMux
    port map (
            O => \N__18699\,
            I => \nx.n10889\
        );

    \I__1653\ : InMux
    port map (
            O => \N__18696\,
            I => \nx.n10890\
        );

    \I__1652\ : InMux
    port map (
            O => \N__18693\,
            I => \N__18689\
        );

    \I__1651\ : InMux
    port map (
            O => \N__18692\,
            I => \N__18686\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__18689\,
            I => \N__18681\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__18686\,
            I => \N__18681\
        );

    \I__1648\ : Odrv4
    port map (
            O => \N__18681\,
            I => \nx.n3106\
        );

    \I__1647\ : InMux
    port map (
            O => \N__18678\,
            I => \N__18675\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__18675\,
            I => \N__18672\
        );

    \I__1645\ : Odrv12
    port map (
            O => \N__18672\,
            I => \nx.n3173\
        );

    \I__1644\ : InMux
    port map (
            O => \N__18669\,
            I => \nx.n10891\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__18666\,
            I => \N__18662\
        );

    \I__1642\ : CascadeMux
    port map (
            O => \N__18665\,
            I => \N__18659\
        );

    \I__1641\ : InMux
    port map (
            O => \N__18662\,
            I => \N__18656\
        );

    \I__1640\ : InMux
    port map (
            O => \N__18659\,
            I => \N__18653\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__18656\,
            I => \N__18650\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__18653\,
            I => \nx.n3105\
        );

    \I__1637\ : Odrv4
    port map (
            O => \N__18650\,
            I => \nx.n3105\
        );

    \I__1636\ : InMux
    port map (
            O => \N__18645\,
            I => \N__18642\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__18642\,
            I => \N__18639\
        );

    \I__1634\ : Odrv4
    port map (
            O => \N__18639\,
            I => \nx.n3172\
        );

    \I__1633\ : InMux
    port map (
            O => \N__18636\,
            I => \nx.n10892\
        );

    \I__1632\ : InMux
    port map (
            O => \N__18633\,
            I => \nx.n10893\
        );

    \I__1631\ : InMux
    port map (
            O => \N__18630\,
            I => \N__18627\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__18627\,
            I => \nx.n3170\
        );

    \I__1629\ : InMux
    port map (
            O => \N__18624\,
            I => \nx.n10894\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__18621\,
            I => \nx.n3100_cascade_\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__18618\,
            I => \nx.n29_adj_697_cascade_\
        );

    \I__1626\ : CascadeMux
    port map (
            O => \N__18615\,
            I => \nx.n12331_cascade_\
        );

    \I__1625\ : InMux
    port map (
            O => \N__18612\,
            I => \N__18609\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__18609\,
            I => \nx.n12335\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__18606\,
            I => \nx.n37_adj_695_cascade_\
        );

    \I__1622\ : InMux
    port map (
            O => \N__18603\,
            I => \N__18600\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__18600\,
            I => \nx.n12333\
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__18597\,
            I => \nx.n31_adj_691_cascade_\
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__18594\,
            I => \nx.n49_adj_693_cascade_\
        );

    \I__1618\ : InMux
    port map (
            O => \N__18591\,
            I => \N__18588\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__18588\,
            I => \nx.n48_adj_692\
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__18585\,
            I => \nx.n2908_cascade_\
        );

    \I__1615\ : CascadeMux
    port map (
            O => \N__18582\,
            I => \nx.n3007_cascade_\
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__18579\,
            I => \nx.n3106_cascade_\
        );

    \I__1613\ : InMux
    port map (
            O => \N__18576\,
            I => \N__18573\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__18573\,
            I => \nx.n19_adj_698\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__18570\,
            I => \nx.n3105_cascade_\
        );

    \I__1610\ : InMux
    port map (
            O => \N__18567\,
            I => \N__18564\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__18564\,
            I => \nx.n13271\
        );

    \I__1608\ : CascadeMux
    port map (
            O => \N__18561\,
            I => \nx.n12369_cascade_\
        );

    \I__1607\ : InMux
    port map (
            O => \N__18558\,
            I => \N__18552\
        );

    \I__1606\ : InMux
    port map (
            O => \N__18557\,
            I => \N__18552\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__18552\,
            I => neo_pixel_transmitter_t0_15
        );

    \I__1604\ : InMux
    port map (
            O => \N__18549\,
            I => \N__18543\
        );

    \I__1603\ : InMux
    port map (
            O => \N__18548\,
            I => \N__18543\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__18543\,
            I => neo_pixel_transmitter_t0_8
        );

    \I__1601\ : CascadeMux
    port map (
            O => \N__18540\,
            I => \nx.n9700_cascade_\
        );

    \I__1600\ : InMux
    port map (
            O => \N__18537\,
            I => \N__18534\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__18534\,
            I => \N__18531\
        );

    \I__1598\ : Odrv4
    port map (
            O => \N__18531\,
            I => \nx.n7131\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__18528\,
            I => \nx.n12117_cascade_\
        );

    \I__1596\ : CascadeMux
    port map (
            O => \N__18525\,
            I => \n7239_cascade_\
        );

    \I__1595\ : InMux
    port map (
            O => \N__18522\,
            I => \N__18515\
        );

    \I__1594\ : InMux
    port map (
            O => \N__18521\,
            I => \N__18515\
        );

    \I__1593\ : InMux
    port map (
            O => \N__18520\,
            I => \N__18512\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__18515\,
            I => \N__18509\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__18512\,
            I => \nx.n9700\
        );

    \I__1590\ : Odrv4
    port map (
            O => \N__18509\,
            I => \nx.n9700\
        );

    \I__1589\ : InMux
    port map (
            O => \N__18504\,
            I => \N__18498\
        );

    \I__1588\ : InMux
    port map (
            O => \N__18503\,
            I => \N__18498\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__18498\,
            I => \nx.n9702\
        );

    \I__1586\ : InMux
    port map (
            O => \N__18495\,
            I => \N__18492\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__18492\,
            I => \nx.n11606\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__18489\,
            I => \N__18485\
        );

    \I__1583\ : InMux
    port map (
            O => \N__18488\,
            I => \N__18482\
        );

    \I__1582\ : InMux
    port map (
            O => \N__18485\,
            I => \N__18479\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__18482\,
            I => \N__18474\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__18479\,
            I => \N__18474\
        );

    \I__1579\ : Odrv12
    port map (
            O => \N__18474\,
            I => update_color
        );

    \I__1578\ : InMux
    port map (
            O => \N__18471\,
            I => \N__18468\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__18468\,
            I => \N__18465\
        );

    \I__1576\ : Odrv4
    port map (
            O => \N__18465\,
            I => \nx.n10_adj_653\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__18462\,
            I => \nx.n7131_cascade_\
        );

    \I__1574\ : CascadeMux
    port map (
            O => \N__18459\,
            I => \nx.n13263_cascade_\
        );

    \I__1573\ : CascadeMux
    port map (
            O => \N__18456\,
            I => \nx.n7120_cascade_\
        );

    \I__1572\ : CascadeMux
    port map (
            O => \N__18453\,
            I => \nx.n13262_cascade_\
        );

    \I__1571\ : InMux
    port map (
            O => \N__18450\,
            I => \N__18447\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__18447\,
            I => \nx.n3739\
        );

    \I__1569\ : CascadeMux
    port map (
            O => \N__18444\,
            I => \nx.n3739_cascade_\
        );

    \I__1568\ : InMux
    port map (
            O => \N__18441\,
            I => \N__18435\
        );

    \I__1567\ : InMux
    port map (
            O => \N__18440\,
            I => \N__18435\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__18435\,
            I => \N__18429\
        );

    \I__1565\ : InMux
    port map (
            O => \N__18434\,
            I => \N__18424\
        );

    \I__1564\ : InMux
    port map (
            O => \N__18433\,
            I => \N__18424\
        );

    \I__1563\ : InMux
    port map (
            O => \N__18432\,
            I => \N__18421\
        );

    \I__1562\ : Odrv4
    port map (
            O => \N__18429\,
            I => \nx.n7120\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__18424\,
            I => \nx.n7120\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__18421\,
            I => \nx.n7120\
        );

    \I__1559\ : IoInMux
    port map (
            O => \N__18414\,
            I => \N__18411\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__18411\,
            I => \NEOPXL_c\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__18408\,
            I => \nx.n13325_cascade_\
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__18405\,
            I => \nx.n11535_cascade_\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__18402\,
            I => \nx.n11672_cascade_\
        );

    \I__1554\ : InMux
    port map (
            O => \N__18399\,
            I => \N__18396\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__18396\,
            I => \nx.n13326\
        );

    \I__1552\ : CEMux
    port map (
            O => \N__18393\,
            I => \N__18390\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__18390\,
            I => \N__18387\
        );

    \I__1550\ : Odrv12
    port map (
            O => \N__18387\,
            I => \nx.n11692\
        );

    \I__1549\ : SRMux
    port map (
            O => \N__18384\,
            I => \N__18381\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__18381\,
            I => \N__18378\
        );

    \I__1547\ : Span4Mux_s1_h
    port map (
            O => \N__18378\,
            I => \N__18375\
        );

    \I__1546\ : Odrv4
    port map (
            O => \N__18375\,
            I => \nx.n12204\
        );

    \I__1545\ : CascadeMux
    port map (
            O => \N__18372\,
            I => \nx.n11696_cascade_\
        );

    \I__1544\ : IoInMux
    port map (
            O => \N__18369\,
            I => \N__18366\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__18366\,
            I => \N__18363\
        );

    \I__1542\ : IoSpan4Mux
    port map (
            O => \N__18363\,
            I => \N__18360\
        );

    \I__1541\ : IoSpan4Mux
    port map (
            O => \N__18360\,
            I => \N__18357\
        );

    \I__1540\ : IoSpan4Mux
    port map (
            O => \N__18357\,
            I => \N__18354\
        );

    \I__1539\ : Odrv4
    port map (
            O => \N__18354\,
            I => \CLK_pad_gb_input\
        );

    \IN_MUX_bfv_3_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_21_0_\
        );

    \IN_MUX_bfv_3_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10429\,
            carryinitout => \bfn_3_22_0_\
        );

    \IN_MUX_bfv_3_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10436_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_3_23_0_\
        );

    \IN_MUX_bfv_3_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10442_THRU_CRY_1_THRU_CO\,
            carryinitout => \bfn_3_24_0_\
        );

    \IN_MUX_bfv_3_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10448_THRU_CRY_1_THRU_CO\,
            carryinitout => \bfn_3_25_0_\
        );

    \IN_MUX_bfv_3_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_17_0_\
        );

    \IN_MUX_bfv_3_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10486\,
            carryinitout => \bfn_3_18_0_\
        );

    \IN_MUX_bfv_3_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10494\,
            carryinitout => \bfn_3_19_0_\
        );

    \IN_MUX_bfv_3_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10502\,
            carryinitout => \bfn_3_20_0_\
        );

    \IN_MUX_bfv_2_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_31_0_\
        );

    \IN_MUX_bfv_2_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10580\,
            carryinitout => \bfn_2_32_0_\
        );

    \IN_MUX_bfv_1_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_31_0_\
        );

    \IN_MUX_bfv_1_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10460\,
            carryinitout => \bfn_1_32_0_\
        );

    \IN_MUX_bfv_2_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_29_0_\
        );

    \IN_MUX_bfv_5_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_26_0_\
        );

    \IN_MUX_bfv_6_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_28_0_\
        );

    \IN_MUX_bfv_1_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_26_0_\
        );

    \IN_MUX_bfv_1_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10895\,
            carryinitout => \bfn_1_27_0_\
        );

    \IN_MUX_bfv_1_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10903\,
            carryinitout => \bfn_1_28_0_\
        );

    \IN_MUX_bfv_1_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10911\,
            carryinitout => \bfn_1_29_0_\
        );

    \IN_MUX_bfv_3_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_26_0_\
        );

    \IN_MUX_bfv_3_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10869\,
            carryinitout => \bfn_3_27_0_\
        );

    \IN_MUX_bfv_3_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10877\,
            carryinitout => \bfn_3_28_0_\
        );

    \IN_MUX_bfv_3_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10885\,
            carryinitout => \bfn_3_29_0_\
        );

    \IN_MUX_bfv_5_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_22_0_\
        );

    \IN_MUX_bfv_5_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10844\,
            carryinitout => \bfn_5_23_0_\
        );

    \IN_MUX_bfv_5_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10852\,
            carryinitout => \bfn_5_24_0_\
        );

    \IN_MUX_bfv_5_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10860\,
            carryinitout => \bfn_5_25_0_\
        );

    \IN_MUX_bfv_6_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_21_0_\
        );

    \IN_MUX_bfv_6_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10820\,
            carryinitout => \bfn_6_22_0_\
        );

    \IN_MUX_bfv_6_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10828\,
            carryinitout => \bfn_6_23_0_\
        );

    \IN_MUX_bfv_6_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10836\,
            carryinitout => \bfn_6_24_0_\
        );

    \IN_MUX_bfv_7_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_19_0_\
        );

    \IN_MUX_bfv_7_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10797\,
            carryinitout => \bfn_7_20_0_\
        );

    \IN_MUX_bfv_7_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10805\,
            carryinitout => \bfn_7_21_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_10_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10775\,
            carryinitout => \bfn_10_18_0_\
        );

    \IN_MUX_bfv_10_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10783\,
            carryinitout => \bfn_10_19_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_12_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10754\,
            carryinitout => \bfn_12_21_0_\
        );

    \IN_MUX_bfv_12_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10762\,
            carryinitout => \bfn_12_22_0_\
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_21_0_\
        );

    \IN_MUX_bfv_14_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10734\,
            carryinitout => \bfn_14_22_0_\
        );

    \IN_MUX_bfv_14_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10742\,
            carryinitout => \bfn_14_23_0_\
        );

    \IN_MUX_bfv_15_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_23_0_\
        );

    \IN_MUX_bfv_15_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10715\,
            carryinitout => \bfn_15_24_0_\
        );

    \IN_MUX_bfv_15_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10723\,
            carryinitout => \bfn_15_25_0_\
        );

    \IN_MUX_bfv_13_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_23_0_\
        );

    \IN_MUX_bfv_13_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10697\,
            carryinitout => \bfn_13_24_0_\
        );

    \IN_MUX_bfv_13_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10705\,
            carryinitout => \bfn_13_25_0_\
        );

    \IN_MUX_bfv_11_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_23_0_\
        );

    \IN_MUX_bfv_11_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10680\,
            carryinitout => \bfn_11_24_0_\
        );

    \IN_MUX_bfv_11_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10688\,
            carryinitout => \bfn_11_25_0_\
        );

    \IN_MUX_bfv_9_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_23_0_\
        );

    \IN_MUX_bfv_9_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10664\,
            carryinitout => \bfn_9_24_0_\
        );

    \IN_MUX_bfv_9_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10672\,
            carryinitout => \bfn_9_25_0_\
        );

    \IN_MUX_bfv_7_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_25_0_\
        );

    \IN_MUX_bfv_7_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10649\,
            carryinitout => \bfn_7_26_0_\
        );

    \IN_MUX_bfv_10_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_28_0_\
        );

    \IN_MUX_bfv_10_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10622\,
            carryinitout => \bfn_10_29_0_\
        );

    \IN_MUX_bfv_7_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_30_0_\
        );

    \IN_MUX_bfv_7_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10610\,
            carryinitout => \bfn_7_31_0_\
        );

    \IN_MUX_bfv_6_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_31_0_\
        );

    \IN_MUX_bfv_6_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10599\,
            carryinitout => \bfn_6_32_0_\
        );

    \IN_MUX_bfv_3_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_31_0_\
        );

    \IN_MUX_bfv_3_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10589\,
            carryinitout => \bfn_3_32_0_\
        );

    \IN_MUX_bfv_9_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_27_0_\
        );

    \IN_MUX_bfv_9_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10635\,
            carryinitout => \bfn_9_28_0_\
        );

    \IN_MUX_bfv_4_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_27_0_\
        );

    \IN_MUX_bfv_4_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10398\,
            carryinitout => \bfn_4_28_0_\
        );

    \IN_MUX_bfv_4_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10406\,
            carryinitout => \bfn_4_29_0_\
        );

    \IN_MUX_bfv_4_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \nx.n10414\,
            carryinitout => \bfn_4_30_0_\
        );

    \IN_MUX_bfv_12_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_26_0_\
        );

    \IN_MUX_bfv_12_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n10524,
            carryinitout => \bfn_12_27_0_\
        );

    \IN_MUX_bfv_12_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n10532,
            carryinitout => \bfn_12_28_0_\
        );

    \IN_MUX_bfv_12_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n10540,
            carryinitout => \bfn_12_29_0_\
        );

    \IN_MUX_bfv_16_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_15_0_\
        );

    \IN_MUX_bfv_15_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_26_0_\
        );

    \IN_MUX_bfv_15_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n10555,
            carryinitout => \bfn_15_27_0_\
        );

    \IN_MUX_bfv_15_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n10563,
            carryinitout => \bfn_15_28_0_\
        );

    \IN_MUX_bfv_15_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n10571,
            carryinitout => \bfn_15_29_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_17_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__18369\,
            GLOBALBUFFEROUTPUT => \CLK_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \nx.one_wire_108_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19281\,
            lcout => \NEOPXL_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48384\,
            ce => \N__18393\,
            sr => \N__18384\
        );

    \nx.i9488_4_lut_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__19265\,
            in1 => \N__19388\,
            in2 => \N__19604\,
            in3 => \N__19182\,
            lcout => OPEN,
            ltout => \nx.n13325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9478_3_lut_4_lut_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19149\,
            in1 => \N__18440\,
            in2 => \N__18408\,
            in3 => \N__19511\,
            lcout => \nx.n13326\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7775_2_lut_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__18441\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19150\,
            lcout => OPEN,
            ltout => \nx.n11535_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i53_4_lut_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000110010"
        )
    port map (
            in0 => \N__19389\,
            in1 => \N__19512\,
            in2 => \N__18405\,
            in3 => \N__18521\,
            lcout => OPEN,
            ltout => \nx.n11672_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i52_4_lut_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111101111"
        )
    port map (
            in0 => \N__19603\,
            in1 => \N__19267\,
            in2 => \N__18402\,
            in3 => \N__18399\,
            lcout => \nx.n11692\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i3_4_lut_4_lut_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__18522\,
            in1 => \N__19514\,
            in2 => \N__19605\,
            in3 => \N__19266\,
            lcout => \nx.n12204\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i22_4_lut_adj_157_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011100010"
        )
    port map (
            in0 => \N__19387\,
            in1 => \N__19263\,
            in2 => \N__19181\,
            in3 => \N__19595\,
            lcout => OPEN,
            ltout => \nx.n11696_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7914_4_lut_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__19513\,
            in1 => \N__18434\,
            in2 => \N__18372\,
            in3 => \N__19145\,
            lcout => n11683,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.equal_607_i8_2_lut_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__19144\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19262\,
            lcout => \nx.n7131\,
            ltout => \nx.n7131_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9439_3_lut_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18433\,
            in2 => \N__18462\,
            in3 => \N__19174\,
            lcout => OPEN,
            ltout => \nx.n13263_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9551_4_lut_4_lut_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111001101"
        )
    port map (
            in0 => \N__19510\,
            in1 => \N__19594\,
            in2 => \N__18459\,
            in3 => \N__18450\,
            lcout => \nx.n7230\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_153_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21064\,
            in1 => \N__19017\,
            in2 => \N__21134\,
            in3 => \N__21709\,
            lcout => \nx.n7120\,
            ltout => \nx.n7120_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9469_3_lut_4_lut_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111111"
        )
    port map (
            in0 => \N__19143\,
            in1 => \N__19264\,
            in2 => \N__18456\,
            in3 => \N__19378\,
            lcout => OPEN,
            ltout => \nx.n13262_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1393_4_lut_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111110000"
        )
    port map (
            in0 => \N__20171\,
            in1 => \N__18488\,
            in2 => \N__18453\,
            in3 => \N__19480\,
            lcout => \nx.n3739\,
            ltout => \nx.n3739_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5_3_lut_adj_144_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__19586\,
            in1 => \_gnd_net_\,
            in2 => \N__18444\,
            in3 => \N__18471\,
            lcout => \nx.n7411\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \update_color_195_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25014\,
            in1 => \N__19323\,
            in2 => \N__19203\,
            in3 => \N__19305\,
            lcout => update_color,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48386\,
            ce => 'H',
            sr => \N__47115\
        );

    \nx.i7796_4_lut_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001010"
        )
    port map (
            in0 => \N__19173\,
            in1 => \N__19377\,
            in2 => \N__19596\,
            in3 => \N__18432\,
            lcout => \nx.n9702\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6476_4_lut_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__21066\,
            in1 => \N__21167\,
            in2 => \N__21135\,
            in3 => \N__21711\,
            lcout => \nx.n9700\,
            ltout => \nx.n9700_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_3_lut_4_lut_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011111111"
        )
    port map (
            in0 => \N__19282\,
            in1 => \N__19580\,
            in2 => \N__18540\,
            in3 => \N__19495\,
            lcout => OPEN,
            ltout => \nx.n12117_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_131_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010100000"
        )
    port map (
            in0 => \N__19496\,
            in1 => \N__18537\,
            in2 => \N__18528\,
            in3 => \N__18503\,
            lcout => n7239,
            ltout => \n7239_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.state_i1_LC_1_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111111110000"
        )
    port map (
            in0 => \N__20172\,
            in1 => \N__19581\,
            in2 => \N__18525\,
            in3 => \N__19500\,
            lcout => state_1_adj_726,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_adj_145_LC_1_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__18567\,
            in1 => \N__18520\,
            in2 => \N__19515\,
            in3 => \N__18495\,
            lcout => \nx.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_prev_i5_LC_1_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39795\,
            lcout => neopxl_color_prev_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7843_3_lut_LC_1_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__18504\,
            in1 => \_gnd_net_\,
            in2 => \N__19287\,
            in3 => \N__19154\,
            lcout => \nx.n11606\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.state_i0_LC_1_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__23913\,
            in1 => \N__20164\,
            in2 => \N__19668\,
            in3 => \N__19395\,
            lcout => state_0_adj_727,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48395\,
            ce => \N__19431\,
            sr => \N__19419\
        );

    \nx.i4_4_lut_4_lut_LC_1_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19479\,
            in1 => \N__19564\,
            in2 => \N__18489\,
            in3 => \N__20163\,
            lcout => \nx.n10_adj_653\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9438_2_lut_LC_1_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__19565\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19286\,
            lcout => \nx.n13271\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_128_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100100"
        )
    port map (
            in0 => \N__24213\,
            in1 => \N__19727\,
            in2 => \N__18849\,
            in3 => \N__24072\,
            lcout => OPEN,
            ltout => \nx.n12369_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_129_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__19748\,
            in1 => \N__18831\,
            in2 => \N__18561\,
            in3 => \N__24214\,
            lcout => \nx.n12371\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i9_1_lut_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18548\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \nx.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9309_3_lut_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40756\,
            in1 => \N__37434\,
            in2 => \_gnd_net_\,
            in3 => \N__23990\,
            lcout => \nx.n13156\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i15_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18558\,
            in1 => \N__21399\,
            in2 => \_gnd_net_\,
            in3 => \N__28864\,
            lcout => neo_pixel_transmitter_t0_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i16_1_lut_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18557\,
            lcout => \nx.n18_adj_623\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i8_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18549\,
            in1 => \N__28863\,
            in2 => \_gnd_net_\,
            in3 => \N__21198\,
            lcout => neo_pixel_transmitter_t0_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i5_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28862\,
            in1 => \N__20772\,
            in2 => \_gnd_net_\,
            in3 => \N__19064\,
            lcout => neo_pixel_transmitter_t0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2090_3_lut_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27400\,
            in2 => \N__23354\,
            in3 => \N__21963\,
            lcout => \nx.n3095\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1967_3_lut_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30257\,
            in2 => \N__27027\,
            in3 => \N__27003\,
            lcout => \nx.n2908\,
            ltout => \nx.n2908_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2034_3_lut_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25398\,
            in2 => \N__18585\,
            in3 => \N__31874\,
            lcout => \nx.n3007\,
            ltout => \nx.n3007_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2101_3_lut_LC_1_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__21855\,
            in1 => \_gnd_net_\,
            in2 => \N__18582\,
            in3 => \N__27401\,
            lcout => \nx.n3106\,
            ltout => \nx.n3106_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_112_LC_1_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111100"
        )
    port map (
            in0 => \N__18678\,
            in1 => \N__18576\,
            in2 => \N__18579\,
            in3 => \N__24209\,
            lcout => \nx.n12335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2147_3_lut_LC_1_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18897\,
            in2 => \N__24235\,
            in3 => \N__19694\,
            lcout => \nx.n59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2167_3_lut_LC_1_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18645\,
            in2 => \N__18665\,
            in3 => \N__24167\,
            lcout => \nx.n19_adj_698\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2100_3_lut_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23192\,
            in2 => \N__21840\,
            in3 => \N__27387\,
            lcout => \nx.n3105\,
            ltout => \nx.n3105_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i19_4_lut_adj_102_LC_1_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18770\,
            in1 => \N__20101\,
            in2 => \N__18570\,
            in3 => \N__20062\,
            lcout => \nx.n46_adj_688\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2097_3_lut_LC_1_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31733\,
            in2 => \N__22125\,
            in3 => \N__27388\,
            lcout => \nx.n3102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2095_3_lut_LC_1_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__22085\,
            in1 => \_gnd_net_\,
            in2 => \N__27436\,
            in3 => \N__22065\,
            lcout => \nx.n3100\,
            ltout => \nx.n3100_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2162_3_lut_LC_1_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__24168\,
            in1 => \_gnd_net_\,
            in2 => \N__18621\,
            in3 => \N__18759\,
            lcout => OPEN,
            ltout => \nx.n29_adj_697_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_114_LC_1_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__19823\,
            in1 => \N__18714\,
            in2 => \N__18618\,
            in3 => \N__24169\,
            lcout => OPEN,
            ltout => \nx.n12331_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_119_LC_1_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19830\,
            in1 => \N__18603\,
            in2 => \N__18615\,
            in3 => \N__18612\,
            lcout => \nx.n12349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i21_4_lut_adj_107_LC_1_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20221\,
            in1 => \N__20142\,
            in2 => \N__22281\,
            in3 => \N__19674\,
            lcout => \nx.n48_adj_692\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2158_3_lut_LC_1_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__19793\,
            in1 => \_gnd_net_\,
            in2 => \N__18738\,
            in3 => \N__24170\,
            lcout => OPEN,
            ltout => \nx.n37_adj_695_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_111_LC_1_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__24171\,
            in1 => \N__18815\,
            in2 => \N__18606\,
            in3 => \N__18792\,
            lcout => \nx.n12333\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i4_3_lut_adj_105_LC_1_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__24375\,
            in1 => \N__18811\,
            in2 => \_gnd_net_\,
            in3 => \N__19822\,
            lcout => OPEN,
            ltout => \nx.n31_adj_691_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i22_4_lut_adj_108_LC_1_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18693\,
            in1 => \N__19915\,
            in2 => \N__18597\,
            in3 => \N__23748\,
            lcout => OPEN,
            ltout => \nx.n49_adj_693_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i26_4_lut_LC_1_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19773\,
            in1 => \N__25749\,
            in2 => \N__18594\,
            in3 => \N__18591\,
            lcout => \nx.n3116\,
            ltout => \nx.n3116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2165_3_lut_LC_1_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__18630\,
            in1 => \N__19916\,
            in2 => \N__18720\,
            in3 => \_gnd_net_\,
            lcout => \nx.n23_adj_700\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_2_lut_LC_1_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24369\,
            in2 => \_gnd_net_\,
            in3 => \N__18717\,
            lcout => \nx.n3177\,
            ltout => OPEN,
            carryin => \bfn_1_26_0_\,
            carryout => \nx.n10888\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_3_lut_LC_1_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19824\,
            in3 => \N__18702\,
            lcout => \nx.n3176\,
            ltout => OPEN,
            carryin => \nx.n10888\,
            carryout => \nx.n10889\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_4_lut_LC_1_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44706\,
            in2 => \N__20003\,
            in3 => \N__18699\,
            lcout => \nx.n3175\,
            ltout => OPEN,
            carryin => \nx.n10889\,
            carryout => \nx.n10890\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_5_lut_LC_1_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20102\,
            in2 => \N__45093\,
            in3 => \N__18696\,
            lcout => \nx.n3174\,
            ltout => OPEN,
            carryin => \nx.n10890\,
            carryout => \nx.n10891\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_6_lut_LC_1_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18692\,
            in2 => \N__45094\,
            in3 => \N__18669\,
            lcout => \nx.n3173\,
            ltout => OPEN,
            carryin => \nx.n10891\,
            carryout => \nx.n10892\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_7_lut_LC_1_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44714\,
            in2 => \N__18666\,
            in3 => \N__18636\,
            lcout => \nx.n3172\,
            ltout => OPEN,
            carryin => \nx.n10892\,
            carryout => \nx.n10893\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_8_lut_LC_1_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44710\,
            in2 => \N__23777\,
            in3 => \N__18633\,
            lcout => \nx.n3171\,
            ltout => OPEN,
            carryin => \nx.n10893\,
            carryout => \nx.n10894\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_9_lut_LC_1_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44715\,
            in2 => \N__19920\,
            in3 => \N__18624\,
            lcout => \nx.n3170\,
            ltout => OPEN,
            carryin => \nx.n10894\,
            carryout => \nx.n10895\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_10_lut_LC_1_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44665\,
            in2 => \N__18816\,
            in3 => \N__18783\,
            lcout => \nx.n3169\,
            ltout => OPEN,
            carryin => \bfn_1_27_0_\,
            carryout => \nx.n10896\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_11_lut_LC_1_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45671\,
            in2 => \N__19857\,
            in3 => \N__18780\,
            lcout => \nx.n3168\,
            ltout => OPEN,
            carryin => \nx.n10896\,
            carryout => \nx.n10897\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_12_lut_LC_1_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44666\,
            in2 => \N__18777\,
            in3 => \N__18750\,
            lcout => \nx.n3167\,
            ltout => OPEN,
            carryin => \nx.n10897\,
            carryout => \nx.n10898\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_13_lut_LC_1_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45672\,
            in2 => \N__20223\,
            in3 => \N__18747\,
            lcout => \nx.n3166\,
            ltout => OPEN,
            carryin => \nx.n10898\,
            carryout => \nx.n10899\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_14_lut_LC_1_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19973\,
            in2 => \N__45755\,
            in3 => \N__18744\,
            lcout => \nx.n3165\,
            ltout => OPEN,
            carryin => \nx.n10899\,
            carryout => \nx.n10900\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_15_lut_LC_1_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19899\,
            in2 => \N__45029\,
            in3 => \N__18741\,
            lcout => \nx.n3164\,
            ltout => OPEN,
            carryin => \nx.n10900\,
            carryout => \nx.n10901\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_16_lut_LC_1_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44670\,
            in2 => \N__19797\,
            in3 => \N__18726\,
            lcout => \nx.n3163\,
            ltout => OPEN,
            carryin => \nx.n10901\,
            carryout => \nx.n10902\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_17_lut_LC_1_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45676\,
            in2 => \N__20075\,
            in3 => \N__18723\,
            lcout => \nx.n3162\,
            ltout => OPEN,
            carryin => \nx.n10902\,
            carryout => \nx.n10903\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_18_lut_LC_1_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27312\,
            in2 => \N__45758\,
            in3 => \N__18870\,
            lcout => \nx.n3161\,
            ltout => OPEN,
            carryin => \bfn_1_28_0_\,
            carryout => \nx.n10904\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_19_lut_LC_1_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25737\,
            in2 => \N__45761\,
            in3 => \N__18867\,
            lcout => \nx.n3160\,
            ltout => OPEN,
            carryin => \nx.n10904\,
            carryout => \nx.n10905\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_20_lut_LC_1_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25812\,
            in2 => \N__45759\,
            in3 => \N__18864\,
            lcout => \nx.n3159\,
            ltout => OPEN,
            carryin => \nx.n10905\,
            carryout => \nx.n10906\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_21_lut_LC_1_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25783\,
            in2 => \N__45762\,
            in3 => \N__18861\,
            lcout => \nx.n3158\,
            ltout => OPEN,
            carryin => \nx.n10906\,
            carryout => \nx.n10907\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_22_lut_LC_1_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45720\,
            in2 => \N__24288\,
            in3 => \N__18858\,
            lcout => \nx.n3157\,
            ltout => OPEN,
            carryin => \nx.n10907\,
            carryout => \nx.n10908\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_23_lut_LC_1_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24015\,
            in2 => \N__45763\,
            in3 => \N__18855\,
            lcout => \nx.n3156\,
            ltout => OPEN,
            carryin => \nx.n10908\,
            carryout => \nx.n10909\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_24_lut_LC_1_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24105\,
            in2 => \N__45760\,
            in3 => \N__18852\,
            lcout => \nx.n3155\,
            ltout => OPEN,
            carryin => \nx.n10909\,
            carryout => \nx.n10910\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_25_lut_LC_1_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19728\,
            in2 => \N__45764\,
            in3 => \N__18834\,
            lcout => \nx.n3154\,
            ltout => OPEN,
            carryin => \nx.n10910\,
            carryout => \nx.n10911\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_26_lut_LC_1_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19749\,
            in2 => \N__45625\,
            in3 => \N__18819\,
            lcout => \nx.n3153\,
            ltout => OPEN,
            carryin => \bfn_1_29_0_\,
            carryout => \nx.n10912\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_27_lut_LC_1_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19698\,
            in2 => \N__45627\,
            in3 => \N__18888\,
            lcout => \nx.n3152\,
            ltout => OPEN,
            carryin => \nx.n10912\,
            carryout => \nx.n10913\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_28_lut_LC_1_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20137\,
            in2 => \N__45626\,
            in3 => \N__18885\,
            lcout => \nx.n3151\,
            ltout => OPEN,
            carryin => \nx.n10913\,
            carryout => \nx.n10914\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2143_29_lut_LC_1_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__22277\,
            in1 => \N__45292\,
            in2 => \N__24246\,
            in3 => \N__18882\,
            lcout => \nx.n13042\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i744_3_lut_LC_1_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25707\,
            in1 => \N__26231\,
            in2 => \_gnd_net_\,
            in3 => \N__26052\,
            lcout => \nx.n1109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i3_2_lut_adj_30_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26351\,
            in3 => \N__26284\,
            lcout => OPEN,
            ltout => \nx.n10_adj_619_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5_4_lut_LC_1_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__20335\,
            in1 => \N__24460\,
            in2 => \N__18879\,
            in3 => \N__26011\,
            lcout => OPEN,
            ltout => \nx.n12_adj_621_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6_4_lut_LC_1_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25894\,
            in1 => \N__25976\,
            in2 => \N__18876\,
            in3 => \N__25931\,
            lcout => \nx.n1136\,
            ltout => \nx.n1136_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i812_3_lut_LC_1_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20346\,
            in2 => \N__18873\,
            in3 => \N__24461\,
            lcout => \nx.n1209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i806_3_lut_LC_1_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26012\,
            in2 => \N__20283\,
            in3 => \N__20424\,
            lcout => \nx.n1203\,
            ltout => \nx.n1203_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5_4_lut_adj_31_LC_1_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20513\,
            in1 => \N__22396\,
            in2 => \N__18924\,
            in3 => \N__20261\,
            lcout => \nx.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i811_3_lut_LC_1_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20336\,
            in2 => \N__20319\,
            in3 => \N__20423\,
            lcout => \nx.n1208\,
            ltout => \nx.n1208_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i3_3_lut_LC_1_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24542\,
            in2 => \N__18921\,
            in3 => \N__18967\,
            lcout => \nx.n11_adj_624\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_870_2_lut_LC_1_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24543\,
            in2 => \_gnd_net_\,
            in3 => \N__18918\,
            lcout => \nx.n1277\,
            ltout => OPEN,
            carryin => \bfn_1_31_0_\,
            carryout => \nx.n10453\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_870_3_lut_LC_1_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18971\,
            in3 => \N__18915\,
            lcout => \nx.n1276\,
            ltout => OPEN,
            carryin => \nx.n10453\,
            carryout => \nx.n10454\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_870_4_lut_LC_1_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45308\,
            in2 => \N__20448\,
            in3 => \N__18912\,
            lcout => \nx.n1275\,
            ltout => OPEN,
            carryin => \nx.n10454\,
            carryout => \nx.n10455\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_870_5_lut_LC_1_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45311\,
            in2 => \N__20385\,
            in3 => \N__18909\,
            lcout => \nx.n1274\,
            ltout => OPEN,
            carryin => \nx.n10455\,
            carryout => \nx.n10456\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_870_6_lut_LC_1_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45309\,
            in2 => \N__20477\,
            in3 => \N__18906\,
            lcout => \nx.n1273\,
            ltout => OPEN,
            carryin => \nx.n10456\,
            carryout => \nx.n10457\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_870_7_lut_LC_1_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45312\,
            in2 => \N__22403\,
            in3 => \N__18903\,
            lcout => \nx.n1272\,
            ltout => OPEN,
            carryin => \nx.n10457\,
            carryout => \nx.n10458\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_870_8_lut_LC_1_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45310\,
            in2 => \N__20517\,
            in3 => \N__18900\,
            lcout => \nx.n1271\,
            ltout => OPEN,
            carryin => \nx.n10458\,
            carryout => \nx.n10459\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_870_9_lut_LC_1_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45313\,
            in2 => \N__19004\,
            in3 => \N__19011\,
            lcout => \nx.n1270\,
            ltout => OPEN,
            carryin => \nx.n10459\,
            carryout => \nx.n10460\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_870_10_lut_LC_1_32_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__44385\,
            in1 => \N__20268\,
            in2 => \N__22378\,
            in3 => \N__19008\,
            lcout => \nx.n1301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i873_3_lut_LC_1_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19005\,
            in2 => \N__22379\,
            in3 => \N__18987\,
            lcout => \nx.n1302\,
            ltout => \nx.n1302_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_2_lut_adj_34_LC_1_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18981\,
            in3 => \N__20537\,
            lcout => \nx.n10_adj_626\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i879_3_lut_LC_1_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18978\,
            in2 => \N__22380\,
            in3 => \N__18972\,
            lcout => \nx.n1308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i809_3_lut_LC_1_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20301\,
            in2 => \N__25935\,
            in3 => \N__20427\,
            lcout => \nx.n1206\,
            ltout => \nx.n1206_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i876_3_lut_LC_1_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__22377\,
            in1 => \_gnd_net_\,
            in2 => \N__18948\,
            in3 => \N__18945\,
            lcout => \nx.n1305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.start_103_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19122\,
            in2 => \_gnd_net_\,
            in3 => \N__19527\,
            lcout => \nx.start\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48390\,
            ce => \N__18939\,
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i32_1_lut_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20594\,
            lcout => \nx.n2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i24_1_lut_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19049\,
            lcout => \nx.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i23_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19050\,
            in1 => \N__21611\,
            in2 => \_gnd_net_\,
            in3 => \N__28777\,
            lcout => neo_pixel_transmitter_t0_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i24_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28774\,
            in2 => \N__19041\,
            in3 => \N__21555\,
            lcout => neo_pixel_transmitter_t0_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i25_1_lut_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19037\,
            lcout => \nx.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_done_104_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000010001"
        )
    port map (
            in0 => \N__19142\,
            in1 => \N__19523\,
            in2 => \_gnd_net_\,
            in3 => \N__19271\,
            lcout => \nx.neo_pixel_transmitter_done\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48387\,
            ce => \N__19026\,
            sr => \_gnd_net_\
        );

    \nx.i2_2_lut_adj_149_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__21065\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21246\,
            lcout => OPEN,
            ltout => \nx.n7_adj_713_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i4_4_lut_adj_150_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__20787\,
            in1 => \N__20733\,
            in2 => \N__19029\,
            in3 => \N__19089\,
            lcout => \nx.n13491\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_2_lut_adj_151_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20786\,
            in2 => \_gnd_net_\,
            in3 => \N__20729\,
            lcout => OPEN,
            ltout => \nx.n12933_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_152_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21245\,
            in1 => \N__21228\,
            in2 => \N__19020\,
            in3 => \N__21166\,
            lcout => \nx.n12939\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i13_1_lut_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19298\,
            lcout => \nx.n21_adj_620\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i2_2_lut_adj_154_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20907\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20928\,
            lcout => \nx.n10918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i14_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19074\,
            in1 => \N__21440\,
            in2 => \_gnd_net_\,
            in3 => \N__28776\,
            lcout => neo_pixel_transmitter_t0_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i7_1_lut_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19082\,
            lcout => \nx.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7_4_lut_adj_147_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__21130\,
            in1 => \N__19209\,
            in2 => \N__19516\,
            in3 => \N__21168\,
            lcout => OPEN,
            ltout => \nx.n18_adj_711_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9_4_lut_adj_148_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__19155\,
            in1 => \N__21227\,
            in2 => \N__19092\,
            in3 => \N__21710\,
            lcout => \nx.n20_adj_712\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i6_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19083\,
            in1 => \N__28775\,
            in2 => \_gnd_net_\,
            in3 => \N__21282\,
            lcout => neo_pixel_transmitter_t0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i15_1_lut_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19073\,
            lcout => \nx.n19_adj_622\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i6_1_lut_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19065\,
            lcout => \nx.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_221_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__19329\,
            in1 => \N__39794\,
            in2 => \N__25005\,
            in3 => \N__28917\,
            lcout => n10_adj_776,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i4_1_lut_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19313\,
            lcout => \nx.n30_adj_598\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i3_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19314\,
            in1 => \N__28838\,
            in2 => \_gnd_net_\,
            in3 => \N__20876\,
            lcout => neo_pixel_transmitter_t0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__38453\,
            in1 => \N__38427\,
            in2 => \N__43125\,
            in3 => \N__43167\,
            lcout => n12_adj_774,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i12_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21021\,
            in1 => \N__19299\,
            in2 => \_gnd_net_\,
            in3 => \N__28839\,
            lcout => neo_pixel_transmitter_t0_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9545_2_lut_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__19574\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19272\,
            lcout => OPEN,
            ltout => \nx.n11487_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_146_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001110101"
        )
    port map (
            in0 => \N__20906\,
            in1 => \N__20924\,
            in2 => \N__19212\,
            in3 => \N__20849\,
            lcout => \nx.n103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_222_LC_2_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__40889\,
            in1 => \N__19188\,
            in2 => \N__37430\,
            in3 => \N__20199\,
            lcout => n9_adj_777,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_prev_i4_LC_2_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40890\,
            lcout => neopxl_color_prev_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i4155_3_lut_LC_2_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__19582\,
            in1 => \N__19504\,
            in2 => \_gnd_net_\,
            in3 => \N__19430\,
            lcout => \nx.n7392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i26_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28836\,
            in1 => \N__21491\,
            in2 => \_gnd_net_\,
            in3 => \N__19353\,
            lcout => neo_pixel_transmitter_t0_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i16_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21354\,
            in1 => \N__19341\,
            in2 => \_gnd_net_\,
            in3 => \N__28837\,
            lcout => neo_pixel_transmitter_t0_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9308_3_lut_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23991\,
            in1 => \N__40888\,
            in2 => \_gnd_net_\,
            in3 => \N__39793\,
            lcout => \nx.n13155\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.bit_ctr_1__bdd_4_lut_LC_2_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011110000"
        )
    port map (
            in0 => \N__19659\,
            in1 => \N__22851\,
            in2 => \N__23940\,
            in3 => \N__19616\,
            lcout => OPEN,
            ltout => \nx.n13456_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.n13456_bdd_4_lut_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__19617\,
            in1 => \N__19410\,
            in2 => \N__19404\,
            in3 => \N__19401\,
            lcout => \nx.n13459\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_2_lut_adj_156_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20905\,
            in2 => \_gnd_net_\,
            in3 => \N__20848\,
            lcout => \nx.n4_adj_642\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i27_1_lut_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19352\,
            lcout => \nx.n7_adj_597\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i17_1_lut_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19340\,
            lcout => \nx.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9470_3_lut_LC_2_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__20031\,
            in1 => \N__23889\,
            in2 => \_gnd_net_\,
            in3 => \N__19626\,
            lcout => \nx.color_bit_N_571_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9311_3_lut_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28916\,
            in1 => \N__23989\,
            in2 => \_gnd_net_\,
            in3 => \N__38445\,
            lcout => \nx.n13158\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_i12_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101100101010"
        )
    port map (
            in0 => \N__38446\,
            in1 => \N__50079\,
            in2 => \N__49851\,
            in3 => \N__49589\,
            lcout => neopxl_color_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48407\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_130_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19653\,
            in1 => \N__20232\,
            in2 => \N__19647\,
            in3 => \N__19638\,
            lcout => \nx.n10947\,
            ltout => \nx.n10947_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_2_lut_adj_58_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19620\,
            in3 => \N__23888\,
            lcout => \nx.n10975\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2028_3_lut_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30411\,
            in2 => \N__25287\,
            in3 => \N__31852\,
            lcout => \nx.n3001\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2080_3_lut_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27421\,
            in2 => \N__23460\,
            in3 => \N__22308\,
            lcout => \nx.n3085\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2035_3_lut_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29776\,
            in2 => \N__25197\,
            in3 => \N__31851\,
            lcout => \nx.n3008\,
            ltout => \nx.n3008_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i19_4_lut_adj_96_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23347\,
            in1 => \N__22030\,
            in2 => \N__19608\,
            in3 => \N__22084\,
            lcout => \nx.n45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2026_3_lut_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29715\,
            in2 => \N__25578\,
            in3 => \N__31853\,
            lcout => \nx.n2999\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2091_3_lut_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23319\,
            in2 => \N__21981\,
            in3 => \N__27422\,
            lcout => \nx.n3096\,
            ltout => \nx.n3096_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i20_4_lut_adj_109_LC_2_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19966\,
            in1 => \N__19898\,
            in2 => \N__19776\,
            in3 => \N__20004\,
            lcout => \nx.n47_adj_694\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2096_3_lut_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22107\,
            in2 => \N__23534\,
            in3 => \N__27415\,
            lcout => \nx.n3101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i23_4_lut_adj_101_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21869\,
            in1 => \N__23599\,
            in2 => \N__19764\,
            in3 => \N__23427\,
            lcout => OPEN,
            ltout => \nx.n49_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i25_4_lut_LC_2_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23502\,
            in1 => \N__23547\,
            in2 => \N__19755\,
            in3 => \N__22986\,
            lcout => \nx.n3017\,
            ltout => \nx.n3017_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2082_3_lut_LC_2_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23576\,
            in2 => \N__19752\,
            in3 => \N__22155\,
            lcout => \nx.n3087\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2081_3_lut_LC_2_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27420\,
            in2 => \N__23283\,
            in3 => \N__22140\,
            lcout => \nx.n3086\,
            ltout => \nx.n3086_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_adj_103_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19846\,
            in1 => \N__19717\,
            in2 => \N__19701\,
            in3 => \N__19690\,
            lcout => \nx.n42_adj_689\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2093_3_lut_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22031\,
            in2 => \N__22011\,
            in3 => \N__27419\,
            lcout => \nx.n3098\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2098_3_lut_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23600\,
            in2 => \N__27451\,
            in3 => \N__21813\,
            lcout => \nx.n3103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2092_3_lut_LC_2_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23159\,
            in2 => \N__21996\,
            in3 => \N__27399\,
            lcout => \nx.n3097\,
            ltout => \nx.n3097_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2159_3_lut_LC_2_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19881\,
            in2 => \N__19872\,
            in3 => \N__24172\,
            lcout => OPEN,
            ltout => \nx.n35_adj_699_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_113_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__24173\,
            in1 => \N__19869\,
            in2 => \N__19860\,
            in3 => \N__19850\,
            lcout => \nx.n12337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2104_3_lut_LC_2_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__21927\,
            in1 => \_gnd_net_\,
            in2 => \N__27438\,
            in3 => \N__26175\,
            lcout => \nx.n3109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_120_LC_2_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__20027\,
            in1 => \N__23878\,
            in2 => \N__19929\,
            in3 => \N__19803\,
            lcout => \nx.n12353\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2099_3_lut_LC_2_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23246\,
            in2 => \N__27437\,
            in3 => \N__21822\,
            lcout => \nx.n3104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2102_3_lut_LC_2_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21905\,
            in2 => \N__21888\,
            in3 => \N__27389\,
            lcout => \nx.n3107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2103_3_lut_LC_2_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__23493\,
            in1 => \_gnd_net_\,
            in2 => \N__27439\,
            in3 => \N__21915\,
            lcout => \nx.n3108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_115_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111100"
        )
    port map (
            in0 => \N__20118\,
            in1 => \N__20112\,
            in2 => \N__20106\,
            in3 => \N__24174\,
            lcout => OPEN,
            ltout => \nx.n12327_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_117_LC_2_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__24176\,
            in1 => \N__20085\,
            in2 => \N__20079\,
            in3 => \N__20076\,
            lcout => \nx.n12339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2161_3_lut_LC_2_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20222\,
            in2 => \N__20046\,
            in3 => \N__24177\,
            lcout => \nx.n31_adj_702\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2172_3_lut_LC_2_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__24370\,
            in1 => \N__20037\,
            in2 => \N__24208\,
            in3 => \_gnd_net_\,
            lcout => \nx.n3209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2166_3_lut_LC_2_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20016\,
            in2 => \N__23778\,
            in3 => \N__24175\,
            lcout => \nx.n21_adj_701\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2170_3_lut_LC_2_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20010\,
            in2 => \N__24207\,
            in3 => \N__20002\,
            lcout => OPEN,
            ltout => \nx.n13_adj_696_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_116_LC_2_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__19980\,
            in1 => \N__19974\,
            in2 => \N__19953\,
            in3 => \N__24181\,
            lcout => OPEN,
            ltout => \nx.n12325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_118_LC_2_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19950\,
            in1 => \N__19944\,
            in2 => \N__19938\,
            in3 => \N__19935\,
            lcout => \nx.n12347\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2086_3_lut_LC_2_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22173\,
            in2 => \N__23847\,
            in3 => \N__27440\,
            lcout => \nx.n3091\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2146_3_lut_LC_2_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20138\,
            in1 => \N__20241\,
            in2 => \_gnd_net_\,
            in3 => \N__24234\,
            lcout => \nx.n61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2094_3_lut_LC_2_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23390\,
            in2 => \N__22050\,
            in3 => \N__27441\,
            lcout => \nx.n3099\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_prev_i7_LC_2_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37423\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => neopxl_color_prev_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48419\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i26_4_lut_adj_141_LC_2_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25953\,
            in1 => \N__24501\,
            in2 => \N__26406\,
            in3 => \N__22257\,
            lcout => \nx.n54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i21_4_lut_adj_142_LC_2_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34977\,
            in1 => \N__28069\,
            in2 => \N__24462\,
            in3 => \N__28533\,
            lcout => \nx.n49_adj_710\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_adj_140_LC_2_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__23887\,
            in1 => \N__24374\,
            in2 => \N__39846\,
            in3 => \N__32682\,
            lcout => OPEN,
            ltout => \nx.n43_adj_709_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i27_4_lut_LC_2_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20187\,
            in1 => \N__26091\,
            in2 => \N__20181\,
            in3 => \N__20178\,
            lcout => \state_3_N_377_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2079_3_lut_LC_2_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22293\,
            in2 => \N__23127\,
            in3 => \N__27459\,
            lcout => \nx.n3084\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_803_2_lut_LC_2_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24456\,
            in2 => \_gnd_net_\,
            in3 => \N__20340\,
            lcout => \nx.n1177\,
            ltout => OPEN,
            carryin => \bfn_2_29_0_\,
            carryout => \nx.n10461\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_803_3_lut_LC_2_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20337\,
            in3 => \N__20307\,
            lcout => \nx.n1176\,
            ltout => OPEN,
            carryin => \nx.n10461\,
            carryout => \nx.n10462\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_803_4_lut_LC_2_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45280\,
            in2 => \N__26352\,
            in3 => \N__20304\,
            lcout => \nx.n1175\,
            ltout => OPEN,
            carryin => \nx.n10462\,
            carryout => \nx.n10463\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_803_5_lut_LC_2_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45284\,
            in2 => \N__25930\,
            in3 => \N__20292\,
            lcout => \nx.n1174\,
            ltout => OPEN,
            carryin => \nx.n10463\,
            carryout => \nx.n10464\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_803_6_lut_LC_2_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45281\,
            in2 => \N__26292\,
            in3 => \N__20289\,
            lcout => \nx.n1173\,
            ltout => OPEN,
            carryin => \nx.n10464\,
            carryout => \nx.n10465\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_803_7_lut_LC_2_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45285\,
            in2 => \N__25896\,
            in3 => \N__20286\,
            lcout => \nx.n1172\,
            ltout => OPEN,
            carryin => \nx.n10465\,
            carryout => \nx.n10466\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_803_8_lut_LC_2_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45282\,
            in2 => \N__26016\,
            in3 => \N__20274\,
            lcout => \nx.n1171\,
            ltout => OPEN,
            carryin => \nx.n10466\,
            carryout => \nx.n10467\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_803_9_lut_LC_2_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__45283\,
            in1 => \N__20419\,
            in2 => \N__25977\,
            in3 => \N__20271\,
            lcout => \nx.n1202\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i808_3_lut_LC_2_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26291\,
            in2 => \N__20250\,
            in3 => \N__20412\,
            lcout => \nx.n1205\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i807_3_lut_LC_2_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25895\,
            in2 => \N__20425\,
            in3 => \N__20523\,
            lcout => \nx.n1204\,
            ltout => \nx.n1204_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i874_3_lut_LC_2_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20502\,
            in2 => \N__20496\,
            in3 => \N__22367\,
            lcout => \nx.n1303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7_4_lut_adj_32_LC_2_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20381\,
            in1 => \N__20493\,
            in2 => \N__20487\,
            in3 => \N__20478\,
            lcout => \nx.n1235\,
            ltout => \nx.n1235_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i878_3_lut_LC_2_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20457\,
            in2 => \N__20451\,
            in3 => \N__20447\,
            lcout => \nx.n1307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i810_3_lut_LC_2_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20433\,
            in2 => \N__20426\,
            in3 => \N__26347\,
            lcout => \nx.n1207\,
            ltout => \nx.n1207_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i877_3_lut_LC_2_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__20370\,
            in1 => \_gnd_net_\,
            in2 => \N__20364\,
            in3 => \N__22366\,
            lcout => \nx.n1306\,
            ltout => \nx.n1306_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7_4_lut_adj_35_LC_2_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22240\,
            in1 => \N__24733\,
            in2 => \N__20361\,
            in3 => \N__20358\,
            lcout => \nx.n16_adj_627\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_2_lut_LC_2_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32717\,
            in2 => \_gnd_net_\,
            in3 => \N__20349\,
            lcout => \nx.n1377\,
            ltout => OPEN,
            carryin => \bfn_2_31_0_\,
            carryout => \nx.n10573\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_3_lut_LC_2_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22203\,
            in3 => \N__20565\,
            lcout => \nx.n1376\,
            ltout => OPEN,
            carryin => \nx.n10573\,
            carryout => \nx.n10574\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_4_lut_LC_2_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45298\,
            in2 => \N__24734\,
            in3 => \N__20562\,
            lcout => \nx.n1375\,
            ltout => OPEN,
            carryin => \nx.n10574\,
            carryout => \nx.n10575\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_5_lut_LC_2_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22241\,
            in2 => \N__45628\,
            in3 => \N__20559\,
            lcout => \nx.n1374\,
            ltout => OPEN,
            carryin => \nx.n10575\,
            carryout => \nx.n10576\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_6_lut_LC_2_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45302\,
            in2 => \N__24683\,
            in3 => \N__20556\,
            lcout => \nx.n1373\,
            ltout => OPEN,
            carryin => \nx.n10576\,
            carryout => \nx.n10577\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_7_lut_LC_2_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45303\,
            in2 => \N__24631\,
            in3 => \N__20553\,
            lcout => \nx.n1372\,
            ltout => OPEN,
            carryin => \nx.n10577\,
            carryout => \nx.n10578\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_8_lut_LC_2_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24652\,
            in2 => \N__45629\,
            in3 => \N__20550\,
            lcout => \nx.n1371\,
            ltout => OPEN,
            carryin => \nx.n10578\,
            carryout => \nx.n10579\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_9_lut_LC_2_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45307\,
            in2 => \N__22517\,
            in3 => \N__20547\,
            lcout => \nx.n1370\,
            ltout => OPEN,
            carryin => \nx.n10579\,
            carryout => \nx.n10580\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_10_lut_LC_2_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44833\,
            in2 => \N__20625\,
            in3 => \N__20544\,
            lcout => \nx.n1369\,
            ltout => OPEN,
            carryin => \bfn_2_32_0_\,
            carryout => \nx.n10581\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_937_11_lut_LC_2_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__44834\,
            in1 => \N__24589\,
            in2 => \N__20541\,
            in3 => \N__20526\,
            lcout => \nx.n1400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i940_3_lut_LC_2_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20624\,
            in2 => \N__20613\,
            in3 => \N__24588\,
            lcout => \nx.n1401\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i4_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20583\,
            in1 => \N__20817\,
            in2 => \_gnd_net_\,
            in3 => \N__28858\,
            lcout => neo_pixel_transmitter_t0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i1_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28857\,
            in1 => \N__20951\,
            in2 => \_gnd_net_\,
            in3 => \N__20604\,
            lcout => neo_pixel_transmitter_t0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i2_1_lut_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20603\,
            lcout => \nx.n32_adj_651\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i31_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28841\,
            in1 => \N__21765\,
            in2 => \_gnd_net_\,
            in3 => \N__20595\,
            lcout => neo_pixel_transmitter_t0_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i10_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28840\,
            in1 => \N__21096\,
            in2 => \_gnd_net_\,
            in3 => \N__22610\,
            lcout => neo_pixel_transmitter_t0_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i5_1_lut_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20582\,
            lcout => \nx.n29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i0_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28666\,
            in2 => \_gnd_net_\,
            in3 => \N__20571\,
            lcout => timer_0,
            ltout => OPEN,
            carryin => \bfn_3_17_0_\,
            carryout => \nx.n10479\,
            clk => \N__48385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i1_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20947\,
            in2 => \_gnd_net_\,
            in3 => \N__20568\,
            lcout => timer_1,
            ltout => OPEN,
            carryin => \nx.n10479\,
            carryout => \nx.n10480\,
            clk => \N__48385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i2_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22693\,
            in2 => \_gnd_net_\,
            in3 => \N__20655\,
            lcout => timer_2,
            ltout => OPEN,
            carryin => \nx.n10480\,
            carryout => \nx.n10481\,
            clk => \N__48385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i3_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20869\,
            in2 => \_gnd_net_\,
            in3 => \N__20652\,
            lcout => timer_3,
            ltout => OPEN,
            carryin => \nx.n10481\,
            carryout => \nx.n10482\,
            clk => \N__48385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i4_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20803\,
            in2 => \_gnd_net_\,
            in3 => \N__20649\,
            lcout => timer_4,
            ltout => OPEN,
            carryin => \nx.n10482\,
            carryout => \nx.n10483\,
            clk => \N__48385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i5_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20761\,
            in2 => \_gnd_net_\,
            in3 => \N__20646\,
            lcout => timer_5,
            ltout => OPEN,
            carryin => \nx.n10483\,
            carryout => \nx.n10484\,
            clk => \N__48385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i6_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21277\,
            in2 => \_gnd_net_\,
            in3 => \N__20643\,
            lcout => timer_6,
            ltout => OPEN,
            carryin => \nx.n10484\,
            carryout => \nx.n10485\,
            clk => \N__48385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i7_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22870\,
            in2 => \_gnd_net_\,
            in3 => \N__20640\,
            lcout => timer_7,
            ltout => OPEN,
            carryin => \nx.n10485\,
            carryout => \nx.n10486\,
            clk => \N__48385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i8_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21187\,
            in2 => \_gnd_net_\,
            in3 => \N__20637\,
            lcout => timer_8,
            ltout => OPEN,
            carryin => \bfn_3_18_0_\,
            carryout => \nx.n10487\,
            clk => \N__48393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i9_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22630\,
            in2 => \_gnd_net_\,
            in3 => \N__20634\,
            lcout => timer_9,
            ltout => OPEN,
            carryin => \nx.n10487\,
            carryout => \nx.n10488\,
            clk => \N__48393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i10_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21082\,
            in2 => \_gnd_net_\,
            in3 => \N__20631\,
            lcout => timer_10,
            ltout => OPEN,
            carryin => \nx.n10488\,
            carryout => \nx.n10489\,
            clk => \N__48393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i11_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22552\,
            in2 => \_gnd_net_\,
            in3 => \N__20628\,
            lcout => timer_11,
            ltout => OPEN,
            carryin => \nx.n10489\,
            carryout => \nx.n10490\,
            clk => \N__48393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i12_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21016\,
            in2 => \_gnd_net_\,
            in3 => \N__20682\,
            lcout => timer_12,
            ltout => OPEN,
            carryin => \nx.n10490\,
            carryout => \nx.n10491\,
            clk => \N__48393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i13_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22942\,
            in2 => \_gnd_net_\,
            in3 => \N__20679\,
            lcout => timer_13,
            ltout => OPEN,
            carryin => \nx.n10491\,
            carryout => \nx.n10492\,
            clk => \N__48393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i14_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21439\,
            in2 => \_gnd_net_\,
            in3 => \N__20676\,
            lcout => timer_14,
            ltout => OPEN,
            carryin => \nx.n10492\,
            carryout => \nx.n10493\,
            clk => \N__48393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i15_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21388\,
            in2 => \_gnd_net_\,
            in3 => \N__20673\,
            lcout => timer_15,
            ltout => OPEN,
            carryin => \nx.n10493\,
            carryout => \nx.n10494\,
            clk => \N__48393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i16_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21337\,
            in2 => \_gnd_net_\,
            in3 => \N__20670\,
            lcout => timer_16,
            ltout => OPEN,
            carryin => \bfn_3_19_0_\,
            carryout => \nx.n10495\,
            clk => \N__48398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i17_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22729\,
            in2 => \_gnd_net_\,
            in3 => \N__20667\,
            lcout => timer_17,
            ltout => OPEN,
            carryin => \nx.n10495\,
            carryout => \nx.n10496\,
            clk => \N__48398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i18_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22783\,
            in2 => \_gnd_net_\,
            in3 => \N__20664\,
            lcout => timer_18,
            ltout => OPEN,
            carryin => \nx.n10496\,
            carryout => \nx.n10497\,
            clk => \N__48398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i19_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25120\,
            in2 => \_gnd_net_\,
            in3 => \N__20661\,
            lcout => timer_19,
            ltout => OPEN,
            carryin => \nx.n10497\,
            carryout => \nx.n10498\,
            clk => \N__48398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i20_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25168\,
            in2 => \_gnd_net_\,
            in3 => \N__20658\,
            lcout => timer_20,
            ltout => OPEN,
            carryin => \nx.n10498\,
            carryout => \nx.n10499\,
            clk => \N__48398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i21_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22969\,
            in2 => \_gnd_net_\,
            in3 => \N__20709\,
            lcout => timer_21,
            ltout => OPEN,
            carryin => \nx.n10499\,
            carryout => \nx.n10500\,
            clk => \N__48398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i22_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24868\,
            in2 => \_gnd_net_\,
            in3 => \N__20706\,
            lcout => timer_22,
            ltout => OPEN,
            carryin => \nx.n10500\,
            carryout => \nx.n10501\,
            clk => \N__48398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i23_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21598\,
            in2 => \_gnd_net_\,
            in3 => \N__20703\,
            lcout => timer_23,
            ltout => OPEN,
            carryin => \nx.n10501\,
            carryout => \nx.n10502\,
            clk => \N__48398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i24_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21547\,
            in2 => \_gnd_net_\,
            in3 => \N__20700\,
            lcout => timer_24,
            ltout => OPEN,
            carryin => \bfn_3_20_0_\,
            carryout => \nx.n10503\,
            clk => \N__48403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i25_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22807\,
            in2 => \_gnd_net_\,
            in3 => \N__20697\,
            lcout => timer_25,
            ltout => OPEN,
            carryin => \nx.n10503\,
            carryout => \nx.n10504\,
            clk => \N__48403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i26_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21481\,
            in2 => \_gnd_net_\,
            in3 => \N__20694\,
            lcout => timer_26,
            ltout => OPEN,
            carryin => \nx.n10504\,
            carryout => \nx.n10505\,
            clk => \N__48403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i27_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21670\,
            in2 => \_gnd_net_\,
            in3 => \N__20691\,
            lcout => timer_27,
            ltout => OPEN,
            carryin => \nx.n10505\,
            carryout => \nx.n10506\,
            clk => \N__48403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i28_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23029\,
            in2 => \_gnd_net_\,
            in3 => \N__20688\,
            lcout => timer_28,
            ltout => OPEN,
            carryin => \nx.n10506\,
            carryout => \nx.n10507\,
            clk => \N__48403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i29_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22654\,
            in2 => \_gnd_net_\,
            in3 => \N__20685\,
            lcout => timer_29,
            ltout => OPEN,
            carryin => \nx.n10507\,
            carryout => \nx.n10508\,
            clk => \N__48403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i30_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22444\,
            in2 => \_gnd_net_\,
            in3 => \N__20967\,
            lcout => timer_30,
            ltout => OPEN,
            carryin => \nx.n10508\,
            carryout => \nx.n10509\,
            clk => \N__48403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.timer_1102__i31_LC_3_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21757\,
            in2 => \_gnd_net_\,
            in3 => \N__20964\,
            lcout => timer_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48403\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_2_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28635\,
            in2 => \N__28677\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_21_0_\,
            carryout => \nx.n10422\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_3_lut_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__20850\,
            in1 => \N__20961\,
            in2 => \N__20952\,
            in3 => \N__20910\,
            lcout => \nx.n11533\,
            ltout => OPEN,
            carryin => \nx.n10422\,
            carryout => \nx.n10423\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_4_lut_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22764\,
            in2 => \N__22698\,
            in3 => \N__20886\,
            lcout => \nx.one_wire_N_528_2\,
            ltout => OPEN,
            carryin => \nx.n10423\,
            carryout => \nx.n10424\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_5_lut_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20883\,
            in2 => \N__20877\,
            in3 => \N__20829\,
            lcout => \nx.one_wire_N_528_3\,
            ltout => OPEN,
            carryin => \nx.n10424\,
            carryout => \nx.n10425\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_6_lut_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20826\,
            in2 => \N__20816\,
            in3 => \N__20775\,
            lcout => \nx.one_wire_N_528_4\,
            ltout => OPEN,
            carryin => \nx.n10425\,
            carryout => \nx.n10426\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_7_lut_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20771\,
            in2 => \N__20742\,
            in3 => \N__20712\,
            lcout => \nx.one_wire_N_528_5\,
            ltout => OPEN,
            carryin => \nx.n10426\,
            carryout => \nx.n10427\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_8_lut_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21281\,
            in2 => \N__21258\,
            in3 => \N__21231\,
            lcout => \nx.one_wire_N_528_6\,
            ltout => OPEN,
            carryin => \nx.n10427\,
            carryout => \nx.n10428\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_9_lut_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23199\,
            in2 => \N__22881\,
            in3 => \N__21210\,
            lcout => \nx.one_wire_N_528_7\,
            ltout => OPEN,
            carryin => \nx.n10428\,
            carryout => \nx.n10429\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_10_lut_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21207\,
            in2 => \N__21197\,
            in3 => \N__21138\,
            lcout => \nx.one_wire_N_528_8\,
            ltout => OPEN,
            carryin => \bfn_3_22_0_\,
            carryout => \nx.n10430\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_11_lut_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25074\,
            in2 => \N__22635\,
            in3 => \N__21099\,
            lcout => \nx.one_wire_N_528_9\,
            ltout => OPEN,
            carryin => \nx.n10430\,
            carryout => \nx.n10431\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_12_lut_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22596\,
            in2 => \N__21095\,
            in3 => \N__21033\,
            lcout => \nx.one_wire_N_528_10\,
            ltout => OPEN,
            carryin => \nx.n10431\,
            carryout => \nx.n10432\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_13_lut_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22911\,
            in2 => \N__22557\,
            in3 => \N__21030\,
            lcout => \nx.one_wire_N_528_11\,
            ltout => OPEN,
            carryin => \nx.n10432\,
            carryout => \nx.n10433\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_14_lut_LC_3_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21027\,
            in1 => \N__21020\,
            in2 => \N__20997\,
            in3 => \N__20979\,
            lcout => \nx.n12945\,
            ltout => OPEN,
            carryin => \nx.n10433\,
            carryout => \nx.n10434\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_15_lut_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__20976\,
            in1 => \N__22890\,
            in2 => \N__22950\,
            in3 => \N__20970\,
            lcout => \nx.n12947\,
            ltout => OPEN,
            carryin => \nx.n10434\,
            carryout => \nx.n10435\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_16_lut_LC_3_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21462\,
            in1 => \N__21456\,
            in2 => \N__21447\,
            in3 => \N__21420\,
            lcout => \nx.n12949\,
            ltout => OPEN,
            carryin => \nx.n10435\,
            carryout => \nx.n10436\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_16_THRU_CRY_0_LC_3_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45757\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \nx.n10436\,
            carryout => \nx.n10436_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_17_lut_LC_3_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21417\,
            in1 => \N__21411\,
            in2 => \N__21398\,
            in3 => \N__21369\,
            lcout => \nx.n12951\,
            ltout => OPEN,
            carryin => \bfn_3_23_0_\,
            carryout => \nx.n10437\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_18_lut_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21366\,
            in1 => \N__21360\,
            in2 => \N__21350\,
            in3 => \N__21321\,
            lcout => \nx.n12953\,
            ltout => OPEN,
            carryin => \nx.n10437\,
            carryout => \nx.n10438\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_19_lut_LC_3_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21318\,
            in1 => \N__22737\,
            in2 => \N__22752\,
            in3 => \N__21312\,
            lcout => \nx.n12955\,
            ltout => OPEN,
            carryin => \nx.n10438\,
            carryout => \nx.n10439\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_20_lut_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21309\,
            in1 => \N__23046\,
            in2 => \N__22788\,
            in3 => \N__21303\,
            lcout => \nx.n12957\,
            ltout => OPEN,
            carryin => \nx.n10439\,
            carryout => \nx.n10440\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_21_lut_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21300\,
            in1 => \N__25124\,
            in2 => \N__25047\,
            in3 => \N__21294\,
            lcout => \nx.n12959\,
            ltout => OPEN,
            carryin => \nx.n10440\,
            carryout => \nx.n10441\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_22_lut_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21291\,
            in1 => \N__24990\,
            in2 => \N__25179\,
            in3 => \N__21285\,
            lcout => \nx.n12961\,
            ltout => OPEN,
            carryin => \nx.n10441\,
            carryout => \nx.n10442\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_22_THRU_CRY_0_LC_3_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45666\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \nx.n10442\,
            carryout => \nx.n10442_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_22_THRU_CRY_1_LC_3_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__45754\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \nx.n10442_THRU_CRY_0_THRU_CO\,
            carryout => \nx.n10442_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_23_lut_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21651\,
            in1 => \N__22827\,
            in2 => \N__22974\,
            in3 => \N__21645\,
            lcout => \nx.n12963\,
            ltout => OPEN,
            carryin => \bfn_3_24_0_\,
            carryout => \nx.n10443\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_24_lut_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21642\,
            in1 => \N__24872\,
            in2 => \N__29262\,
            in3 => \N__21636\,
            lcout => \nx.n12965\,
            ltout => OPEN,
            carryin => \nx.n10443\,
            carryout => \nx.n10444\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_25_lut_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21633\,
            in1 => \N__21627\,
            in2 => \N__21612\,
            in3 => \N__21579\,
            lcout => \nx.n12967\,
            ltout => OPEN,
            carryin => \nx.n10444\,
            carryout => \nx.n10445\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_26_lut_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21576\,
            in1 => \N__21567\,
            in2 => \N__21554\,
            in3 => \N__21528\,
            lcout => \nx.n12969\,
            ltout => OPEN,
            carryin => \nx.n10445\,
            carryout => \nx.n10446\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_27_lut_LC_3_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21525\,
            in1 => \N__23067\,
            in2 => \N__22815\,
            in3 => \N__21516\,
            lcout => \nx.n12971\,
            ltout => OPEN,
            carryin => \nx.n10446\,
            carryout => \nx.n10447\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_28_lut_LC_3_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21513\,
            in1 => \N__21507\,
            in2 => \N__21492\,
            in3 => \N__21465\,
            lcout => \nx.n12973\,
            ltout => OPEN,
            carryin => \nx.n10447\,
            carryout => \nx.n10448\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_28_THRU_CRY_0_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45635\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \nx.n10448\,
            carryout => \nx.n10448_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_28_THRU_CRY_1_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__45750\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \nx.n10448_THRU_CRY_0_THRU_CO\,
            carryout => \nx.n10448_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_29_lut_LC_3_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21801\,
            in1 => \N__21933\,
            in2 => \N__21675\,
            in3 => \N__21795\,
            lcout => \nx.n12975\,
            ltout => OPEN,
            carryin => \bfn_3_25_0_\,
            carryout => \nx.n10449\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_30_lut_LC_3_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21792\,
            in1 => \N__23034\,
            in2 => \N__23097\,
            in3 => \N__21786\,
            lcout => \nx.n12977\,
            ltout => OPEN,
            carryin => \nx.n10449\,
            carryout => \nx.n10450\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_31_lut_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21783\,
            in1 => \N__22662\,
            in2 => \N__22575\,
            in3 => \N__21777\,
            lcout => \nx.n12979\,
            ltout => OPEN,
            carryin => \nx.n10450\,
            carryout => \nx.n10451\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_32_lut_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__21774\,
            in1 => \N__22454\,
            in2 => \N__22473\,
            in3 => \N__21768\,
            lcout => \nx.n12981\,
            ltout => OPEN,
            carryin => \nx.n10451\,
            carryout => \nx.n10452\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_add_2_33_lut_LC_3_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__21764\,
            in1 => \N__21738\,
            in2 => \N__21723\,
            in3 => \N__21714\,
            lcout => \nx.n7181\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i27_LC_3_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21942\,
            in1 => \N__21674\,
            in2 => \_gnd_net_\,
            in3 => \N__28876\,
            lcout => neo_pixel_transmitter_t0_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48416\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i28_1_lut_LC_3_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21941\,
            lcout => \nx.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_2_lut_LC_3_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26162\,
            in2 => \_gnd_net_\,
            in3 => \N__21918\,
            lcout => \nx.n3077\,
            ltout => OPEN,
            carryin => \bfn_3_26_0_\,
            carryout => \nx.n10862\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_3_lut_LC_3_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23485\,
            in3 => \N__21909\,
            lcout => \nx.n3076\,
            ltout => OPEN,
            carryin => \nx.n10862\,
            carryout => \nx.n10863\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_4_lut_LC_3_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45632\,
            in2 => \N__21906\,
            in3 => \N__21879\,
            lcout => \nx.n3075\,
            ltout => OPEN,
            carryin => \nx.n10863\,
            carryout => \nx.n10864\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_5_lut_LC_3_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45090\,
            in2 => \N__21876\,
            in3 => \N__21843\,
            lcout => \nx.n3074\,
            ltout => OPEN,
            carryin => \nx.n10864\,
            carryout => \nx.n10865\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_6_lut_LC_3_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45633\,
            in2 => \N__23193\,
            in3 => \N__21825\,
            lcout => \nx.n3073\,
            ltout => OPEN,
            carryin => \nx.n10865\,
            carryout => \nx.n10866\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_7_lut_LC_3_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45091\,
            in2 => \N__23247\,
            in3 => \N__21816\,
            lcout => \nx.n3072\,
            ltout => OPEN,
            carryin => \nx.n10866\,
            carryout => \nx.n10867\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_8_lut_LC_3_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45634\,
            in2 => \N__23601\,
            in3 => \N__21804\,
            lcout => \nx.n3071\,
            ltout => OPEN,
            carryin => \nx.n10867\,
            carryout => \nx.n10868\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_9_lut_LC_3_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45092\,
            in2 => \N__31734\,
            in3 => \N__22110\,
            lcout => \nx.n3070\,
            ltout => OPEN,
            carryin => \nx.n10868\,
            carryout => \nx.n10869\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_10_lut_LC_3_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45392\,
            in2 => \N__23535\,
            in3 => \N__22095\,
            lcout => \nx.n3069\,
            ltout => OPEN,
            carryin => \bfn_3_27_0_\,
            carryout => \nx.n10870\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_11_lut_LC_3_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45399\,
            in2 => \N__22092\,
            in3 => \N__22053\,
            lcout => \nx.n3068\,
            ltout => OPEN,
            carryin => \nx.n10870\,
            carryout => \nx.n10871\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_12_lut_LC_3_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45393\,
            in2 => \N__23391\,
            in3 => \N__22041\,
            lcout => \nx.n3067\,
            ltout => OPEN,
            carryin => \nx.n10871\,
            carryout => \nx.n10872\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_13_lut_LC_3_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45400\,
            in2 => \N__22038\,
            in3 => \N__21999\,
            lcout => \nx.n3066\,
            ltout => OPEN,
            carryin => \nx.n10872\,
            carryout => \nx.n10873\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_14_lut_LC_3_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45394\,
            in2 => \N__23160\,
            in3 => \N__21984\,
            lcout => \nx.n3065\,
            ltout => OPEN,
            carryin => \nx.n10873\,
            carryout => \nx.n10874\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_15_lut_LC_3_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45401\,
            in2 => \N__23318\,
            in3 => \N__21966\,
            lcout => \nx.n3064\,
            ltout => OPEN,
            carryin => \nx.n10874\,
            carryout => \nx.n10875\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_16_lut_LC_3_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45395\,
            in2 => \N__23355\,
            in3 => \N__21948\,
            lcout => \nx.n3063\,
            ltout => OPEN,
            carryin => \nx.n10875\,
            carryout => \nx.n10876\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_17_lut_LC_3_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27503\,
            in2 => \N__45670\,
            in3 => \N__21945\,
            lcout => \nx.n3062\,
            ltout => OPEN,
            carryin => \nx.n10876\,
            carryout => \nx.n10877\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_18_lut_LC_3_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23729\,
            in2 => \N__45631\,
            in3 => \N__22179\,
            lcout => \nx.n3061\,
            ltout => OPEN,
            carryin => \bfn_3_28_0_\,
            carryout => \nx.n10878\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_19_lut_LC_3_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45322\,
            in2 => \N__25848\,
            in3 => \N__22176\,
            lcout => \nx.n3060\,
            ltout => OPEN,
            carryin => \nx.n10878\,
            carryout => \nx.n10879\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_20_lut_LC_3_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45504\,
            in2 => \N__23846\,
            in3 => \N__22167\,
            lcout => \nx.n3059\,
            ltout => OPEN,
            carryin => \nx.n10879\,
            carryout => \nx.n10880\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_21_lut_LC_3_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45323\,
            in2 => \N__23709\,
            in3 => \N__22164\,
            lcout => \nx.n3058\,
            ltout => OPEN,
            carryin => \nx.n10880\,
            carryout => \nx.n10881\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_22_lut_LC_3_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45505\,
            in2 => \N__24057\,
            in3 => \N__22161\,
            lcout => \nx.n3057\,
            ltout => OPEN,
            carryin => \nx.n10881\,
            carryout => \nx.n10882\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_23_lut_LC_3_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45324\,
            in2 => \N__23817\,
            in3 => \N__22158\,
            lcout => \nx.n3056\,
            ltout => OPEN,
            carryin => \nx.n10882\,
            carryout => \nx.n10883\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_24_lut_LC_3_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45506\,
            in2 => \N__23577\,
            in3 => \N__22143\,
            lcout => \nx.n3055\,
            ltout => OPEN,
            carryin => \nx.n10883\,
            carryout => \nx.n10884\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_25_lut_LC_3_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45325\,
            in2 => \N__23282\,
            in3 => \N__22128\,
            lcout => \nx.n3054\,
            ltout => OPEN,
            carryin => \nx.n10884\,
            carryout => \nx.n10885\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_26_lut_LC_3_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23456\,
            in2 => \N__45630\,
            in3 => \N__22296\,
            lcout => \nx.n3053\,
            ltout => OPEN,
            carryin => \bfn_3_29_0_\,
            carryout => \nx.n10886\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_27_lut_LC_3_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45317\,
            in2 => \N__23126\,
            in3 => \N__22287\,
            lcout => \nx.n3052\,
            ltout => OPEN,
            carryin => \nx.n10886\,
            carryout => \nx.n10887\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2076_28_lut_LC_3_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__45318\,
            in1 => \N__25605\,
            in2 => \N__27465\,
            in3 => \N__22284\,
            lcout => \nx.n3083\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i17_4_lut_adj_138_LC_3_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24968\,
            in1 => \N__31003\,
            in2 => \N__26559\,
            in3 => \N__36895\,
            lcout => \nx.n45_adj_707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i2_3_lut_adj_36_LC_3_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32708\,
            in2 => \N__22516\,
            in3 => \N__22202\,
            lcout => OPEN,
            ltout => \nx.n11_adj_628_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i8_4_lut_LC_3_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24653\,
            in1 => \N__24635\,
            in2 => \N__22251\,
            in3 => \N__22248\,
            lcout => \nx.n1334\,
            ltout => \nx.n1334_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i945_3_lut_LC_3_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__22242\,
            in1 => \_gnd_net_\,
            in2 => \N__22224\,
            in3 => \N__22221\,
            lcout => \nx.n1406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i880_3_lut_LC_3_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24533\,
            in1 => \N__22215\,
            in2 => \_gnd_net_\,
            in3 => \N__22364\,
            lcout => \nx.n1309\,
            ltout => \nx.n1309_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i947_3_lut_LC_3_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22188\,
            in2 => \N__22182\,
            in3 => \N__24587\,
            lcout => \nx.n1408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i875_3_lut_LC_3_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22416\,
            in2 => \N__22404\,
            in3 => \N__22365\,
            lcout => \nx.n1304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i948_3_lut_LC_3_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22335\,
            in1 => \N__32709\,
            in2 => \_gnd_net_\,
            in3 => \N__24586\,
            lcout => \nx.n1409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_2_lut_LC_3_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24970\,
            in2 => \_gnd_net_\,
            in3 => \N__22329\,
            lcout => \nx.n1477\,
            ltout => OPEN,
            carryin => \bfn_3_31_0_\,
            carryout => \nx.n10582\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_3_lut_LC_3_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28247\,
            in3 => \N__22326\,
            lcout => \nx.n1476\,
            ltout => OPEN,
            carryin => \nx.n10582\,
            carryout => \nx.n10583\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_4_lut_LC_3_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44926\,
            in2 => \N__26791\,
            in3 => \N__22323\,
            lcout => \nx.n1475\,
            ltout => OPEN,
            carryin => \nx.n10583\,
            carryout => \nx.n10584\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_5_lut_LC_3_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44929\,
            in2 => \N__26850\,
            in3 => \N__22320\,
            lcout => \nx.n1474\,
            ltout => OPEN,
            carryin => \nx.n10584\,
            carryout => \nx.n10585\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_6_lut_LC_3_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44927\,
            in2 => \N__26677\,
            in3 => \N__22317\,
            lcout => \nx.n1473\,
            ltout => OPEN,
            carryin => \nx.n10585\,
            carryout => \nx.n10586\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_7_lut_LC_3_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44930\,
            in2 => \N__26721\,
            in3 => \N__22314\,
            lcout => \nx.n1472\,
            ltout => OPEN,
            carryin => \nx.n10586\,
            carryout => \nx.n10587\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_8_lut_LC_3_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44928\,
            in2 => \N__24489\,
            in3 => \N__22311\,
            lcout => \nx.n1471\,
            ltout => OPEN,
            carryin => \nx.n10587\,
            carryout => \nx.n10588\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_9_lut_LC_3_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44931\,
            in2 => \N__26462\,
            in3 => \N__22533\,
            lcout => \nx.n1470\,
            ltout => OPEN,
            carryin => \nx.n10588\,
            carryout => \nx.n10589\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_10_lut_LC_3_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44828\,
            in2 => \N__24903\,
            in3 => \N__22530\,
            lcout => \nx.n1469\,
            ltout => OPEN,
            carryin => \bfn_3_32_0_\,
            carryout => \nx.n10590\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_11_lut_LC_3_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26761\,
            in2 => \N__45279\,
            in3 => \N__22527\,
            lcout => \nx.n1468\,
            ltout => OPEN,
            carryin => \nx.n10590\,
            carryout => \nx.n10591\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1004_12_lut_LC_3_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__44832\,
            in1 => \N__22482\,
            in2 => \N__28203\,
            in3 => \N__22524\,
            lcout => \nx.n1499\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i941_3_lut_LC_3_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22521\,
            in2 => \N__22491\,
            in3 => \N__24590\,
            lcout => \nx.n1402\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6_4_lut_adj_37_LC_3_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22481\,
            in1 => \N__26455\,
            in2 => \N__26765\,
            in3 => \N__24898\,
            lcout => \nx.n16_adj_629\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i31_1_lut_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22424\,
            lcout => \nx.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i30_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22455\,
            in1 => \N__22425\,
            in2 => \_gnd_net_\,
            in3 => \N__28842\,
            lcout => neo_pixel_transmitter_t0_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48399\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_prev_i15_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26651\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => neopxl_color_prev_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i3_1_lut_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22673\,
            lcout => \nx.n31_adj_650\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i18_1_lut_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22706\,
            lcout => \nx.n16_adj_661\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i17_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28843\,
            in2 => \N__22710\,
            in3 => \N__22736\,
            lcout => neo_pixel_transmitter_t0_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i2_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__22674\,
            in1 => \N__22694\,
            in2 => \N__28873\,
            in3 => \_gnd_net_\,
            lcout => neo_pixel_transmitter_t0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i29_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28833\,
            in1 => \N__22661\,
            in2 => \_gnd_net_\,
            in3 => \N__22584\,
            lcout => neo_pixel_transmitter_t0_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i9_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28834\,
            in1 => \N__22631\,
            in2 => \_gnd_net_\,
            in3 => \N__25086\,
            lcout => neo_pixel_transmitter_t0_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i11_1_lut_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22611\,
            lcout => \nx.n23_adj_617\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i30_1_lut_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22583\,
            lcout => \nx.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i11_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22553\,
            in1 => \N__28835\,
            in2 => \_gnd_net_\,
            in3 => \N__22923\,
            lcout => neo_pixel_transmitter_t0_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i21_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28850\,
            in2 => \N__22839\,
            in3 => \N__22970\,
            lcout => neo_pixel_transmitter_t0_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i13_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22899\,
            in1 => \N__22943\,
            in2 => \_gnd_net_\,
            in3 => \N__28855\,
            lcout => neo_pixel_transmitter_t0_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i12_1_lut_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22922\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \nx.n22_adj_618\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i14_1_lut_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22898\,
            lcout => \nx.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i7_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23214\,
            in1 => \N__22877\,
            in2 => \_gnd_net_\,
            in3 => \N__28856\,
            lcout => neo_pixel_transmitter_t0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9312_3_lut_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26647\,
            in1 => \N__23979\,
            in2 => \_gnd_net_\,
            in3 => \N__43160\,
            lcout => \nx.n13159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i22_1_lut_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22835\,
            lcout => \nx.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i25_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22808\,
            in2 => \N__23079\,
            in3 => \N__28851\,
            lcout => neo_pixel_transmitter_t0_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i18_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__23055\,
            in1 => \N__22784\,
            in2 => \N__28875\,
            in3 => \_gnd_net_\,
            lcout => neo_pixel_transmitter_t0_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i29_1_lut_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23006\,
            lcout => \nx.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i26_1_lut_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23075\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \nx.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i19_1_lut_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23054\,
            lcout => \nx.n15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i28_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__23030\,
            in1 => \_gnd_net_\,
            in2 => \N__23010\,
            in3 => \N__28878\,
            lcout => neo_pixel_transmitter_t0_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i18_4_lut_adj_86_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25372\,
            in1 => \N__31906\,
            in2 => \N__30368\,
            in3 => \N__25492\,
            lcout => \nx.n43_adj_677\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i18_4_lut_adj_93_LC_4_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23182\,
            in1 => \N__23143\,
            in2 => \N__23311\,
            in3 => \N__23233\,
            lcout => \nx.n44_adj_681\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2022_3_lut_LC_4_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25452\,
            in2 => \N__25470\,
            in3 => \N__31858\,
            lcout => \nx.n2995\,
            ltout => \nx.n2995_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7_3_lut_adj_94_LC_4_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26171\,
            in2 => \N__22998\,
            in3 => \N__23492\,
            lcout => OPEN,
            ltout => \nx.n33_adj_682_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i22_4_lut_adj_98_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22995\,
            in1 => \N__23386\,
            in2 => \N__22989\,
            in3 => \N__31732\,
            lcout => \nx.n48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2032_3_lut_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25326\,
            in2 => \N__31875\,
            in3 => \N__25346\,
            lcout => \nx.n3005\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i8_1_lut_LC_4_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23213\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \nx.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9508_3_lut_LC_4_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25356\,
            in2 => \N__25382\,
            in3 => \N__31854\,
            lcout => \nx.n3006\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2013_3_lut_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25632\,
            in1 => \N__31838\,
            in2 => \_gnd_net_\,
            in3 => \N__29589\,
            lcout => \nx.n2986\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1958_3_lut_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27173\,
            in2 => \N__27147\,
            in3 => \N__30301\,
            lcout => \nx.n2899\,
            ltout => \nx.n2899_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9504_3_lut_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31837\,
            in2 => \N__23163\,
            in3 => \N__25548\,
            lcout => \nx.n2998\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1953_3_lut_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27285\,
            in2 => \N__27258\,
            in3 => \N__30302\,
            lcout => \nx.n2894\,
            ltout => \nx.n2894_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_adj_87_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29650\,
            in1 => \N__27543\,
            in2 => \N__23130\,
            in3 => \N__29518\,
            lcout => \nx.n40_adj_678\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2012_3_lut_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31839\,
            in2 => \N__29967\,
            in3 => \N__25620\,
            lcout => \nx.n2985\,
            ltout => \nx.n2985_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i14_4_lut_adj_95_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25601\,
            in1 => \N__23263\,
            in2 => \N__23463\,
            in3 => \N__23443\,
            lcout => \nx.n40_adj_683\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i22_4_lut_adj_92_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29450\,
            in1 => \N__29707\,
            in2 => \N__23415\,
            in3 => \N__23361\,
            lcout => OPEN,
            ltout => \nx.n47_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i24_4_lut_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25221\,
            in1 => \N__23403\,
            in2 => \N__23397\,
            in3 => \N__30462\,
            lcout => \nx.n2918\,
            ltout => \nx.n2918_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2027_3_lut_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25245\,
            in2 => \N__23394\,
            in3 => \N__25268\,
            lcout => \nx.n3000\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_3_lut_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27579\,
            in2 => \N__30409\,
            in3 => \N__29956\,
            lcout => \nx.n38_adj_676\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2023_3_lut_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__31834\,
            in1 => \_gnd_net_\,
            in2 => \N__25506\,
            in3 => \N__25479\,
            lcout => \nx.n2996\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9502_3_lut_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__25538\,
            in1 => \_gnd_net_\,
            in2 => \N__25518\,
            in3 => \N__31833\,
            lcout => \nx.n2997\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2018_3_lut_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31836\,
            in1 => \N__29528\,
            in2 => \_gnd_net_\,
            in3 => \N__25680\,
            lcout => \nx.n2991\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2014_3_lut_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25641\,
            in2 => \N__30495\,
            in3 => \N__31835\,
            lcout => \nx.n2987\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9506_3_lut_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25317\,
            in2 => \N__31863\,
            in3 => \N__29451\,
            lcout => \nx.n3004\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2029_3_lut_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30361\,
            in2 => \N__25302\,
            in3 => \N__31822\,
            lcout => \nx.n3002\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2016_3_lut_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__29571\,
            in1 => \_gnd_net_\,
            in2 => \N__31865\,
            in3 => \N__25659\,
            lcout => \nx.n2989\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2017_3_lut_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27542\,
            in2 => \N__25671\,
            in3 => \N__31826\,
            lcout => \nx.n2990\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2015_3_lut_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30144\,
            in2 => \N__31866\,
            in3 => \N__25650\,
            lcout => \nx.n2988\,
            ltout => \nx.n2988_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_adj_100_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24043\,
            in1 => \N__23695\,
            in2 => \N__23550\,
            in3 => \N__23803\,
            lcout => \nx.n41_adj_686\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2021_3_lut_LC_4_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25440\,
            in2 => \N__31864\,
            in3 => \N__29874\,
            lcout => \nx.n2994\,
            ltout => \nx.n2994_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i16_4_lut_adj_97_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23828\,
            in1 => \N__25841\,
            in2 => \N__23538\,
            in3 => \N__23521\,
            lcout => \nx.n42_adj_684\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2036_3_lut_LC_4_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25212\,
            in1 => \N__26134\,
            in2 => \_gnd_net_\,
            in3 => \N__31859\,
            lcout => \nx.n3009\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2019_3_lut_LC_4_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29652\,
            in2 => \N__31876\,
            in3 => \N__25428\,
            lcout => \nx.n2992\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2083_3_lut_LC_4_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__27456\,
            in1 => \_gnd_net_\,
            in2 => \N__23813\,
            in3 => \N__23787\,
            lcout => \nx.n3088\,
            ltout => \nx.n3088_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i17_4_lut_adj_104_LC_4_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24004\,
            in1 => \N__23776\,
            in2 => \N__23751\,
            in3 => \N__24277\,
            lcout => \nx.n44_adj_690\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2088_3_lut_LC_4_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23739\,
            in2 => \N__23730\,
            in3 => \N__27452\,
            lcout => \nx.n3093\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2085_3_lut_LC_4_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23705\,
            in2 => \N__27464\,
            in3 => \N__23682\,
            lcout => \nx.n3090\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_121_LC_4_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101100"
        )
    port map (
            in0 => \N__23673\,
            in1 => \N__27311\,
            in2 => \N__24236\,
            in3 => \N__23661\,
            lcout => \nx.n12355\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_122_LC_4_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__25733\,
            in1 => \N__24237\,
            in2 => \N__23652\,
            in3 => \N__23637\,
            lcout => OPEN,
            ltout => \nx.n12357_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_123_LC_4_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__24238\,
            in1 => \N__25808\,
            in2 => \N__23631\,
            in3 => \N__23628\,
            lcout => OPEN,
            ltout => \nx.n12359_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_124_LC_4_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__25794\,
            in1 => \N__23616\,
            in2 => \N__23604\,
            in3 => \N__24239\,
            lcout => OPEN,
            ltout => \nx.n12361_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_125_LC_4_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__24240\,
            in1 => \N__24303\,
            in2 => \N__24291\,
            in3 => \N__24281\,
            lcout => OPEN,
            ltout => \nx.n12363_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_126_LC_4_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111000"
        )
    port map (
            in0 => \N__24261\,
            in1 => \N__24241\,
            in2 => \N__24249\,
            in3 => \N__24014\,
            lcout => OPEN,
            ltout => \nx.n12365_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_127_LC_4_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__24242\,
            in1 => \N__24101\,
            in2 => \N__24087\,
            in3 => \N__24084\,
            lcout => \nx.n12367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2084_3_lut_LC_4_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24053\,
            in2 => \N__24027\,
            in3 => \N__27463\,
            lcout => \nx.n3089\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.bit_ctr__i0_LC_4_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23959\,
            in2 => \_gnd_net_\,
            in3 => \N__23943\,
            lcout => \nx.bit_ctr_0\,
            ltout => OPEN,
            carryin => \bfn_4_27_0_\,
            carryout => \nx.n10391\,
            clk => \N__48423\,
            ce => \N__24840\,
            sr => \N__24768\
        );

    \nx.bit_ctr__i1_LC_4_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23927\,
            in2 => \_gnd_net_\,
            in3 => \N__23916\,
            lcout => \nx.bit_ctr_1\,
            ltout => OPEN,
            carryin => \nx.n10391\,
            carryout => \nx.n10392\,
            clk => \N__48423\,
            ce => \N__24840\,
            sr => \N__24768\
        );

    \nx.bit_ctr__i2_LC_4_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23903\,
            in2 => \_gnd_net_\,
            in3 => \N__23892\,
            lcout => \nx.bit_ctr_2\,
            ltout => OPEN,
            carryin => \nx.n10392\,
            carryout => \nx.n10393\,
            clk => \N__48423\,
            ce => \N__24840\,
            sr => \N__24768\
        );

    \nx.bit_ctr__i3_LC_4_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23877\,
            in2 => \_gnd_net_\,
            in3 => \N__23850\,
            lcout => \nx.bit_ctr_3\,
            ltout => OPEN,
            carryin => \nx.n10393\,
            carryout => \nx.n10394\,
            clk => \N__48423\,
            ce => \N__24840\,
            sr => \N__24768\
        );

    \nx.bit_ctr__i4_LC_4_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24356\,
            in2 => \_gnd_net_\,
            in3 => \N__24330\,
            lcout => \nx.bit_ctr_4\,
            ltout => OPEN,
            carryin => \nx.n10394\,
            carryout => \nx.n10395\,
            clk => \N__48423\,
            ce => \N__24840\,
            sr => \N__24768\
        );

    \nx.bit_ctr__i5_LC_4_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26170\,
            in2 => \_gnd_net_\,
            in3 => \N__24327\,
            lcout => \nx.bit_ctr_5\,
            ltout => OPEN,
            carryin => \nx.n10395\,
            carryout => \nx.n10396\,
            clk => \N__48423\,
            ce => \N__24840\,
            sr => \N__24768\
        );

    \nx.bit_ctr__i6_LC_4_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26119\,
            in2 => \_gnd_net_\,
            in3 => \N__24324\,
            lcout => \nx.bit_ctr_6\,
            ltout => OPEN,
            carryin => \nx.n10396\,
            carryout => \nx.n10397\,
            clk => \N__48423\,
            ce => \N__24840\,
            sr => \N__24768\
        );

    \nx.bit_ctr__i7_LC_4_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29808\,
            in2 => \_gnd_net_\,
            in3 => \N__24321\,
            lcout => \nx.bit_ctr_7\,
            ltout => OPEN,
            carryin => \nx.n10397\,
            carryout => \nx.n10398\,
            clk => \N__48423\,
            ce => \N__24840\,
            sr => \N__24768\
        );

    \nx.bit_ctr__i8_LC_4_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28523\,
            in2 => \_gnd_net_\,
            in3 => \N__24318\,
            lcout => \nx.bit_ctr_8\,
            ltout => OPEN,
            carryin => \bfn_4_28_0_\,
            carryout => \nx.n10399\,
            clk => \N__48426\,
            ce => \N__24844\,
            sr => \N__24778\
        );

    \nx.bit_ctr__i9_LC_4_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35881\,
            in2 => \_gnd_net_\,
            in3 => \N__24315\,
            lcout => \nx.bit_ctr_9\,
            ltout => OPEN,
            carryin => \nx.n10399\,
            carryout => \nx.n10400\,
            clk => \N__48426\,
            ce => \N__24844\,
            sr => \N__24778\
        );

    \nx.bit_ctr__i10_LC_4_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37859\,
            in2 => \_gnd_net_\,
            in3 => \N__24312\,
            lcout => \nx.bit_ctr_10\,
            ltout => OPEN,
            carryin => \nx.n10400\,
            carryout => \nx.n10401\,
            clk => \N__48426\,
            ce => \N__24844\,
            sr => \N__24778\
        );

    \nx.bit_ctr__i11_LC_4_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41258\,
            in2 => \_gnd_net_\,
            in3 => \N__24309\,
            lcout => \nx.bit_ctr_11\,
            ltout => OPEN,
            carryin => \nx.n10401\,
            carryout => \nx.n10402\,
            clk => \N__48426\,
            ce => \N__24844\,
            sr => \N__24778\
        );

    \nx.bit_ctr__i12_LC_4_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43539\,
            in2 => \_gnd_net_\,
            in3 => \N__24306\,
            lcout => \nx.bit_ctr_12\,
            ltout => OPEN,
            carryin => \nx.n10402\,
            carryout => \nx.n10403\,
            clk => \N__48426\,
            ce => \N__24844\,
            sr => \N__24778\
        );

    \nx.bit_ctr__i13_LC_4_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39828\,
            in2 => \_gnd_net_\,
            in3 => \N__24402\,
            lcout => \nx.bit_ctr_13\,
            ltout => OPEN,
            carryin => \nx.n10403\,
            carryout => \nx.n10404\,
            clk => \N__48426\,
            ce => \N__24844\,
            sr => \N__24778\
        );

    \nx.bit_ctr__i14_LC_4_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36901\,
            in2 => \_gnd_net_\,
            in3 => \N__24399\,
            lcout => \nx.bit_ctr_14\,
            ltout => OPEN,
            carryin => \nx.n10404\,
            carryout => \nx.n10405\,
            clk => \N__48426\,
            ce => \N__24844\,
            sr => \N__24778\
        );

    \nx.bit_ctr__i15_LC_4_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34064\,
            in2 => \_gnd_net_\,
            in3 => \N__24396\,
            lcout => \nx.bit_ctr_15\,
            ltout => OPEN,
            carryin => \nx.n10405\,
            carryout => \nx.n10406\,
            clk => \N__48426\,
            ce => \N__24844\,
            sr => \N__24778\
        );

    \nx.bit_ctr__i16_LC_4_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30096\,
            in2 => \_gnd_net_\,
            in3 => \N__24393\,
            lcout => \nx.bit_ctr_16\,
            ltout => OPEN,
            carryin => \bfn_4_29_0_\,
            carryout => \nx.n10407\,
            clk => \N__48432\,
            ce => \N__24846\,
            sr => \N__24783\
        );

    \nx.bit_ctr__i17_LC_4_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32745\,
            in2 => \_gnd_net_\,
            in3 => \N__24390\,
            lcout => \nx.bit_ctr_17\,
            ltout => OPEN,
            carryin => \nx.n10407\,
            carryout => \nx.n10408\,
            clk => \N__48432\,
            ce => \N__24846\,
            sr => \N__24783\
        );

    \nx.bit_ctr__i18_LC_4_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34952\,
            in2 => \_gnd_net_\,
            in3 => \N__24387\,
            lcout => \nx.bit_ctr_18\,
            ltout => OPEN,
            carryin => \nx.n10408\,
            carryout => \nx.n10409\,
            clk => \N__48432\,
            ce => \N__24846\,
            sr => \N__24783\
        );

    \nx.bit_ctr__i19_LC_4_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30995\,
            in2 => \_gnd_net_\,
            in3 => \N__24384\,
            lcout => \nx.bit_ctr_19\,
            ltout => OPEN,
            carryin => \nx.n10409\,
            carryout => \nx.n10410\,
            clk => \N__48432\,
            ce => \N__24846\,
            sr => \N__24783\
        );

    \nx.bit_ctr__i20_LC_4_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30836\,
            in2 => \_gnd_net_\,
            in3 => \N__24381\,
            lcout => \nx.bit_ctr_20\,
            ltout => OPEN,
            carryin => \nx.n10410\,
            carryout => \nx.n10411\,
            clk => \N__48432\,
            ce => \N__24846\,
            sr => \N__24783\
        );

    \nx.bit_ctr__i21_LC_4_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24969\,
            in2 => \_gnd_net_\,
            in3 => \N__24378\,
            lcout => \nx.bit_ctr_21\,
            ltout => OPEN,
            carryin => \nx.n10411\,
            carryout => \nx.n10412\,
            clk => \N__48432\,
            ce => \N__24846\,
            sr => \N__24783\
        );

    \nx.bit_ctr__i22_LC_4_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32710\,
            in2 => \_gnd_net_\,
            in3 => \N__24468\,
            lcout => \nx.bit_ctr_22\,
            ltout => OPEN,
            carryin => \nx.n10412\,
            carryout => \nx.n10413\,
            clk => \N__48432\,
            ce => \N__24846\,
            sr => \N__24783\
        );

    \nx.bit_ctr__i23_LC_4_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24534\,
            in2 => \_gnd_net_\,
            in3 => \N__24465\,
            lcout => \nx.bit_ctr_23\,
            ltout => OPEN,
            carryin => \nx.n10413\,
            carryout => \nx.n10414\,
            clk => \N__48432\,
            ce => \N__24846\,
            sr => \N__24783\
        );

    \nx.bit_ctr__i24_LC_4_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24444\,
            in2 => \_gnd_net_\,
            in3 => \N__24423\,
            lcout => \nx.bit_ctr_24\,
            ltout => OPEN,
            carryin => \bfn_4_30_0_\,
            carryout => \nx.n10415\,
            clk => \N__48437\,
            ce => \N__24845\,
            sr => \N__24779\
        );

    \nx.bit_ctr__i25_LC_4_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26219\,
            in2 => \_gnd_net_\,
            in3 => \N__24420\,
            lcout => \nx.bit_ctr_25\,
            ltout => OPEN,
            carryin => \nx.n10415\,
            carryout => \nx.n10416\,
            clk => \N__48437\,
            ce => \N__24845\,
            sr => \N__24779\
        );

    \nx.bit_ctr__i26_LC_4_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28056\,
            in2 => \_gnd_net_\,
            in3 => \N__24417\,
            lcout => \nx.bit_ctr_26\,
            ltout => OPEN,
            carryin => \nx.n10416\,
            carryout => \nx.n10417\,
            clk => \N__48437\,
            ce => \N__24845\,
            sr => \N__24779\
        );

    \nx.bit_ctr__i27_LC_4_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27732\,
            in2 => \_gnd_net_\,
            in3 => \N__24414\,
            lcout => \nx.bit_ctr_27\,
            ltout => OPEN,
            carryin => \nx.n10417\,
            carryout => \nx.n10418\,
            clk => \N__48437\,
            ce => \N__24845\,
            sr => \N__24779\
        );

    \nx.bit_ctr__i28_LC_4_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27678\,
            in2 => \_gnd_net_\,
            in3 => \N__24411\,
            lcout => \nx.bit_ctr_28\,
            ltout => OPEN,
            carryin => \nx.n10418\,
            carryout => \nx.n10419\,
            clk => \N__48437\,
            ce => \N__24845\,
            sr => \N__24779\
        );

    \nx.bit_ctr__i29_LC_4_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26504\,
            in2 => \_gnd_net_\,
            in3 => \N__24408\,
            lcout => \nx.bit_ctr_29\,
            ltout => OPEN,
            carryin => \nx.n10419\,
            carryout => \nx.n10420\,
            clk => \N__48437\,
            ce => \N__24845\,
            sr => \N__24779\
        );

    \nx.bit_ctr__i30_LC_4_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26437\,
            in2 => \_gnd_net_\,
            in3 => \N__24405\,
            lcout => \nx.bit_ctr_30\,
            ltout => OPEN,
            carryin => \nx.n10420\,
            carryout => \nx.n10421\,
            clk => \N__48437\,
            ce => \N__24845\,
            sr => \N__24779\
        );

    \nx.bit_ctr__i31_LC_4_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26557\,
            in2 => \_gnd_net_\,
            in3 => \N__24849\,
            lcout => \nx.bit_ctr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48437\,
            ce => \N__24845\,
            sr => \N__24779\
        );

    \nx.mod_5_i946_3_lut_LC_4_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24738\,
            in2 => \N__24708\,
            in3 => \N__24581\,
            lcout => \nx.n1407\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i944_3_lut_LC_4_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24696\,
            in2 => \N__24591\,
            in3 => \N__24687\,
            lcout => \nx.n1405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i942_3_lut_LC_4_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24666\,
            in2 => \N__24657\,
            in3 => \N__24580\,
            lcout => \nx.n1403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i943_3_lut_LC_4_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24636\,
            in2 => \N__24603\,
            in3 => \N__24585\,
            lcout => \nx.n1404\,
            ltout => \nx.n1404_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i3_3_lut_adj_38_LC_4_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24971\,
            in2 => \N__24546\,
            in3 => \N__28243\,
            lcout => \nx.n13_adj_631\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i19_4_lut_adj_137_LC_4_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34074\,
            in1 => \N__24541\,
            in2 => \N__26505\,
            in3 => \N__43548\,
            lcout => \nx.n47_adj_706\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1010_3_lut_LC_4_32_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24488\,
            in2 => \N__28202\,
            in3 => \N__24474\,
            lcout => \nx.n1503\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1016_3_lut_LC_4_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24975\,
            in1 => \N__24939\,
            in2 => \_gnd_net_\,
            in3 => \N__28182\,
            lcout => \nx.n1509\,
            ltout => \nx.n1509_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6448_2_lut_LC_4_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24933\,
            in3 => \N__30837\,
            lcout => \nx.n9672\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i8_3_lut_LC_4_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26792\,
            in2 => \N__26684\,
            in3 => \N__24930\,
            lcout => OPEN,
            ltout => \nx.n18_adj_630_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9_4_lut_LC_4_32_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26719\,
            in1 => \N__26848\,
            in2 => \N__24924\,
            in3 => \N__24921\,
            lcout => \nx.n1433\,
            ltout => \nx.n1433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1008_3_lut_LC_4_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24915\,
            in2 => \N__24906\,
            in3 => \N__24902\,
            lcout => \nx.n1501\,
            ltout => \nx.n1501_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7_4_lut_adj_39_LC_4_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28351\,
            in1 => \N__31016\,
            in2 => \N__24885\,
            in3 => \N__24882\,
            lcout => \nx.n18_adj_632\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i22_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24876\,
            in1 => \N__29276\,
            in2 => \_gnd_net_\,
            in3 => \N__28865\,
            lcout => neo_pixel_transmitter_t0_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48405\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9323_3_lut_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__49091\,
            in1 => \N__47015\,
            in2 => \_gnd_net_\,
            in3 => \N__48993\,
            lcout => n13170,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9324_3_lut_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39149\,
            in1 => \N__47084\,
            in2 => \_gnd_net_\,
            in3 => \N__48992\,
            lcout => n13171,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i19_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__25128\,
            in1 => \N__28866\,
            in2 => \_gnd_net_\,
            in3 => \N__25059\,
            lcout => neo_pixel_transmitter_t0_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_pin_1__bdd_4_lut_9609_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__25101\,
            in1 => \N__25092\,
            in2 => \N__50574\,
            in3 => \N__50356\,
            lcout => n13450,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i10_1_lut_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25085\,
            lcout => \nx.n24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i20_1_lut_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25058\,
            lcout => \nx.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_prev_i6_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40758\,
            lcout => neopxl_color_prev_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6_3_lut_adj_19_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28543\,
            in2 => \N__29069\,
            in3 => \N__31454\,
            lcout => \nx.n29_adj_607\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__25029\,
            in1 => \N__40757\,
            in2 => \N__26652\,
            in3 => \N__25023\,
            lcout => n11_adj_775,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_prev_i13_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28915\,
            lcout => neopxl_color_prev_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i21_1_lut_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25148\,
            lcout => \nx.n13_adj_649\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1896_3_lut_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29033\,
            in2 => \N__29013\,
            in3 => \N__36569\,
            lcout => \nx.n2805\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i20_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25175\,
            in1 => \N__25149\,
            in2 => \_gnd_net_\,
            in3 => \N__28877\,
            lcout => neo_pixel_transmitter_t0_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_adj_26_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27121\,
            in1 => \N__27271\,
            in2 => \N__26953\,
            in3 => \N__29668\,
            lcout => \nx.n39_adj_614\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1891_rep_18_3_lut_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__29244\,
            in1 => \_gnd_net_\,
            in2 => \N__36593\,
            in3 => \N__31599\,
            lcout => \nx.n2800\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1900_3_lut_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28491\,
            in1 => \N__28544\,
            in2 => \_gnd_net_\,
            in3 => \N__36565\,
            lcout => \nx.n2809\,
            ltout => \nx.n2809_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7_3_lut_adj_25_LC_5_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__29826\,
            in1 => \_gnd_net_\,
            in2 => \N__25140\,
            in3 => \N__29890\,
            lcout => OPEN,
            ltout => \nx.n31_adj_613_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i20_4_lut_LC_5_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26986\,
            in1 => \N__27163\,
            in2 => \N__25137\,
            in3 => \N__25134\,
            lcout => \nx.n44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1956_3_lut_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27094\,
            in2 => \N__30303\,
            in3 => \N__27072\,
            lcout => \nx.n2897\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1966_3_lut_LC_5_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__26987\,
            in1 => \_gnd_net_\,
            in2 => \N__26970\,
            in3 => \N__30286\,
            lcout => \nx.n2907\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1963_3_lut_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26892\,
            in2 => \N__26919\,
            in3 => \N__30294\,
            lcout => \nx.n2904\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1955_3_lut_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27059\,
            in2 => \N__30305\,
            in3 => \N__27042\,
            lcout => \nx.n2896\,
            ltout => \nx.n2896_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7_3_lut_adj_84_LC_5_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26135\,
            in2 => \N__25236\,
            in3 => \N__29777\,
            lcout => \nx.n32_adj_674\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1965_3_lut_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__26931\,
            in1 => \_gnd_net_\,
            in2 => \N__30304\,
            in3 => \N__26957\,
            lcout => \nx.n2906\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1960_3_lut_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27186\,
            in2 => \N__27216\,
            in3 => \N__30293\,
            lcout => \nx.n2901\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1957_3_lut_LC_5_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27131\,
            in2 => \N__30306\,
            in3 => \N__27108\,
            lcout => \nx.n2898\,
            ltout => \nx.n2898_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i17_4_lut_adj_85_LC_5_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25342\,
            in1 => \N__25258\,
            in2 => \N__25233\,
            in3 => \N__25415\,
            lcout => OPEN,
            ltout => \nx.n42_adj_675_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i21_4_lut_adj_88_LC_5_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25559\,
            in1 => \N__29872\,
            in2 => \N__25230\,
            in3 => \N__25227\,
            lcout => \nx.n46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_2_lut_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26136\,
            in2 => \_gnd_net_\,
            in3 => \N__25200\,
            lcout => \nx.n2977\,
            ltout => OPEN,
            carryin => \bfn_5_22_0_\,
            carryout => \nx.n10837\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_3_lut_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29781\,
            in3 => \N__25182\,
            lcout => \nx.n2976\,
            ltout => OPEN,
            carryin => \nx.n10837\,
            carryout => \nx.n10838\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_4_lut_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45557\,
            in2 => \N__25419\,
            in3 => \N__25386\,
            lcout => \nx.n2975\,
            ltout => OPEN,
            carryin => \nx.n10838\,
            carryout => \nx.n10839\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_5_lut_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45563\,
            in2 => \N__25383\,
            in3 => \N__25350\,
            lcout => \nx.n2974\,
            ltout => OPEN,
            carryin => \nx.n10839\,
            carryout => \nx.n10840\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_6_lut_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45558\,
            in2 => \N__25347\,
            in3 => \N__25320\,
            lcout => \nx.n2973\,
            ltout => OPEN,
            carryin => \nx.n10840\,
            carryout => \nx.n10841\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_7_lut_LC_5_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29443\,
            in2 => \N__45730\,
            in3 => \N__25308\,
            lcout => \nx.n2972\,
            ltout => OPEN,
            carryin => \nx.n10841\,
            carryout => \nx.n10842\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_8_lut_LC_5_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45562\,
            in2 => \N__31913\,
            in3 => \N__25305\,
            lcout => \nx.n2971\,
            ltout => OPEN,
            carryin => \nx.n10842\,
            carryout => \nx.n10843\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_9_lut_LC_5_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45564\,
            in2 => \N__30369\,
            in3 => \N__25290\,
            lcout => \nx.n2970\,
            ltout => OPEN,
            carryin => \nx.n10843\,
            carryout => \nx.n10844\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_10_lut_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45551\,
            in2 => \N__30410\,
            in3 => \N__25272\,
            lcout => \nx.n2969\,
            ltout => OPEN,
            carryin => \bfn_5_23_0_\,
            carryout => \nx.n10845\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_11_lut_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45659\,
            in2 => \N__25269\,
            in3 => \N__25239\,
            lcout => \nx.n2968\,
            ltout => OPEN,
            carryin => \nx.n10845\,
            carryout => \nx.n10846\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_12_lut_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45552\,
            in2 => \N__29714\,
            in3 => \N__25566\,
            lcout => \nx.n2967\,
            ltout => OPEN,
            carryin => \nx.n10846\,
            carryout => \nx.n10847\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_13_lut_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45660\,
            in2 => \N__25563\,
            in3 => \N__25542\,
            lcout => \nx.n2966\,
            ltout => OPEN,
            carryin => \nx.n10847\,
            carryout => \nx.n10848\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_14_lut_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45553\,
            in2 => \N__25539\,
            in3 => \N__25509\,
            lcout => \nx.n2965\,
            ltout => OPEN,
            carryin => \nx.n10848\,
            carryout => \nx.n10849\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_15_lut_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45661\,
            in2 => \N__25505\,
            in3 => \N__25473\,
            lcout => \nx.n2964\,
            ltout => OPEN,
            carryin => \nx.n10849\,
            carryout => \nx.n10850\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_16_lut_LC_5_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25469\,
            in2 => \N__45753\,
            in3 => \N__25443\,
            lcout => \nx.n2963\,
            ltout => OPEN,
            carryin => \nx.n10850\,
            carryout => \nx.n10851\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_17_lut_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45665\,
            in2 => \N__29873\,
            in3 => \N__25434\,
            lcout => \nx.n2962\,
            ltout => OPEN,
            carryin => \nx.n10851\,
            carryout => \nx.n10852\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_18_lut_LC_5_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45540\,
            in2 => \N__25869\,
            in3 => \N__25431\,
            lcout => \nx.n2961\,
            ltout => OPEN,
            carryin => \bfn_5_24_0_\,
            carryout => \nx.n10853\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_19_lut_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45565\,
            in2 => \N__29651\,
            in3 => \N__25422\,
            lcout => \nx.n2960\,
            ltout => OPEN,
            carryin => \nx.n10853\,
            carryout => \nx.n10854\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_20_lut_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45541\,
            in2 => \N__29529\,
            in3 => \N__25674\,
            lcout => \nx.n2959\,
            ltout => OPEN,
            carryin => \nx.n10854\,
            carryout => \nx.n10855\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_21_lut_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45566\,
            in2 => \N__27541\,
            in3 => \N__25662\,
            lcout => \nx.n2958\,
            ltout => OPEN,
            carryin => \nx.n10855\,
            carryout => \nx.n10856\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_22_lut_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45542\,
            in2 => \N__29570\,
            in3 => \N__25653\,
            lcout => \nx.n2957\,
            ltout => OPEN,
            carryin => \nx.n10856\,
            carryout => \nx.n10857\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_23_lut_LC_5_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45567\,
            in2 => \N__30143\,
            in3 => \N__25644\,
            lcout => \nx.n2956\,
            ltout => OPEN,
            carryin => \nx.n10857\,
            carryout => \nx.n10858\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_24_lut_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45543\,
            in2 => \N__30488\,
            in3 => \N__25635\,
            lcout => \nx.n2955\,
            ltout => OPEN,
            carryin => \nx.n10858\,
            carryout => \nx.n10859\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_25_lut_LC_5_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29585\,
            in2 => \N__45729\,
            in3 => \N__25623\,
            lcout => \nx.n2954\,
            ltout => OPEN,
            carryin => \nx.n10859\,
            carryout => \nx.n10860\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_26_lut_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29966\,
            in2 => \N__45727\,
            in3 => \N__25611\,
            lcout => \nx.n2953\,
            ltout => OPEN,
            carryin => \bfn_5_25_0_\,
            carryout => \nx.n10861\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_2009_27_lut_LC_5_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__45526\,
            in1 => \N__31867\,
            in2 => \N__27578\,
            in3 => \N__25608\,
            lcout => \nx.n2984\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2020_3_lut_LC_5_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__25584\,
            in1 => \_gnd_net_\,
            in2 => \N__31877\,
            in3 => \N__25868\,
            lcout => \nx.n2993\,
            ltout => \nx.n2993_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2087_3_lut_LC_5_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25827\,
            in2 => \N__25815\,
            in3 => \N__27458\,
            lcout => \nx.n3092\,
            ltout => \nx.n3092_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i23_4_lut_adj_106_LC_5_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25793\,
            in1 => \N__25713\,
            in2 => \N__25764\,
            in3 => \N__25761\,
            lcout => \nx.n50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9_2_lut_LC_5_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27307\,
            in3 => \N__25729\,
            lcout => \nx.n36_adj_687\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_736_2_lut_LC_5_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26230\,
            in2 => \_gnd_net_\,
            in3 => \N__25695\,
            lcout => \nx.n1077\,
            ltout => OPEN,
            carryin => \bfn_5_26_0_\,
            carryout => \nx.n10468\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_736_3_lut_LC_5_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26253\,
            in3 => \N__25692\,
            lcout => \nx.n1076\,
            ltout => OPEN,
            carryin => \nx.n10468\,
            carryout => \nx.n10469\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_736_4_lut_LC_5_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26391\,
            in2 => \N__45704\,
            in3 => \N__25689\,
            lcout => \nx.n1075\,
            ltout => OPEN,
            carryin => \nx.n10469\,
            carryout => \nx.n10470\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_736_5_lut_LC_5_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45501\,
            in2 => \N__26316\,
            in3 => \N__25686\,
            lcout => \nx.n1074\,
            ltout => OPEN,
            carryin => \nx.n10470\,
            carryout => \nx.n10471\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_736_6_lut_LC_5_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45525\,
            in2 => \N__27767\,
            in3 => \N__25683\,
            lcout => \nx.n1073\,
            ltout => OPEN,
            carryin => \nx.n10471\,
            carryout => \nx.n10472\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_736_7_lut_LC_5_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45502\,
            in2 => \N__26082\,
            in3 => \N__25983\,
            lcout => \nx.n1072\,
            ltout => OPEN,
            carryin => \nx.n10472\,
            carryout => \nx.n10473\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_736_8_lut_LC_5_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__45503\,
            in1 => \N__26048\,
            in2 => \N__27891\,
            in3 => \N__25980\,
            lcout => \nx.n1103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_2_lut_LC_5_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45497\,
            in2 => \_gnd_net_\,
            in3 => \N__32763\,
            lcout => \nx.n1877\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i18_4_lut_adj_136_LC_5_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35880\,
            in1 => \N__27737\,
            in2 => \N__26235\,
            in3 => \N__37881\,
            lcout => \nx.n46_adj_705\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i742_3_lut_LC_5_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25941\,
            in1 => \N__26390\,
            in2 => \_gnd_net_\,
            in3 => \N__26046\,
            lcout => \nx.n1107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9571_2_lut_LC_5_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27972\,
            in3 => \N__30639\,
            lcout => \nx.n1007\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i740_3_lut_LC_5_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25902\,
            in2 => \N__27768\,
            in3 => \N__26047\,
            lcout => \nx.n1105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1219_3_lut_LC_5_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34887\,
            in2 => \N__34916\,
            in3 => \N__35148\,
            lcout => \nx.n1808\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7853_3_lut_LC_5_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27956\,
            in2 => \N__30645\,
            in3 => \N__27971\,
            lcout => OPEN,
            ltout => \nx.n11617_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i4_4_lut_LC_5_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__26389\,
            in1 => \N__26181\,
            in2 => \N__26364\,
            in3 => \N__27884\,
            lcout => \nx.n1037\,
            ltout => \nx.n1037_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i743_3_lut_LC_5_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26361\,
            in2 => \N__26355\,
            in3 => \N__26249\,
            lcout => \nx.n1108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i741_3_lut_LC_5_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26315\,
            in1 => \N__26301\,
            in2 => \_gnd_net_\,
            in3 => \N__26044\,
            lcout => \nx.n1106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i676_3_lut_LC_5_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__30625\,
            in1 => \N__28023\,
            in2 => \N__28070\,
            in3 => \_gnd_net_\,
            lcout => \nx.n1009\,
            ltout => \nx.n1009_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i2_3_lut_LC_5_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26223\,
            in2 => \N__26184\,
            in3 => \N__26075\,
            lcout => \nx.n7_adj_616\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i16_4_lut_adj_139_LC_5_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27689\,
            in1 => \N__26169\,
            in2 => \N__41268\,
            in3 => \N__26118\,
            lcout => \nx.n44_adj_708\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i672_3_lut_LC_5_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30627\,
            in2 => \N__27939\,
            in3 => \N__27915\,
            lcout => \nx.n1005\,
            ltout => \nx.n1005_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i739_3_lut_LC_5_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26064\,
            in2 => \N__26055\,
            in3 => \N__26045\,
            lcout => \nx.n1104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i675_3_lut_LC_5_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28013\,
            in2 => \N__27999\,
            in3 => \N__30626\,
            lcout => \nx.n1008\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_2_lut_adj_158_LC_5_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27736\,
            in3 => \N__27816\,
            lcout => \nx.n7082\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9585_4_lut_LC_5_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27873\,
            in1 => \N__27853\,
            in2 => \N__27825\,
            in3 => \N__26573\,
            lcout => \nx.n13064\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9228_4_lut_LC_5_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101101001"
        )
    port map (
            in0 => \N__27724\,
            in1 => \N__27674\,
            in2 => \N__27636\,
            in3 => \N__27815\,
            lcout => \nx.n7342\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_2_lut_adj_29_LC_5_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27682\,
            in3 => \N__27631\,
            lcout => OPEN,
            ltout => \nx.n7084_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_27_LC_5_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__27723\,
            in1 => \N__26572\,
            in2 => \N__26373\,
            in3 => \N__27841\,
            lcout => \nx.n838\,
            ltout => \nx.n838_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_3_lut_4_lut_adj_143_LC_5_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111011"
        )
    port map (
            in0 => \N__27728\,
            in1 => \N__28052\,
            in2 => \N__26370\,
            in3 => \N__27983\,
            lcout => OPEN,
            ltout => \nx.n12595_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_adj_28_LC_5_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__27794\,
            in1 => \N__27905\,
            in2 => \N__26367\,
            in3 => \N__27931\,
            lcout => \nx.n10994\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i605_4_lut_LC_5_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000001"
        )
    port map (
            in0 => \N__27872\,
            in1 => \N__27854\,
            in2 => \N__27824\,
            in3 => \N__26574\,
            lcout => \nx.n906\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6377_2_lut_LC_5_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26558\,
            in3 => \N__26428\,
            lcout => \nx.n608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_3_lut_LC_5_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26548\,
            in2 => \N__26438\,
            in3 => \N__26497\,
            lcout => \nx.n9618\,
            ltout => \nx.n9618_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9471_4_lut_4_lut_LC_5_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001001101100"
        )
    port map (
            in0 => \N__26498\,
            in1 => \N__26432\,
            in2 => \N__26613\,
            in3 => \N__26552\,
            lcout => \nx.n708\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7854_rep_2_3_lut_4_lut_LC_5_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101000"
        )
    port map (
            in0 => \N__27666\,
            in1 => \N__26499\,
            in2 => \N__26610\,
            in3 => \N__26518\,
            lcout => \nx.n11738\,
            ltout => \nx.n11738_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_4_lut_LC_5_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__26609\,
            in1 => \N__26522\,
            in2 => \N__26595\,
            in3 => \N__26591\,
            lcout => \nx.n739\,
            ltout => \nx.n739_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i538_3_lut_LC_5_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100101"
        )
    port map (
            in0 => \N__26592\,
            in1 => \_gnd_net_\,
            in2 => \N__26583\,
            in3 => \N__26580\,
            lcout => \nx.n807\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6508_rep_3_2_lut_3_lut_LC_5_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26553\,
            in2 => \N__26523\,
            in3 => \N__26433\,
            lcout => OPEN,
            ltout => \nx.n11771_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9479_4_lut_LC_5_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110010010110"
        )
    port map (
            in0 => \N__27667\,
            in1 => \N__26500\,
            in2 => \N__26475\,
            in3 => \N__27627\,
            lcout => \nx.n11559\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1009_3_lut_LC_5_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26472\,
            in2 => \N__26463\,
            in3 => \N__28186\,
            lcout => \nx.n1502\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i20_4_lut_adj_135_LC_5_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29827\,
            in1 => \N__30846\,
            in2 => \N__30115\,
            in3 => \N__26439\,
            lcout => \nx.n48_adj_704\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1013_3_lut_LC_5_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26849\,
            in2 => \N__26829\,
            in3 => \N__28188\,
            lcout => \nx.n1506\,
            ltout => \nx.n1506_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9_4_lut_adj_40_LC_5_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28279\,
            in1 => \N__28937\,
            in2 => \N__26817\,
            in3 => \N__26814\,
            lcout => \nx.n20_adj_634\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1014_3_lut_LC_5_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26808\,
            in2 => \N__26799\,
            in3 => \N__28187\,
            lcout => \nx.n1507\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1007_3_lut_LC_5_32_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26766\,
            in2 => \N__28207\,
            in3 => \N__26742\,
            lcout => \nx.n1500\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1011_3_lut_LC_5_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__26733\,
            in1 => \_gnd_net_\,
            in2 => \N__28208\,
            in3 => \N__26720\,
            lcout => \nx.n1504\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1012_3_lut_LC_5_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26700\,
            in2 => \N__26688\,
            in3 => \N__28195\,
            lcout => \nx.n1505\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_i15_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100010000"
        )
    port map (
            in0 => \N__50075\,
            in1 => \N__49843\,
            in2 => \N__49600\,
            in3 => \N__26646\,
            lcout => neopxl_color_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1830_3_lut_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35826\,
            in2 => \N__36209\,
            in3 => \N__33441\,
            lcout => \nx.n2707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1823_3_lut_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37668\,
            in2 => \N__33588\,
            in3 => \N__36206\,
            lcout => \nx.n2700\,
            ltout => \nx.n2700_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i17_4_lut_adj_21_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28969\,
            in1 => \N__29032\,
            in2 => \N__26856\,
            in3 => \N__29101\,
            lcout => \nx.n40_adj_609\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1831_3_lut_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35928\,
            in2 => \N__33459\,
            in3 => \N__36199\,
            lcout => \nx.n2708\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1829_3_lut_LC_6_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33426\,
            in2 => \N__36210\,
            in3 => \N__39423\,
            lcout => \nx.n2706\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1892_3_lut_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28953\,
            in2 => \N__28976\,
            in3 => \N__36575\,
            lcout => \nx.n2801\,
            ltout => \nx.n2801_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i18_4_lut_adj_42_LC_6_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27202\,
            in1 => \N__26911\,
            in2 => \N__26853\,
            in3 => \N__27095\,
            lcout => \nx.n42_adj_635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1893_3_lut_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28986\,
            in2 => \N__36590\,
            in3 => \N__31482\,
            lcout => \nx.n2802\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1887_3_lut_LC_6_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31282\,
            in2 => \N__29184\,
            in3 => \N__36550\,
            lcout => \nx.n2796\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1898_3_lut_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__36549\,
            in1 => \N__29082\,
            in2 => \N__29106\,
            in3 => \_gnd_net_\,
            lcout => \nx.n2807\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1890_rep_19_3_lut_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29211\,
            in2 => \N__29232\,
            in3 => \N__36548\,
            lcout => \nx.n2799\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i14_4_lut_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31537\,
            in1 => \N__33853\,
            in2 => \N__31286\,
            in3 => \N__31312\,
            lcout => OPEN,
            ltout => \nx.n37_adj_608_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i19_4_lut_LC_6_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26880\,
            in1 => \N__29167\,
            in2 => \N__26874\,
            in3 => \N__31564\,
            lcout => OPEN,
            ltout => \nx.n42_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i22_4_lut_LC_6_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31491\,
            in1 => \N__26871\,
            in2 => \N__26865\,
            in3 => \N__33978\,
            lcout => \nx.n2720\,
            ltout => \nx.n2720_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1885_3_lut_LC_6_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31538\,
            in2 => \N__26862\,
            in3 => \N__29130\,
            lcout => \nx.n2794\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1886_3_lut_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29171\,
            in2 => \N__29142\,
            in3 => \N__36554\,
            lcout => \nx.n2795\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1879_3_lut_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__31688\,
            in1 => \_gnd_net_\,
            in2 => \N__36591\,
            in3 => \N__29298\,
            lcout => \nx.n2788\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1888_3_lut_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29193\,
            in2 => \N__31515\,
            in3 => \N__36564\,
            lcout => \nx.n2797\,
            ltout => \nx.n2797_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i17_4_lut_adj_49_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36043\,
            in1 => \N__30442\,
            in2 => \N__26859\,
            in3 => \N__29470\,
            lcout => \nx.n41_adj_643\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1889_3_lut_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29202\,
            in2 => \N__33813\,
            in3 => \N__36556\,
            lcout => \nx.n2798\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1897_rep_21_3_lut_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__36560\,
            in1 => \N__29043\,
            in2 => \N__29073\,
            in3 => \_gnd_net_\,
            lcout => \nx.n2806\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1899_rep_16_3_lut_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36555\,
            in2 => \N__29118\,
            in3 => \N__31455\,
            lcout => \nx.n2808\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1894_3_lut_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28995\,
            in2 => \N__36592\,
            in3 => \N__31569\,
            lcout => \nx.n2803\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_2_lut_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29828\,
            in2 => \_gnd_net_\,
            in3 => \N__27030\,
            lcout => \nx.n2877\,
            ltout => OPEN,
            carryin => \bfn_6_21_0_\,
            carryout => \nx.n10813\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_3_lut_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27020\,
            in3 => \N__26991\,
            lcout => \nx.n2876\,
            ltout => OPEN,
            carryin => \nx.n10813\,
            carryout => \nx.n10814\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_4_lut_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45554\,
            in2 => \N__26988\,
            in3 => \N__26961\,
            lcout => \nx.n2875\,
            ltout => OPEN,
            carryin => \nx.n10814\,
            carryout => \nx.n10815\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_5_lut_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45656\,
            in2 => \N__26958\,
            in3 => \N__26925\,
            lcout => \nx.n2874\,
            ltout => OPEN,
            carryin => \nx.n10815\,
            carryout => \nx.n10816\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_6_lut_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45555\,
            in2 => \N__29474\,
            in3 => \N__26922\,
            lcout => \nx.n2873\,
            ltout => OPEN,
            carryin => \nx.n10816\,
            carryout => \nx.n10817\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_7_lut_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45657\,
            in2 => \N__26918\,
            in3 => \N__26886\,
            lcout => \nx.n2872\,
            ltout => OPEN,
            carryin => \nx.n10817\,
            carryout => \nx.n10818\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_8_lut_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45556\,
            in2 => \N__36047\,
            in3 => \N__26883\,
            lcout => \nx.n2871\,
            ltout => OPEN,
            carryin => \nx.n10818\,
            carryout => \nx.n10819\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_9_lut_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45658\,
            in2 => \N__30446\,
            in3 => \N__27219\,
            lcout => \nx.n2870\,
            ltout => OPEN,
            carryin => \nx.n10819\,
            carryout => \nx.n10820\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_10_lut_LC_6_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45547\,
            in2 => \N__27215\,
            in3 => \N__27180\,
            lcout => \nx.n2869\,
            ltout => OPEN,
            carryin => \bfn_6_22_0_\,
            carryout => \nx.n10821\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_11_lut_LC_6_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45645\,
            in2 => \N__29738\,
            in3 => \N__27177\,
            lcout => \nx.n2868\,
            ltout => OPEN,
            carryin => \nx.n10821\,
            carryout => \nx.n10822\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_12_lut_LC_6_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45548\,
            in2 => \N__27174\,
            in3 => \N__27135\,
            lcout => \nx.n2867\,
            ltout => OPEN,
            carryin => \nx.n10822\,
            carryout => \nx.n10823\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_13_lut_LC_6_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45646\,
            in2 => \N__27132\,
            in3 => \N__27102\,
            lcout => \nx.n2866\,
            ltout => OPEN,
            carryin => \nx.n10823\,
            carryout => \nx.n10824\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_14_lut_LC_6_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45549\,
            in2 => \N__27099\,
            in3 => \N__27063\,
            lcout => \nx.n2865\,
            ltout => OPEN,
            carryin => \nx.n10824\,
            carryout => \nx.n10825\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_15_lut_LC_6_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45647\,
            in2 => \N__27060\,
            in3 => \N__27036\,
            lcout => \nx.n2864\,
            ltout => OPEN,
            carryin => \nx.n10825\,
            carryout => \nx.n10826\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_16_lut_LC_6_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45550\,
            in2 => \N__29903\,
            in3 => \N__27033\,
            lcout => \nx.n2863\,
            ltout => OPEN,
            carryin => \nx.n10826\,
            carryout => \nx.n10827\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_17_lut_LC_6_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45648\,
            in2 => \N__27284\,
            in3 => \N__27246\,
            lcout => \nx.n2862\,
            ltout => OPEN,
            carryin => \nx.n10827\,
            carryout => \nx.n10828\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_18_lut_LC_6_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45530\,
            in2 => \N__29681\,
            in3 => \N__27243\,
            lcout => \nx.n2861\,
            ltout => OPEN,
            carryin => \bfn_6_23_0_\,
            carryout => \nx.n10829\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_19_lut_LC_6_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45533\,
            in2 => \N__29427\,
            in3 => \N__27240\,
            lcout => \nx.n2860\,
            ltout => OPEN,
            carryin => \nx.n10829\,
            carryout => \nx.n10830\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_20_lut_LC_6_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45531\,
            in2 => \N__29396\,
            in3 => \N__27237\,
            lcout => \nx.n2859\,
            ltout => OPEN,
            carryin => \nx.n10830\,
            carryout => \nx.n10831\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_21_lut_LC_6_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45534\,
            in2 => \N__29412\,
            in3 => \N__27234\,
            lcout => \nx.n2858\,
            ltout => OPEN,
            carryin => \nx.n10831\,
            carryout => \nx.n10832\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_22_lut_LC_6_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45532\,
            in2 => \N__30329\,
            in3 => \N__27231\,
            lcout => \nx.n2857\,
            ltout => OPEN,
            carryin => \nx.n10832\,
            carryout => \nx.n10833\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_23_lut_LC_6_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45535\,
            in2 => \N__29934\,
            in3 => \N__27228\,
            lcout => \nx.n2856\,
            ltout => OPEN,
            carryin => \nx.n10833\,
            carryout => \nx.n10834\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_24_lut_LC_6_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29618\,
            in2 => \N__45728\,
            in3 => \N__27225\,
            lcout => \nx.n2855\,
            ltout => OPEN,
            carryin => \nx.n10834\,
            carryout => \nx.n10835\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_25_lut_LC_6_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45539\,
            in2 => \N__36465\,
            in3 => \N__27222\,
            lcout => \nx.n2854\,
            ltout => OPEN,
            carryin => \nx.n10835\,
            carryout => \nx.n10836\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1942_26_lut_LC_6_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__45338\,
            in1 => \N__29370\,
            in2 => \N__30283\,
            in3 => \N__27582\,
            lcout => \nx.n2885\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1882_3_lut_LC_6_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29325\,
            in2 => \N__33906\,
            in3 => \N__36595\,
            lcout => \nx.n2791\,
            ltout => \nx.n2791_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1949_3_lut_LC_6_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__30246\,
            in1 => \N__27558\,
            in2 => \N__27552\,
            in3 => \_gnd_net_\,
            lcout => \nx.n2890\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1819_3_lut_LC_6_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33753\,
            in2 => \N__37704\,
            in3 => \N__36208\,
            lcout => \nx.n2696\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1950_3_lut_LC_6_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29397\,
            in2 => \N__30284\,
            in3 => \N__27549\,
            lcout => \nx.n2891\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1880_3_lut_LC_6_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36594\,
            in2 => \N__31668\,
            in3 => \N__29310\,
            lcout => \nx.n2789\,
            ltout => \nx.n2789_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1947_3_lut_LC_6_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__30250\,
            in1 => \N__27513\,
            in2 => \N__27507\,
            in3 => \_gnd_net_\,
            lcout => \nx.n2888\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_2_lut_LC_6_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30573\,
            in3 => \N__30519\,
            lcout => \nx.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2089_3_lut_LC_6_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27504\,
            in2 => \N__27480\,
            in3 => \N__27457\,
            lcout => \nx.n3094\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_4_lut_adj_64_LC_6_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30547\,
            in1 => \N__30687\,
            in2 => \N__27777\,
            in3 => \N__32409\,
            lcout => OPEN,
            ltout => \nx.n28_adj_660_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i14_4_lut_adj_81_LC_6_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32449\,
            in1 => \N__27594\,
            in2 => \N__27609\,
            in3 => \N__27606\,
            lcout => \nx.n1928\,
            ltout => \nx.n1928_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9586_1_lut_LC_6_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27600\,
            in3 => \_gnd_net_\,
            lcout => \nx.n13435\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1283_3_lut_LC_6_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32538\,
            in2 => \N__32511\,
            in3 => \N__32887\,
            lcout => \nx.n1904\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1287_3_lut_LC_6_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__32643\,
            in1 => \_gnd_net_\,
            in2 => \N__32900\,
            in3 => \N__32662\,
            lcout => \nx.n1908\,
            ltout => \nx.n1908_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9_4_lut_adj_55_LC_6_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30658\,
            in1 => \N__30007\,
            in2 => \N__27597\,
            in3 => \N__32356\,
            lcout => \nx.n24_adj_648\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1286_3_lut_LC_6_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32607\,
            in2 => \N__32899\,
            in3 => \N__32624\,
            lcout => \nx.n1907\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1288_3_lut_LC_6_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27588\,
            in1 => \N__32764\,
            in2 => \_gnd_net_\,
            in3 => \N__32874\,
            lcout => \nx.n1909\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_4_lut_adj_16_LC_6_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32588\,
            in1 => \N__32623\,
            in2 => \N__32400\,
            in3 => \N__27744\,
            lcout => \nx.n1829\,
            ltout => \nx.n1829_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1282_3_lut_LC_6_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__32486\,
            in1 => \N__32472\,
            in2 => \N__27783\,
            in3 => \_gnd_net_\,
            lcout => \nx.n1903\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1285_3_lut_LC_6_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__32878\,
            in1 => \_gnd_net_\,
            in2 => \N__32592\,
            in3 => \N__32568\,
            lcout => \nx.n1906\,
            ltout => \nx.n1906_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7_3_lut_LC_6_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30108\,
            in2 => \N__27780\,
            in3 => \N__30061\,
            lcout => \nx.n22_adj_605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9569_2_lut_LC_6_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27957\,
            in3 => \N__30643\,
            lcout => \nx.n1006\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1215_3_lut_LC_6_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34716\,
            in2 => \N__34749\,
            in3 => \N__35151\,
            lcout => \nx.n1804\,
            ltout => \nx.n1804_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5_3_lut_adj_132_LC_6_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32769\,
            in2 => \N__27750\,
            in3 => \N__32666\,
            lcout => OPEN,
            ltout => \nx.n19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i12_4_lut_adj_15_LC_6_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34613\,
            in1 => \N__32530\,
            in2 => \N__27747\,
            in3 => \N__30861\,
            lcout => \nx.n26_adj_600\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i2045_2_lut_3_lut_LC_6_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27738\,
            in2 => \N__27690\,
            in3 => \N__27635\,
            lcout => \nx.n5260\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1278_3_lut_LC_6_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__33020\,
            in1 => \_gnd_net_\,
            in2 => \N__33000\,
            in3 => \N__32882\,
            lcout => \nx.n1899\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_669_2_lut_LC_6_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28071\,
            in3 => \N__28017\,
            lcout => \nx.n977\,
            ltout => OPEN,
            carryin => \bfn_6_28_0_\,
            carryout => \nx.n10474\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_669_3_lut_LC_6_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28014\,
            in3 => \N__27990\,
            lcout => \nx.n976\,
            ltout => OPEN,
            carryin => \nx.n10474\,
            carryout => \nx.n10475\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_669_4_lut_LC_6_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45099\,
            in2 => \N__27987\,
            in3 => \N__27960\,
            lcout => \nx.n975\,
            ltout => OPEN,
            carryin => \nx.n10475\,
            carryout => \nx.n10476\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_669_5_lut_LC_6_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45104\,
            in2 => \N__27798\,
            in3 => \N__27942\,
            lcout => \nx.n974\,
            ltout => OPEN,
            carryin => \nx.n10476\,
            carryout => \nx.n10477\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_669_6_lut_LC_6_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45100\,
            in2 => \N__27938\,
            in3 => \N__27909\,
            lcout => \nx.n973\,
            ltout => OPEN,
            carryin => \nx.n10477\,
            carryout => \nx.n10478\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_669_7_lut_LC_6_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__27906\,
            in1 => \N__30597\,
            in2 => \N__45496\,
            in3 => \N__27894\,
            lcout => \nx.n4_adj_596\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1152_3_lut_LC_6_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30957\,
            in1 => \N__31005\,
            in2 => \_gnd_net_\,
            in3 => \N__34480\,
            lcout => \nx.n1709\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i606_3_lut_LC_6_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27871\,
            in2 => \N__27855\,
            in3 => \N__27823\,
            lcout => \nx.n11674\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i10_4_lut_adj_41_LC_6_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28475\,
            in1 => \N__28143\,
            in2 => \N__28398\,
            in3 => \N__28098\,
            lcout => \nx.n1532\,
            ltout => \nx.n1532_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1078_3_lut_LC_6_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28397\,
            in2 => \N__28089\,
            in3 => \N__28371\,
            lcout => \nx.n1603\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1081_3_lut_LC_6_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__28476\,
            in1 => \_gnd_net_\,
            in2 => \N__28455\,
            in3 => \N__33263\,
            lcout => \nx.n1606\,
            ltout => \nx.n1606_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i10_4_lut_adj_54_LC_6_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31156\,
            in1 => \N__28077\,
            in2 => \N__28086\,
            in3 => \N__30801\,
            lcout => OPEN,
            ltout => \nx.n22_adj_647_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i11_4_lut_adj_80_LC_6_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33172\,
            in1 => \N__30910\,
            in2 => \N__28083\,
            in3 => \N__33321\,
            lcout => \nx.n1631\,
            ltout => \nx.n1631_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1147_3_lut_LC_6_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33203\,
            in2 => \N__28080\,
            in3 => \N__30876\,
            lcout => \nx.n1704\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1082_3_lut_LC_6_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28110\,
            in2 => \N__28128\,
            in3 => \N__33262\,
            lcout => \nx.n1607\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1079_3_lut_LC_6_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__28410\,
            in1 => \_gnd_net_\,
            in2 => \N__33275\,
            in3 => \N__28437\,
            lcout => \nx.n1604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7_4_lut_LC_6_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31109\,
            in1 => \N__33385\,
            in2 => \N__31070\,
            in3 => \N__31089\,
            lcout => \nx.n19_adj_602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1076_3_lut_LC_6_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28355\,
            in2 => \N__33272\,
            in3 => \N__28335\,
            lcout => \nx.n1601\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1075_3_lut_LC_6_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__28323\,
            in1 => \_gnd_net_\,
            in2 => \N__28302\,
            in3 => \N__33255\,
            lcout => \nx.n1600\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1015_3_lut_LC_6_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28248\,
            in2 => \N__28224\,
            in3 => \N__28209\,
            lcout => \nx.n1508\,
            ltout => \nx.n1508_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5_2_lut_LC_6_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28146\,
            in3 => \N__28433\,
            lcout => \nx.n16_adj_633\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i7_3_lut_adj_91_LC_6_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35063\,
            in2 => \N__35425\,
            in3 => \N__35185\,
            lcout => \nx.n20_adj_680\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1074_3_lut_LC_6_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28287\,
            in2 => \N__28263\,
            in3 => \N__33251\,
            lcout => \nx.n1599\,
            ltout => \nx.n1599_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1141_3_lut_LC_6_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34499\,
            in2 => \N__28137\,
            in3 => \N__31098\,
            lcout => \nx.n1698\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_2_lut_LC_6_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30845\,
            in2 => \_gnd_net_\,
            in3 => \N__28134\,
            lcout => \nx.n1577\,
            ltout => OPEN,
            carryin => \bfn_6_31_0_\,
            carryout => \nx.n10592\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_3_lut_LC_6_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33362\,
            in3 => \N__28131\,
            lcout => \nx.n1576\,
            ltout => OPEN,
            carryin => \nx.n10592\,
            carryout => \nx.n10593\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_4_lut_LC_6_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44869\,
            in2 => \N__28127\,
            in3 => \N__28101\,
            lcout => \nx.n1575\,
            ltout => OPEN,
            carryin => \nx.n10593\,
            carryout => \nx.n10594\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_5_lut_LC_6_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44923\,
            in2 => \N__28474\,
            in3 => \N__28443\,
            lcout => \nx.n1574\,
            ltout => OPEN,
            carryin => \nx.n10594\,
            carryout => \nx.n10595\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_6_lut_LC_6_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44870\,
            in2 => \N__33308\,
            in3 => \N__28440\,
            lcout => \nx.n1573\,
            ltout => OPEN,
            carryin => \nx.n10595\,
            carryout => \nx.n10596\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_7_lut_LC_6_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44924\,
            in2 => \N__28432\,
            in3 => \N__28401\,
            lcout => \nx.n1572\,
            ltout => OPEN,
            carryin => \nx.n10596\,
            carryout => \nx.n10597\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_8_lut_LC_6_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44871\,
            in2 => \N__28393\,
            in3 => \N__28362\,
            lcout => \nx.n1571\,
            ltout => OPEN,
            carryin => \nx.n10597\,
            carryout => \nx.n10598\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_9_lut_LC_6_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44925\,
            in2 => \N__31032\,
            in3 => \N__28359\,
            lcout => \nx.n1570\,
            ltout => OPEN,
            carryin => \nx.n10598\,
            carryout => \nx.n10599\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_10_lut_LC_6_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44483\,
            in2 => \N__28356\,
            in3 => \N__28326\,
            lcout => \nx.n1569\,
            ltout => OPEN,
            carryin => \bfn_6_32_0_\,
            carryout => \nx.n10600\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_11_lut_LC_6_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44486\,
            in2 => \N__28322\,
            in3 => \N__28290\,
            lcout => \nx.n1568\,
            ltout => OPEN,
            carryin => \nx.n10600\,
            carryout => \nx.n10601\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_12_lut_LC_6_32_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44484\,
            in2 => \N__28286\,
            in3 => \N__28251\,
            lcout => \nx.n1567\,
            ltout => OPEN,
            carryin => \nx.n10601\,
            carryout => \nx.n10602\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1071_13_lut_LC_6_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__44485\,
            in1 => \N__28941\,
            in2 => \N__33276\,
            in3 => \N__28920\,
            lcout => \nx.n1598\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i0_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__31254\,
            in1 => \N__35472\,
            in2 => \N__28613\,
            in3 => \N__46536\,
            lcout => pin_out_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48411\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1825_3_lut_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__36687\,
            in1 => \_gnd_net_\,
            in2 => \N__33615\,
            in3 => \N__36207\,
            lcout => \nx.n2702\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_i13_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111100000100"
        )
    port map (
            in0 => \N__49842\,
            in1 => \N__49593\,
            in2 => \N__50077\,
            in3 => \N__28897\,
            lcout => neopxl_color_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48406\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.neo_pixel_transmitter_t0_i0_i0_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28874\,
            in1 => \N__28673\,
            in2 => \_gnd_net_\,
            in3 => \N__28647\,
            lcout => neo_pixel_transmitter_t0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48406\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i1_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__31242\,
            in1 => \N__33105\,
            in2 => \N__28571\,
            in3 => \N__46515\,
            lcout => pin_out_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48406\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i1_1_lut_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28646\,
            lcout => \nx.n33_adj_652\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9299_3_lut_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28612\,
            in1 => \N__28564\,
            in2 => \_gnd_net_\,
            in3 => \N__49041\,
            lcout => n13146,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_2_lut_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28548\,
            in2 => \_gnd_net_\,
            in3 => \N__28479\,
            lcout => \nx.n2777\,
            ltout => OPEN,
            carryin => \bfn_7_19_0_\,
            carryout => \nx.n10790\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_3_lut_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31453\,
            in3 => \N__29109\,
            lcout => \nx.n2776\,
            ltout => OPEN,
            carryin => \nx.n10790\,
            carryout => \nx.n10791\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_4_lut_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45695\,
            in2 => \N__29105\,
            in3 => \N__29076\,
            lcout => \nx.n2775\,
            ltout => OPEN,
            carryin => \nx.n10791\,
            carryout => \nx.n10792\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_5_lut_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45698\,
            in2 => \N__29068\,
            in3 => \N__29037\,
            lcout => \nx.n2774\,
            ltout => OPEN,
            carryin => \nx.n10792\,
            carryout => \nx.n10793\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_6_lut_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45696\,
            in2 => \N__29034\,
            in3 => \N__29001\,
            lcout => \nx.n2773\,
            ltout => OPEN,
            carryin => \nx.n10793\,
            carryout => \nx.n10794\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_7_lut_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45699\,
            in2 => \N__36081\,
            in3 => \N__28998\,
            lcout => \nx.n2772\,
            ltout => OPEN,
            carryin => \nx.n10794\,
            carryout => \nx.n10795\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_8_lut_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45697\,
            in2 => \N__31568\,
            in3 => \N__28989\,
            lcout => \nx.n2771\,
            ltout => OPEN,
            carryin => \nx.n10795\,
            carryout => \nx.n10796\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_9_lut_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45700\,
            in2 => \N__31481\,
            in3 => \N__28980\,
            lcout => \nx.n2770\,
            ltout => OPEN,
            carryin => \nx.n10796\,
            carryout => \nx.n10797\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_10_lut_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45016\,
            in2 => \N__28977\,
            in3 => \N__28944\,
            lcout => \nx.n2769\,
            ltout => OPEN,
            carryin => \bfn_7_20_0_\,
            carryout => \nx.n10798\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_11_lut_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45649\,
            in2 => \N__31598\,
            in3 => \N__29235\,
            lcout => \nx.n2768\,
            ltout => OPEN,
            carryin => \nx.n10798\,
            carryout => \nx.n10799\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_12_lut_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45017\,
            in2 => \N__29231\,
            in3 => \N__29205\,
            lcout => \nx.n2767\,
            ltout => OPEN,
            carryin => \nx.n10799\,
            carryout => \nx.n10800\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_13_lut_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45650\,
            in2 => \N__33809\,
            in3 => \N__29196\,
            lcout => \nx.n2766\,
            ltout => OPEN,
            carryin => \nx.n10800\,
            carryout => \nx.n10801\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_14_lut_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31511\,
            in2 => \N__45752\,
            in3 => \N__29187\,
            lcout => \nx.n2765\,
            ltout => OPEN,
            carryin => \nx.n10801\,
            carryout => \nx.n10802\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_15_lut_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45654\,
            in2 => \N__31287\,
            in3 => \N__29175\,
            lcout => \nx.n2764\,
            ltout => OPEN,
            carryin => \nx.n10802\,
            carryout => \nx.n10803\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_16_lut_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45018\,
            in2 => \N__29172\,
            in3 => \N__29133\,
            lcout => \nx.n2763\,
            ltout => OPEN,
            carryin => \nx.n10803\,
            carryout => \nx.n10804\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_17_lut_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45655\,
            in2 => \N__31542\,
            in3 => \N__29124\,
            lcout => \nx.n2762\,
            ltout => OPEN,
            carryin => \nx.n10804\,
            carryout => \nx.n10805\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_18_lut_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31316\,
            in2 => \N__45751\,
            in3 => \N__29121\,
            lcout => \nx.n2761\,
            ltout => OPEN,
            carryin => \bfn_7_21_0_\,
            carryout => \nx.n10806\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_19_lut_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45642\,
            in2 => \N__33858\,
            in3 => \N__29328\,
            lcout => \nx.n2760\,
            ltout => OPEN,
            carryin => \nx.n10806\,
            carryout => \nx.n10807\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_20_lut_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45691\,
            in2 => \N__33902\,
            in3 => \N__29316\,
            lcout => \nx.n2759\,
            ltout => OPEN,
            carryin => \nx.n10807\,
            carryout => \nx.n10808\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_21_lut_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45643\,
            in2 => \N__31628\,
            in3 => \N__29313\,
            lcout => \nx.n2758\,
            ltout => OPEN,
            carryin => \nx.n10808\,
            carryout => \nx.n10809\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_22_lut_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45692\,
            in2 => \N__31667\,
            in3 => \N__29301\,
            lcout => \nx.n2757\,
            ltout => OPEN,
            carryin => \nx.n10809\,
            carryout => \nx.n10810\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_23_lut_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45644\,
            in2 => \N__31692\,
            in3 => \N__29292\,
            lcout => \nx.n2756\,
            ltout => OPEN,
            carryin => \nx.n10810\,
            carryout => \nx.n10811\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_24_lut_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45693\,
            in2 => \N__36636\,
            in3 => \N__29289\,
            lcout => \nx.n2755\,
            ltout => OPEN,
            carryin => \nx.n10811\,
            carryout => \nx.n10812\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1875_25_lut_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__45694\,
            in1 => \N__36601\,
            in2 => \N__33789\,
            in3 => \N__29286\,
            lcout => \nx.n2786\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9_4_lut_adj_70_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32182\,
            in1 => \N__34375\,
            in2 => \N__34339\,
            in3 => \N__32129\,
            lcout => \nx.n25_adj_666\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.sub_14_inv_0_i23_1_lut_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29283\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \nx.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1884_3_lut_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__31317\,
            in1 => \N__36596\,
            in2 => \N__29547\,
            in3 => \_gnd_net_\,
            lcout => \nx.n2793\,
            ltout => \nx.n2793_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1951_3_lut_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29538\,
            in2 => \N__29532\,
            in3 => \N__30251\,
            lcout => \nx.n2892\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1881_3_lut_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__29493\,
            in1 => \_gnd_net_\,
            in2 => \N__31629\,
            in3 => \N__36600\,
            lcout => \nx.n2790\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1883_3_lut_LC_7_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__33857\,
            in1 => \_gnd_net_\,
            in2 => \N__36605\,
            in3 => \N__29487\,
            lcout => \nx.n2792\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9505_3_lut_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29481\,
            in2 => \N__30285\,
            in3 => \N__29475\,
            lcout => \nx.n2905\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_4_lut_adj_63_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41060\,
            in1 => \N__41153\,
            in2 => \N__41427\,
            in3 => \N__43199\,
            lcout => \nx.n33_adj_659\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i14_4_lut_adj_33_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29423\,
            in1 => \N__29408\,
            in2 => \N__29395\,
            in3 => \N__30322\,
            lcout => OPEN,
            ltout => \nx.n38_adj_625_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i19_4_lut_adj_43_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29369\,
            in1 => \N__36457\,
            in2 => \N__29355\,
            in3 => \N__29916\,
            lcout => OPEN,
            ltout => \nx.n43_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i23_4_lut_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29352\,
            in1 => \N__29340\,
            in2 => \N__29331\,
            in3 => \N__29988\,
            lcout => \nx.n2819\,
            ltout => \nx.n2819_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1945_3_lut_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__29976\,
            in1 => \_gnd_net_\,
            in2 => \N__29970\,
            in3 => \N__36458\,
            lcout => \nx.n2886\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i2_2_lut_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29933\,
            in3 => \N__29617\,
            lcout => \nx.n26_adj_615\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1954_3_lut_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29910\,
            in2 => \N__30255\,
            in3 => \N__29904\,
            lcout => \nx.n2895\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1968_3_lut_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29841\,
            in1 => \N__29829\,
            in2 => \_gnd_net_\,
            in3 => \N__30211\,
            lcout => \nx.n2909\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1959_3_lut_LC_7_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29745\,
            in2 => \N__30256\,
            in3 => \N__29739\,
            lcout => \nx.n2900\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1952_3_lut_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29688\,
            in2 => \N__30275\,
            in3 => \N__29682\,
            lcout => \nx.n2893\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1946_3_lut_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29619\,
            in2 => \N__30277\,
            in3 => \N__29595\,
            lcout => \nx.n2887\,
            ltout => \nx.n2887_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i14_4_lut_adj_90_LC_7_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29563\,
            in1 => \N__30481\,
            in2 => \N__30465\,
            in3 => \N__30130\,
            lcout => \nx.n39_adj_679\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1961_3_lut_LC_7_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30450\,
            in2 => \N__30274\,
            in3 => \N__30423\,
            lcout => \nx.n2902\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1962_3_lut_LC_7_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30378\,
            in2 => \N__36048\,
            in3 => \N__30227\,
            lcout => \nx.n2903\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1948_3_lut_LC_7_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30330\,
            in2 => \N__30276\,
            in3 => \N__30150\,
            lcout => \nx.n2889\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i12_4_lut_adj_67_LC_7_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31984\,
            in1 => \N__34276\,
            in2 => \N__32089\,
            in3 => \N__32032\,
            lcout => \nx.n28_adj_663\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_2_lut_LC_7_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__30117\,
            in1 => \N__30116\,
            in2 => \N__30044\,
            in3 => \N__30066\,
            lcout => \nx.n2009\,
            ltout => OPEN,
            carryin => \bfn_7_25_0_\,
            carryout => \nx.n10642\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_3_lut_LC_7_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__30063\,
            in1 => \N__30062\,
            in2 => \N__30045\,
            in3 => \N__30027\,
            lcout => \nx.n2008\,
            ltout => OPEN,
            carryin => \nx.n10642\,
            carryout => \nx.n10643\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_4_lut_LC_7_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__30024\,
            in1 => \N__30023\,
            in2 => \N__30773\,
            in3 => \N__30012\,
            lcout => \nx.n2007\,
            ltout => OPEN,
            carryin => \nx.n10643\,
            carryout => \nx.n10644\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_5_lut_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__30009\,
            in1 => \N__30008\,
            in2 => \N__30776\,
            in3 => \N__29991\,
            lcout => \nx.n2006\,
            ltout => OPEN,
            carryin => \nx.n10644\,
            carryout => \nx.n10645\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_6_lut_LC_7_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__30591\,
            in1 => \N__30590\,
            in2 => \N__30774\,
            in3 => \N__30579\,
            lcout => \nx.n2005\,
            ltout => OPEN,
            carryin => \nx.n10645\,
            carryout => \nx.n10646\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_7_lut_LC_7_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__32430\,
            in1 => \N__32429\,
            in2 => \N__30777\,
            in3 => \N__30576\,
            lcout => \nx.n2004\,
            ltout => OPEN,
            carryin => \nx.n10646\,
            carryout => \nx.n10647\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_8_lut_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__30572\,
            in1 => \N__30571\,
            in2 => \N__30775\,
            in3 => \N__30552\,
            lcout => \nx.n2003\,
            ltout => OPEN,
            carryin => \nx.n10647\,
            carryout => \nx.n10648\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_9_lut_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__30549\,
            in1 => \N__30548\,
            in2 => \N__30778\,
            in3 => \N__30531\,
            lcout => \nx.n2002\,
            ltout => OPEN,
            carryin => \nx.n10648\,
            carryout => \nx.n10649\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_10_lut_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__30666\,
            in1 => \N__30665\,
            in2 => \N__30779\,
            in3 => \N__30528\,
            lcout => \nx.n2001\,
            ltout => OPEN,
            carryin => \bfn_7_26_0_\,
            carryout => \nx.n10650\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_11_lut_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__32457\,
            in1 => \N__32456\,
            in2 => \N__30783\,
            in3 => \N__30525\,
            lcout => \nx.n2000\,
            ltout => OPEN,
            carryin => \nx.n10650\,
            carryout => \nx.n10651\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_12_lut_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__32388\,
            in1 => \N__32387\,
            in2 => \N__30780\,
            in3 => \N__30522\,
            lcout => \nx.n1999\,
            ltout => OPEN,
            carryin => \nx.n10651\,
            carryout => \nx.n10652\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_13_lut_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__30518\,
            in1 => \N__30517\,
            in2 => \N__30784\,
            in3 => \N__30498\,
            lcout => \nx.n1998\,
            ltout => OPEN,
            carryin => \nx.n10652\,
            carryout => \nx.n10653\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_14_lut_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__32364\,
            in1 => \N__32363\,
            in2 => \N__30781\,
            in3 => \N__30795\,
            lcout => \nx.n1997\,
            ltout => OPEN,
            carryin => \nx.n10653\,
            carryout => \nx.n10654\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_15_lut_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__30686\,
            in1 => \N__30685\,
            in2 => \N__30785\,
            in3 => \N__30792\,
            lcout => \nx.n1996\,
            ltout => OPEN,
            carryin => \nx.n10654\,
            carryout => \nx.n10655\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_16_lut_LC_7_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__32793\,
            in1 => \N__32792\,
            in2 => \N__30782\,
            in3 => \N__30789\,
            lcout => \nx.n1995\,
            ltout => OPEN,
            carryin => \nx.n10655\,
            carryout => \nx.n10656\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1339_17_lut_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__32819\,
            in1 => \N__32820\,
            in2 => \N__30786\,
            in3 => \N__30690\,
            lcout => \nx.n1994\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1220_3_lut_LC_7_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34932\,
            in1 => \N__34976\,
            in2 => \_gnd_net_\,
            in3 => \N__35149\,
            lcout => \nx.n1809\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i4_3_lut_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41279\,
            in2 => \N__41208\,
            in3 => \N__41883\,
            lcout => \nx.n24_adj_654\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1216_3_lut_LC_7_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34764\,
            in1 => \N__34780\,
            in2 => \_gnd_net_\,
            in3 => \N__35150\,
            lcout => \nx.n1805\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1276_3_lut_LC_7_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34578\,
            in2 => \N__32901\,
            in3 => \N__32955\,
            lcout => \nx.n1897\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1281_3_lut_LC_7_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__32883\,
            in1 => \N__33087\,
            in2 => \N__34617\,
            in3 => \_gnd_net_\,
            lcout => \nx.n1902\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9576_1_lut_LC_7_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30644\,
            lcout => \nx.n13425\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1144_3_lut_LC_7_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34482\,
            in2 => \N__31160\,
            in3 => \N__31131\,
            lcout => \nx.n1701\,
            ltout => \nx.n1701_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1211_3_lut_LC_7_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__35298\,
            in1 => \_gnd_net_\,
            in2 => \N__30867\,
            in3 => \N__35146\,
            lcout => \nx.n1800\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1212_3_lut_LC_7_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35357\,
            in2 => \N__35343\,
            in3 => \N__35147\,
            lcout => \nx.n1801\,
            ltout => \nx.n1801_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9_4_lut_adj_133_LC_7_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33016\,
            in1 => \N__35006\,
            in2 => \N__30864\,
            in3 => \N__34434\,
            lcout => \nx.n23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i3_3_lut_adj_82_LC_7_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34965\,
            in2 => \N__34912\,
            in3 => \N__35356\,
            lcout => \nx.n16_adj_672\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1149_3_lut_LC_7_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30891\,
            in2 => \N__30915\,
            in3 => \N__34481\,
            lcout => \nx.n1706\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_i7_LC_7_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000111100001000"
        )
    port map (
            in0 => \N__50076\,
            in1 => \N__49850\,
            in2 => \N__49601\,
            in3 => \N__37395\,
            lcout => neopxl_color_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48443\,
            ce => 'H',
            sr => \N__37371\
        );

    \nx.mod_5_i1084_3_lut_LC_7_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30855\,
            in2 => \N__33273\,
            in3 => \N__30844\,
            lcout => \nx.n1609\,
            ltout => \nx.n1609_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i4_3_lut_adj_89_LC_7_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31186\,
            in2 => \N__30804\,
            in3 => \N__30999\,
            lcout => \nx.n16_adj_646\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1151_3_lut_LC_7_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__30927\,
            in1 => \_gnd_net_\,
            in2 => \N__34500\,
            in3 => \N__30941\,
            lcout => \nx.n1708\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1145_3_lut_LC_7_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__31187\,
            in1 => \_gnd_net_\,
            in2 => \N__31173\,
            in3 => \N__34476\,
            lcout => \nx.n1702\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1077_3_lut_LC_7_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31041\,
            in2 => \N__33274\,
            in3 => \N__31031\,
            lcout => \nx.n1602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_2_lut_LC_7_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31004\,
            in2 => \_gnd_net_\,
            in3 => \N__30945\,
            lcout => \nx.n1677\,
            ltout => OPEN,
            carryin => \bfn_7_30_0_\,
            carryout => \nx.n10603\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_3_lut_LC_7_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30942\,
            in3 => \N__30921\,
            lcout => \nx.n1676\,
            ltout => OPEN,
            carryin => \nx.n10603\,
            carryout => \nx.n10604\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_4_lut_LC_7_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44932\,
            in2 => \N__34554\,
            in3 => \N__30918\,
            lcout => \nx.n1675\,
            ltout => OPEN,
            carryin => \nx.n10604\,
            carryout => \nx.n10605\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_5_lut_LC_7_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44935\,
            in2 => \N__30914\,
            in3 => \N__30882\,
            lcout => \nx.n1674\,
            ltout => OPEN,
            carryin => \nx.n10605\,
            carryout => \nx.n10606\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_6_lut_LC_7_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44933\,
            in2 => \N__33137\,
            in3 => \N__30879\,
            lcout => \nx.n1673\,
            ltout => OPEN,
            carryin => \nx.n10606\,
            carryout => \nx.n10607\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_7_lut_LC_7_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44936\,
            in2 => \N__33207\,
            in3 => \N__30870\,
            lcout => \nx.n1672\,
            ltout => OPEN,
            carryin => \nx.n10607\,
            carryout => \nx.n10608\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_8_lut_LC_7_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44934\,
            in2 => \N__33176\,
            in3 => \N__31194\,
            lcout => \nx.n1671\,
            ltout => OPEN,
            carryin => \nx.n10608\,
            carryout => \nx.n10609\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_9_lut_LC_7_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44937\,
            in2 => \N__31191\,
            in3 => \N__31164\,
            lcout => \nx.n1670\,
            ltout => OPEN,
            carryin => \nx.n10609\,
            carryout => \nx.n10610\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_10_lut_LC_7_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44518\,
            in2 => \N__31161\,
            in3 => \N__31122\,
            lcout => \nx.n1669\,
            ltout => OPEN,
            carryin => \bfn_7_31_0_\,
            carryout => \nx.n10611\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_11_lut_LC_7_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44520\,
            in2 => \N__33392\,
            in3 => \N__31119\,
            lcout => \nx.n1668\,
            ltout => OPEN,
            carryin => \nx.n10611\,
            carryout => \nx.n10612\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_12_lut_LC_7_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44519\,
            in2 => \N__31071\,
            in3 => \N__31116\,
            lcout => \nx.n1667\,
            ltout => OPEN,
            carryin => \nx.n10612\,
            carryout => \nx.n10613\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_13_lut_LC_7_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44521\,
            in2 => \N__31113\,
            in3 => \N__31092\,
            lcout => \nx.n1666\,
            ltout => OPEN,
            carryin => \nx.n10613\,
            carryout => \nx.n10614\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1138_14_lut_LC_7_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__44522\,
            in1 => \N__31088\,
            in2 => \N__34515\,
            in3 => \N__31074\,
            lcout => \nx.n1697\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1142_3_lut_LC_7_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31069\,
            in2 => \N__31050\,
            in3 => \N__34504\,
            lcout => \nx.n1699\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_210_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000101010"
        )
    port map (
            in0 => \N__47504\,
            in1 => \N__47995\,
            in2 => \N__37584\,
            in3 => \N__35502\,
            lcout => OPEN,
            ltout => \n7258_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i2_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__37583\,
            in1 => \N__31360\,
            in2 => \N__31257\,
            in3 => \N__46534\,
            lcout => pin_out_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48417\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_202_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101010"
        )
    port map (
            in0 => \N__47502\,
            in1 => \N__35471\,
            in2 => \N__42645\,
            in3 => \N__35504\,
            lcout => n7236,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_159_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001001100"
        )
    port map (
            in0 => \N__35525\,
            in1 => \N__47503\,
            in2 => \N__42702\,
            in3 => \N__37493\,
            lcout => OPEN,
            ltout => \n7270_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i5_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__35526\,
            in1 => \N__31214\,
            in2 => \N__31245\,
            in3 => \N__46519\,
            lcout => pin_out_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48412\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_206_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011001100"
        )
    port map (
            in0 => \N__35503\,
            in1 => \N__47501\,
            in2 => \N__42701\,
            in3 => \N__33098\,
            lcout => n7254,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_232_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__50328\,
            in1 => \_gnd_net_\,
            in2 => \N__49050\,
            in3 => \_gnd_net_\,
            lcout => n6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9305_3_lut_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49043\,
            in1 => \N__31213\,
            in2 => \_gnd_net_\,
            in3 => \N__35951\,
            lcout => OPEN,
            ltout => \n13152_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_pin_1__bdd_4_lut_9614_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__50562\,
            in1 => \N__50327\,
            in2 => \N__31197\,
            in3 => \N__31407\,
            lcout => OPEN,
            ltout => \n13462_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n13462_bdd_4_lut_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__31422\,
            in1 => \N__50563\,
            in2 => \N__31410\,
            in3 => \N__31341\,
            lcout => n13465,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9321_3_lut_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__40478\,
            in1 => \N__49044\,
            in2 => \_gnd_net_\,
            in3 => \N__40544\,
            lcout => n13168,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9306_3_lut_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49042\,
            in1 => \N__33502\,
            in2 => \_gnd_net_\,
            in3 => \N__33541\,
            lcout => n13153,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i3_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__33525\,
            in1 => \N__31388\,
            in2 => \N__37521\,
            in3 => \N__46530\,
            lcout => pin_out_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48413\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9300_3_lut_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31387\,
            in1 => \N__31361\,
            in2 => \_gnd_net_\,
            in3 => \N__49030\,
            lcout => n13147,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9320_3_lut_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40517\,
            in1 => \N__39221\,
            in2 => \_gnd_net_\,
            in3 => \N__49031\,
            lcout => OPEN,
            ltout => \n13167_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n13450_bdd_4_lut_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__31335\,
            in1 => \N__50568\,
            in2 => \N__31329\,
            in3 => \N__31326\,
            lcout => n13453,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1817_3_lut_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__33699\,
            in1 => \_gnd_net_\,
            in2 => \N__36194\,
            in3 => \N__33719\,
            lcout => \nx.n2694\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1820_3_lut_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36306\,
            in2 => \N__33765\,
            in3 => \N__36158\,
            lcout => \nx.n2697\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1827_3_lut_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37928\,
            in2 => \N__36191\,
            in3 => \N__33639\,
            lcout => \nx.n2704\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1818_3_lut_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36387\,
            in2 => \N__33735\,
            in3 => \N__36151\,
            lcout => \nx.n2695\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1821_3_lut_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36369\,
            in2 => \N__36193\,
            in3 => \N__33570\,
            lcout => \nx.n2698\,
            ltout => \nx.n2698_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i16_4_lut_adj_23_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31585\,
            in1 => \N__36080\,
            in2 => \N__31494\,
            in3 => \N__31474\,
            lcout => \nx.n39_adj_610\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1826_3_lut_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33627\,
            in2 => \N__36192\,
            in3 => \N__36339\,
            lcout => \nx.n2703\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1832_3_lut_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35907\,
            in1 => \N__33471\,
            in2 => \_gnd_net_\,
            in3 => \N__36144\,
            lcout => \nx.n2709\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1696_3_lut_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41226\,
            in1 => \N__41275\,
            in2 => \_gnd_net_\,
            in3 => \N__41593\,
            lcout => \nx.n2509\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1813_3_lut_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36411\,
            in2 => \N__36197\,
            in3 => \N__33660\,
            lcout => \nx.n2690\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1747_3_lut_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38295\,
            in2 => \N__39548\,
            in3 => \N__38271\,
            lcout => \nx.n2592\,
            ltout => \nx.n2592_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1814_3_lut_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__36166\,
            in1 => \N__33669\,
            in2 => \N__31425\,
            in3 => \_gnd_net_\,
            lcout => \nx.n2691\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1812_rep_23_3_lut_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36170\,
            in2 => \N__36438\,
            in3 => \N__33651\,
            lcout => \nx.n2689\,
            ltout => \nx.n2689_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_4_lut_adj_20_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31648\,
            in1 => \N__33884\,
            in2 => \N__31632\,
            in3 => \N__31610\,
            lcout => \nx.n36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1824_3_lut_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33600\,
            in2 => \N__36270\,
            in3 => \N__36171\,
            lcout => \nx.n2701\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1419_3_lut_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32013\,
            in2 => \N__32049\,
            in3 => \N__34160\,
            lcout => \nx.n2104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1420_3_lut_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__32061\,
            in1 => \_gnd_net_\,
            in2 => \N__34190\,
            in3 => \N__32097\,
            lcout => \nx.n2105\,
            ltout => \nx.n2105_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9_3_lut_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36737\,
            in2 => \N__31572\,
            in3 => \N__37316\,
            lcout => \nx.n26_adj_667\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1410_3_lut_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32196\,
            in2 => \N__32157\,
            in3 => \N__34159\,
            lcout => \nx.n2095\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1686_3_lut_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41385\,
            in2 => \N__43698\,
            in3 => \N__41612\,
            lcout => \nx.n2499\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1750_3_lut_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37972\,
            in2 => \N__37947\,
            in3 => \N__39544\,
            lcout => \nx.n2595\,
            ltout => \nx.n2595_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_4_lut_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36009\,
            in1 => \N__36713\,
            in2 => \N__31950\,
            in3 => \N__33680\,
            lcout => \nx.n35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1418_3_lut_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31965\,
            in2 => \N__32001\,
            in3 => \N__34164\,
            lcout => \nx.n2103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i10_4_lut_adj_68_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32332\,
            in1 => \N__32287\,
            in2 => \N__32247\,
            in3 => \N__34233\,
            lcout => OPEN,
            ltout => \nx.n26_adj_664_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_adj_71_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31947\,
            in1 => \N__33990\,
            in2 => \N__31935\,
            in3 => \N__31932\,
            lcout => \nx.n2027\,
            ltout => \nx.n2027_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1413_3_lut_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__32245\,
            in1 => \N__32214\,
            in2 => \N__31923\,
            in3 => \_gnd_net_\,
            lcout => \nx.n2098\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1414_3_lut_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32259\,
            in2 => \N__32292\,
            in3 => \N__34168\,
            lcout => \nx.n2099\,
            ltout => \nx.n2099_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i11_4_lut_adj_73_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37097\,
            in1 => \N__36976\,
            in2 => \N__31920\,
            in3 => \N__37027\,
            lcout => \nx.n28_adj_669\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i2030_3_lut_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31917\,
            in2 => \N__31890\,
            in3 => \N__31878\,
            lcout => \nx.n3003\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1415_3_lut_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__32333\,
            in1 => \_gnd_net_\,
            in2 => \N__34191\,
            in3 => \N__32304\,
            lcout => \nx.n2100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_2_lut_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34075\,
            in2 => \_gnd_net_\,
            in3 => \N__32109\,
            lcout => \nx.n2077\,
            ltout => OPEN,
            carryin => \bfn_9_23_0_\,
            carryout => \nx.n10657\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_3_lut_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34016\,
            in3 => \N__32106\,
            lcout => \nx.n2076\,
            ltout => OPEN,
            carryin => \nx.n10657\,
            carryout => \nx.n10658\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_4_lut_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44631\,
            in2 => \N__34290\,
            in3 => \N__32103\,
            lcout => \nx.n2075\,
            ltout => OPEN,
            carryin => \nx.n10658\,
            carryout => \nx.n10659\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_5_lut_LC_9_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44634\,
            in2 => \N__34691\,
            in3 => \N__32100\,
            lcout => \nx.n2074\,
            ltout => OPEN,
            carryin => \nx.n10659\,
            carryout => \nx.n10660\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_6_lut_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44632\,
            in2 => \N__32096\,
            in3 => \N__32052\,
            lcout => \nx.n2073\,
            ltout => OPEN,
            carryin => \nx.n10660\,
            carryout => \nx.n10661\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_7_lut_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44635\,
            in2 => \N__32048\,
            in3 => \N__32004\,
            lcout => \nx.n2072\,
            ltout => OPEN,
            carryin => \nx.n10661\,
            carryout => \nx.n10662\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_8_lut_LC_9_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44633\,
            in2 => \N__32000\,
            in3 => \N__31959\,
            lcout => \nx.n2071\,
            ltout => OPEN,
            carryin => \nx.n10662\,
            carryout => \nx.n10663\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_9_lut_LC_9_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44636\,
            in2 => \N__34041\,
            in3 => \N__31956\,
            lcout => \nx.n2070\,
            ltout => OPEN,
            carryin => \nx.n10663\,
            carryout => \nx.n10664\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_10_lut_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45134\,
            in2 => \N__34658\,
            in3 => \N__31953\,
            lcout => \nx.n2069\,
            ltout => OPEN,
            carryin => \bfn_9_24_0_\,
            carryout => \nx.n10665\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_11_lut_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45138\,
            in2 => \N__32334\,
            in3 => \N__32295\,
            lcout => \nx.n2068\,
            ltout => OPEN,
            carryin => \nx.n10665\,
            carryout => \nx.n10666\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_12_lut_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45135\,
            in2 => \N__32291\,
            in3 => \N__32250\,
            lcout => \nx.n2067\,
            ltout => OPEN,
            carryin => \nx.n10666\,
            carryout => \nx.n10667\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_13_lut_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45139\,
            in2 => \N__32246\,
            in3 => \N__32205\,
            lcout => \nx.n2066\,
            ltout => OPEN,
            carryin => \nx.n10667\,
            carryout => \nx.n10668\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_14_lut_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45136\,
            in2 => \N__34231\,
            in3 => \N__32202\,
            lcout => \nx.n2065\,
            ltout => OPEN,
            carryin => \nx.n10668\,
            carryout => \nx.n10669\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_15_lut_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45140\,
            in2 => \N__34388\,
            in3 => \N__32199\,
            lcout => \nx.n2064\,
            ltout => OPEN,
            carryin => \nx.n10669\,
            carryout => \nx.n10670\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_16_lut_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45137\,
            in2 => \N__32195\,
            in3 => \N__32142\,
            lcout => \nx.n2063\,
            ltout => OPEN,
            carryin => \nx.n10670\,
            carryout => \nx.n10671\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_17_lut_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45141\,
            in2 => \N__34346\,
            in3 => \N__32139\,
            lcout => \nx.n2062\,
            ltout => OPEN,
            carryin => \nx.n10671\,
            carryout => \nx.n10672\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1406_18_lut_LC_9_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__44630\,
            in1 => \N__34192\,
            in2 => \N__32136\,
            in3 => \N__32112\,
            lcout => \nx.n2093\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1280_3_lut_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__33075\,
            in1 => \_gnd_net_\,
            in2 => \N__35007\,
            in3 => \N__32903\,
            lcout => \nx.n1901\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9518_3_lut_LC_9_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34433\,
            in2 => \N__32553\,
            in3 => \N__32902\,
            lcout => \nx.n1905\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i10_4_lut_LC_9_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32422\,
            in1 => \N__32380\,
            in2 => \N__32791\,
            in3 => \N__32812\,
            lcout => \nx.n25_adj_606\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i8_4_lut_adj_155_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32978\,
            in1 => \N__34570\,
            in2 => \N__35049\,
            in3 => \N__32933\,
            lcout => \nx.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1279_3_lut_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33063\,
            in2 => \N__33039\,
            in3 => \N__32896\,
            lcout => \nx.n1900\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1210_3_lut_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35262\,
            in1 => \N__35283\,
            in2 => \_gnd_net_\,
            in3 => \N__35125\,
            lcout => \nx.n1799\,
            ltout => \nx.n1799_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1277_3_lut_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32967\,
            in2 => \N__32367\,
            in3 => \N__32898\,
            lcout => \nx.n1898\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1218_3_lut_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__35127\,
            in1 => \_gnd_net_\,
            in2 => \N__34869\,
            in3 => \N__34830\,
            lcout => \nx.n1807\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1208_3_lut_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35205\,
            in2 => \N__35169\,
            in3 => \N__35126\,
            lcout => \nx.n1797\,
            ltout => \nx.n1797_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1275_3_lut_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32897\,
            in2 => \N__32337\,
            in3 => \N__32922\,
            lcout => \nx.n1896\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i2_2_lut_adj_134_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32765\,
            in2 => \_gnd_net_\,
            in3 => \N__32721\,
            lcout => \nx.n30_adj_703\,
            ltout => OPEN,
            carryin => \bfn_9_27_0_\,
            carryout => \nx.n10628\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_3_lut_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32667\,
            in3 => \N__32631\,
            lcout => \nx.n1876\,
            ltout => OPEN,
            carryin => \nx.n10628\,
            carryout => \nx.n10629\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_4_lut_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44956\,
            in2 => \N__32628\,
            in3 => \N__32595\,
            lcout => \nx.n1875\,
            ltout => OPEN,
            carryin => \nx.n10629\,
            carryout => \nx.n10630\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_5_lut_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45296\,
            in2 => \N__32587\,
            in3 => \N__32556\,
            lcout => \nx.n1874\,
            ltout => OPEN,
            carryin => \nx.n10630\,
            carryout => \nx.n10631\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_6_lut_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44957\,
            in2 => \N__34432\,
            in3 => \N__32541\,
            lcout => \nx.n1873\,
            ltout => OPEN,
            carryin => \nx.n10631\,
            carryout => \nx.n10632\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_7_lut_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45297\,
            in2 => \N__32537\,
            in3 => \N__32493\,
            lcout => \nx.n1872\,
            ltout => OPEN,
            carryin => \nx.n10632\,
            carryout => \nx.n10633\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_8_lut_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44958\,
            in2 => \N__32490\,
            in3 => \N__32460\,
            lcout => \nx.n1871\,
            ltout => OPEN,
            carryin => \nx.n10633\,
            carryout => \nx.n10634\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_9_lut_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34612\,
            in2 => \N__45391\,
            in3 => \N__33078\,
            lcout => \nx.n1870\,
            ltout => OPEN,
            carryin => \nx.n10634\,
            carryout => \nx.n10635\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_10_lut_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44717\,
            in2 => \N__35005\,
            in3 => \N__33066\,
            lcout => \nx.n1869\,
            ltout => OPEN,
            carryin => \bfn_9_28_0_\,
            carryout => \nx.n10636\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_11_lut_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45096\,
            in2 => \N__33062\,
            in3 => \N__33027\,
            lcout => \nx.n1868\,
            ltout => OPEN,
            carryin => \nx.n10636\,
            carryout => \nx.n10637\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_12_lut_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44718\,
            in2 => \N__33024\,
            in3 => \N__32985\,
            lcout => \nx.n1867\,
            ltout => OPEN,
            carryin => \nx.n10637\,
            carryout => \nx.n10638\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_13_lut_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32982\,
            in2 => \N__45095\,
            in3 => \N__32958\,
            lcout => \nx.n1866\,
            ltout => OPEN,
            carryin => \nx.n10638\,
            carryout => \nx.n10639\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_14_lut_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44722\,
            in2 => \N__34577\,
            in3 => \N__32943\,
            lcout => \nx.n1865\,
            ltout => OPEN,
            carryin => \nx.n10639\,
            carryout => \nx.n10640\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_15_lut_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45097\,
            in2 => \N__32940\,
            in3 => \N__32913\,
            lcout => \nx.n1864\,
            ltout => OPEN,
            carryin => \nx.n10640\,
            carryout => \nx.n10641\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1272_16_lut_LC_9_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__45098\,
            in1 => \N__35045\,
            in2 => \N__32910\,
            in3 => \N__32823\,
            lcout => \nx.n1895\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1143_3_lut_LC_9_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33411\,
            in2 => \N__33399\,
            in3 => \N__34518\,
            lcout => \nx.n1700\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_i4_LC_9_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000111100001000"
        )
    port map (
            in0 => \N__49829\,
            in1 => \N__50078\,
            in2 => \N__49602\,
            in3 => \N__40864\,
            lcout => neopxl_color_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48446\,
            ce => 'H',
            sr => \N__40842\
        );

    \nx.mod_5_i1083_3_lut_LC_9_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33369\,
            in2 => \N__33339\,
            in3 => \N__33270\,
            lcout => \nx.n1608\,
            ltout => \nx.n1608_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6_2_lut_LC_9_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33324\,
            in3 => \N__33196\,
            lcout => \nx.n18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1080_3_lut_LC_9_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33312\,
            in2 => \N__33291\,
            in3 => \N__33271\,
            lcout => \nx.n1605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1146_3_lut_LC_9_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33177\,
            in2 => \N__33153\,
            in3 => \N__34511\,
            lcout => \nx.n1703\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1148_3_lut_LC_9_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__33138\,
            in1 => \_gnd_net_\,
            in2 => \N__34517\,
            in3 => \N__33120\,
            lcout => \nx.n1705\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_1096_i21_2_lut_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50554\,
            in2 => \_gnd_net_\,
            in3 => \N__50357\,
            lcout => n21,
            ltout => \n21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2930_3_lut_4_lut_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__40441\,
            in1 => \N__46965\,
            in2 => \N__33108\,
            in3 => \N__40352\,
            lcout => n6150,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i6_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__33477\,
            in1 => \N__46523\,
            in2 => \N__33548\,
            in3 => \N__33486\,
            lcout => pin_out_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48415\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_213_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000100"
        )
    port map (
            in0 => \N__37517\,
            in1 => \N__47495\,
            in2 => \N__35508\,
            in3 => \N__43293\,
            lcout => n7262,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i7_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__35445\,
            in1 => \N__35454\,
            in2 => \N__33509\,
            in3 => \N__46524\,
            lcout => pin_out_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48415\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__50126\,
            in1 => \N__40444\,
            in2 => \N__46959\,
            in3 => \N__46683\,
            lcout => n8_adj_780,
            ltout => \n8_adj_780_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_161_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000101010"
        )
    port map (
            in0 => \N__47496\,
            in1 => \N__37494\,
            in2 => \N__33480\,
            in3 => \N__47981\,
            lcout => n7274,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_2_lut_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35906\,
            in2 => \_gnd_net_\,
            in3 => \N__33462\,
            lcout => \nx.n2677\,
            ltout => OPEN,
            carryin => \bfn_10_17_0_\,
            carryout => \nx.n10768\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_3_lut_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35924\,
            in3 => \N__33444\,
            lcout => \nx.n2676\,
            ltout => OPEN,
            carryin => \nx.n10768\,
            carryout => \nx.n10769\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_4_lut_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45685\,
            in2 => \N__35825\,
            in3 => \N__33429\,
            lcout => \nx.n2675\,
            ltout => OPEN,
            carryin => \nx.n10769\,
            carryout => \nx.n10770\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_5_lut_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45688\,
            in2 => \N__39422\,
            in3 => \N__33414\,
            lcout => \nx.n2674\,
            ltout => OPEN,
            carryin => \nx.n10770\,
            carryout => \nx.n10771\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_6_lut_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45686\,
            in2 => \N__36240\,
            in3 => \N__33642\,
            lcout => \nx.n2673\,
            ltout => OPEN,
            carryin => \nx.n10771\,
            carryout => \nx.n10772\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_7_lut_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45689\,
            in2 => \N__37932\,
            in3 => \N__33630\,
            lcout => \nx.n2672\,
            ltout => OPEN,
            carryin => \nx.n10772\,
            carryout => \nx.n10773\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_8_lut_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45687\,
            in2 => \N__36335\,
            in3 => \N__33618\,
            lcout => \nx.n2671\,
            ltout => OPEN,
            carryin => \nx.n10773\,
            carryout => \nx.n10774\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_9_lut_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45690\,
            in2 => \N__36686\,
            in3 => \N__33603\,
            lcout => \nx.n2670\,
            ltout => OPEN,
            carryin => \nx.n10774\,
            carryout => \nx.n10775\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_10_lut_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45742\,
            in2 => \N__36263\,
            in3 => \N__33591\,
            lcout => \nx.n2669\,
            ltout => OPEN,
            carryin => \bfn_10_18_0_\,
            carryout => \nx.n10776\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_11_lut_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45746\,
            in2 => \N__37667\,
            in3 => \N__33576\,
            lcout => \nx.n2668\,
            ltout => OPEN,
            carryin => \nx.n10776\,
            carryout => \nx.n10777\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_12_lut_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45743\,
            in2 => \N__37617\,
            in3 => \N__33573\,
            lcout => \nx.n2667\,
            ltout => OPEN,
            carryin => \nx.n10777\,
            carryout => \nx.n10778\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_13_lut_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45747\,
            in2 => \N__36365\,
            in3 => \N__33564\,
            lcout => \nx.n2666\,
            ltout => OPEN,
            carryin => \nx.n10778\,
            carryout => \nx.n10779\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_14_lut_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45744\,
            in2 => \N__36301\,
            in3 => \N__33756\,
            lcout => \nx.n2665\,
            ltout => OPEN,
            carryin => \nx.n10779\,
            carryout => \nx.n10780\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_15_lut_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45748\,
            in2 => \N__37694\,
            in3 => \N__33738\,
            lcout => \nx.n2664\,
            ltout => OPEN,
            carryin => \nx.n10780\,
            carryout => \nx.n10781\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_16_lut_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45745\,
            in2 => \N__36386\,
            in3 => \N__33726\,
            lcout => \nx.n2663\,
            ltout => OPEN,
            carryin => \nx.n10781\,
            carryout => \nx.n10782\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_17_lut_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45749\,
            in2 => \N__33723\,
            in3 => \N__33693\,
            lcout => \nx.n2662\,
            ltout => OPEN,
            carryin => \nx.n10782\,
            carryout => \nx.n10783\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_18_lut_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45733\,
            in2 => \N__36008\,
            in3 => \N__33690\,
            lcout => \nx.n2661\,
            ltout => OPEN,
            carryin => \bfn_10_19_0_\,
            carryout => \nx.n10784\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_19_lut_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36714\,
            in2 => \N__45765\,
            in3 => \N__33687\,
            lcout => \nx.n2660\,
            ltout => OPEN,
            carryin => \nx.n10784\,
            carryout => \nx.n10785\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_20_lut_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45737\,
            in2 => \N__33684\,
            in3 => \N__33663\,
            lcout => \nx.n2659\,
            ltout => OPEN,
            carryin => \nx.n10785\,
            carryout => \nx.n10786\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_21_lut_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45739\,
            in2 => \N__36410\,
            in3 => \N__33654\,
            lcout => \nx.n2658\,
            ltout => OPEN,
            carryin => \nx.n10786\,
            carryout => \nx.n10787\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_22_lut_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45738\,
            in2 => \N__36434\,
            in3 => \N__33645\,
            lcout => \nx.n2657\,
            ltout => OPEN,
            carryin => \nx.n10787\,
            carryout => \nx.n10788\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_23_lut_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45740\,
            in2 => \N__36657\,
            in3 => \N__33921\,
            lcout => \nx.n2656\,
            ltout => OPEN,
            carryin => \nx.n10788\,
            carryout => \nx.n10789\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1808_24_lut_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__45741\,
            in1 => \N__38169\,
            in2 => \N__36198\,
            in3 => \N__33918\,
            lcout => \nx.n2687\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1815_3_lut_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36712\,
            in2 => \N__33915\,
            in3 => \N__36159\,
            lcout => \nx.n2692\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i12_4_lut_adj_17_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36427\,
            in1 => \N__36403\,
            in2 => \N__36656\,
            in3 => \N__38168\,
            lcout => OPEN,
            ltout => \nx.n34_adj_603_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i17_3_lut_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37615\,
            in2 => \N__33873\,
            in3 => \N__36676\,
            lcout => OPEN,
            ltout => \nx.n39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i21_4_lut_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36312\,
            in1 => \N__36276\,
            in2 => \N__33870\,
            in3 => \N__35835\,
            lcout => \nx.n2621\,
            ltout => \nx.n2621_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1816_3_lut_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__36004\,
            in1 => \_gnd_net_\,
            in2 => \N__33867\,
            in3 => \N__33864\,
            lcout => \nx.n2693\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1822_3_lut_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__37616\,
            in1 => \_gnd_net_\,
            in2 => \N__36196\,
            in3 => \N__33822\,
            lcout => \nx.n2699\,
            ltout => \nx.n2699_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i18_4_lut_adj_22_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33779\,
            in1 => \N__36625\,
            in2 => \N__33768\,
            in3 => \N__33984\,
            lcout => \nx.n41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1811_3_lut_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__36652\,
            in1 => \_gnd_net_\,
            in2 => \N__36195\,
            in3 => \N__33966\,
            lcout => \nx.n2688\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1683_3_lut_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__41316\,
            in1 => \_gnd_net_\,
            in2 => \N__41661\,
            in3 => \N__43200\,
            lcout => \nx.n2496\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i11_4_lut_adj_59_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41722\,
            in1 => \N__44010\,
            in2 => \N__41478\,
            in3 => \N__41764\,
            lcout => OPEN,
            ltout => \nx.n31_adj_655_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i16_4_lut_adj_60_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41804\,
            in1 => \N__41843\,
            in2 => \N__33960\,
            in3 => \N__33957\,
            lcout => OPEN,
            ltout => \nx.n36_adj_656_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i19_4_lut_adj_65_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43641\,
            in1 => \N__39702\,
            in2 => \N__33942\,
            in3 => \N__33939\,
            lcout => \nx.n2423\,
            ltout => \nx.n2423_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1677_3_lut_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41477\,
            in2 => \N__33927\,
            in3 => \N__41685\,
            lcout => \nx.n2490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1678_3_lut_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__41723\,
            in1 => \_gnd_net_\,
            in2 => \N__41703\,
            in3 => \N__41636\,
            lcout => \nx.n2491\,
            ltout => \nx.n2491_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i12_4_lut_adj_56_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38248\,
            in1 => \N__38315\,
            in2 => \N__33924\,
            in3 => \N__38284\,
            lcout => \nx.n33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1679_3_lut_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41765\,
            in2 => \N__41748\,
            in3 => \N__41635\,
            lcout => \nx.n2492\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1611_3_lut_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45828\,
            in2 => \N__45848\,
            in3 => \N__44122\,
            lcout => \nx.n2392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1612_3_lut_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45890\,
            in2 => \N__44129\,
            in3 => \N__45870\,
            lcout => \nx.n2393\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1613_3_lut_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45938\,
            in2 => \N__45918\,
            in3 => \N__44118\,
            lcout => \nx.n2394\,
            ltout => \nx.n2394_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1680_3_lut_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41611\,
            in2 => \N__34113\,
            in3 => \N__41790\,
            lcout => \nx.n2493\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1424_3_lut_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34110\,
            in1 => \N__34083\,
            in2 => \_gnd_net_\,
            in3 => \N__34189\,
            lcout => \nx.n2109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1417_3_lut_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__34040\,
            in1 => \_gnd_net_\,
            in2 => \N__34197\,
            in3 => \N__34104\,
            lcout => \nx.n2102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1416_3_lut_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__34659\,
            in1 => \_gnd_net_\,
            in2 => \N__34098\,
            in3 => \N__34183\,
            lcout => \nx.n2101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1423_3_lut_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34089\,
            in2 => \N__34195\,
            in3 => \N__34015\,
            lcout => \nx.n2108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i11_4_lut_adj_69_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__34076\,
            in1 => \N__34039\,
            in2 => \N__34017\,
            in3 => \N__34626\,
            lcout => \nx.n27_adj_665\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1421_3_lut_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34404\,
            in2 => \N__34196\,
            in3 => \N__34687\,
            lcout => \nx.n2106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1411_3_lut_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34398\,
            in2 => \N__34392\,
            in3 => \N__34184\,
            lcout => \nx.n2096\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1409_3_lut_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34356\,
            in2 => \N__34350\,
            in3 => \N__34185\,
            lcout => \nx.n2094\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_4_lut_adj_72_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__37081\,
            in1 => \N__36910\,
            in2 => \N__36873\,
            in3 => \N__34311\,
            lcout => OPEN,
            ltout => \nx.n30_adj_668_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i16_4_lut_adj_76_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34245\,
            in1 => \N__34698\,
            in2 => \N__34302\,
            in3 => \N__34299\,
            lcout => \nx.n2126\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1422_3_lut_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34289\,
            in2 => \N__34257\,
            in3 => \N__34193\,
            lcout => \nx.n2107\,
            ltout => \nx.n2107_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i12_4_lut_adj_74_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36826\,
            in1 => \N__36790\,
            in2 => \N__34248\,
            in3 => \N__37294\,
            lcout => \nx.n29_adj_670\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1412_3_lut_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34239\,
            in2 => \N__34232\,
            in3 => \N__34194\,
            lcout => \nx.n2097\,
            ltout => \nx.n2097_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i10_4_lut_adj_75_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37060\,
            in1 => \N__36940\,
            in2 => \N__34701\,
            in3 => \N__37270\,
            lcout => \nx.n27_adj_671\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9587_1_lut_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37193\,
            lcout => \nx.n13436\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6_2_lut_adj_66_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34692\,
            in3 => \N__34645\,
            lcout => \nx.n22_adj_662\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1214_3_lut_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35439\,
            in2 => \N__35128\,
            in3 => \N__35403\,
            lcout => \nx.n1803\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9_4_lut_adj_83_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34787\,
            in1 => \N__34741\,
            in2 => \N__34818\,
            in3 => \N__35318\,
            lcout => OPEN,
            ltout => \nx.n22_adj_673_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i11_4_lut_adj_99_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35278\,
            in1 => \N__35242\,
            in2 => \N__34593\,
            in3 => \N__34590\,
            lcout => \nx.n24_adj_685\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1209_3_lut_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35217\,
            in2 => \N__35249\,
            in3 => \N__35108\,
            lcout => \nx.n1798\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1150_rep_76_3_lut_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34550\,
            in2 => \N__34533\,
            in3 => \N__34516\,
            lcout => \nx.n1707\,
            ltout => \nx.n1707_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9517_3_lut_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34803\,
            in2 => \N__34437\,
            in3 => \N__35107\,
            lcout => \nx.n1806\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i12_4_lut_adj_110_LC_10_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35393\,
            in1 => \N__34868\,
            in2 => \N__35031\,
            in3 => \N__35016\,
            lcout => \nx.n1730\,
            ltout => \nx.n1730_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1213_3_lut_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__35373\,
            in1 => \_gnd_net_\,
            in2 => \N__35010\,
            in3 => \N__35394\,
            lcout => \nx.n1802\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_2_lut_LC_10_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34975\,
            in2 => \_gnd_net_\,
            in3 => \N__34920\,
            lcout => \nx.n1777\,
            ltout => OPEN,
            carryin => \bfn_10_28_0_\,
            carryout => \nx.n10615\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_3_lut_LC_10_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34917\,
            in3 => \N__34872\,
            lcout => \nx.n1776\,
            ltout => OPEN,
            carryin => \nx.n10615\,
            carryout => \nx.n10616\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_4_lut_LC_10_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44596\,
            in2 => \N__34867\,
            in3 => \N__34821\,
            lcout => \nx.n1775\,
            ltout => OPEN,
            carryin => \nx.n10616\,
            carryout => \nx.n10617\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_5_lut_LC_10_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34814\,
            in2 => \N__44955\,
            in3 => \N__34797\,
            lcout => \nx.n1774\,
            ltout => OPEN,
            carryin => \nx.n10617\,
            carryout => \nx.n10618\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_6_lut_LC_10_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44600\,
            in2 => \N__34794\,
            in3 => \N__34752\,
            lcout => \nx.n1773\,
            ltout => OPEN,
            carryin => \nx.n10618\,
            carryout => \nx.n10619\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_7_lut_LC_10_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44862\,
            in2 => \N__34742\,
            in3 => \N__34704\,
            lcout => \nx.n1772\,
            ltout => OPEN,
            carryin => \nx.n10619\,
            carryout => \nx.n10620\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_8_lut_LC_10_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44601\,
            in2 => \N__35438\,
            in3 => \N__35397\,
            lcout => \nx.n1771\,
            ltout => OPEN,
            carryin => \nx.n10620\,
            carryout => \nx.n10621\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_9_lut_LC_10_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44863\,
            in2 => \N__35392\,
            in3 => \N__35367\,
            lcout => \nx.n1770\,
            ltout => OPEN,
            carryin => \nx.n10621\,
            carryout => \nx.n10622\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_10_lut_LC_10_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44433\,
            in2 => \N__35364\,
            in3 => \N__35325\,
            lcout => \nx.n1769\,
            ltout => OPEN,
            carryin => \bfn_10_29_0_\,
            carryout => \nx.n10623\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_11_lut_LC_10_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44436\,
            in2 => \N__35322\,
            in3 => \N__35286\,
            lcout => \nx.n1768\,
            ltout => OPEN,
            carryin => \nx.n10623\,
            carryout => \nx.n10624\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_12_lut_LC_10_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35279\,
            in2 => \N__44716\,
            in3 => \N__35253\,
            lcout => \nx.n1767\,
            ltout => OPEN,
            carryin => \nx.n10624\,
            carryout => \nx.n10625\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_13_lut_LC_10_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44440\,
            in2 => \N__35250\,
            in3 => \N__35208\,
            lcout => \nx.n1766\,
            ltout => OPEN,
            carryin => \nx.n10625\,
            carryout => \nx.n10626\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_14_lut_LC_10_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44434\,
            in2 => \N__35204\,
            in3 => \N__35154\,
            lcout => \nx.n1765\,
            ltout => OPEN,
            carryin => \nx.n10626\,
            carryout => \nx.n10627\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1205_15_lut_LC_10_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__44435\,
            in1 => \N__35145\,
            in2 => \N__35073\,
            in3 => \N__35052\,
            lcout => \nx.n1796\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_enable__i1_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__50067\,
            in1 => \N__49838\,
            in2 => \_gnd_net_\,
            in3 => \N__49570\,
            lcout => pin_oe_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48421\,
            ce => \N__37338\,
            sr => \_gnd_net_\
        );

    \i2938_3_lut_4_lut_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__38906\,
            in1 => \N__40401\,
            in2 => \N__49048\,
            in3 => \N__46964\,
            lcout => n6158,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_290_i8_2_lut_3_lut_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__48701\,
            in1 => \_gnd_net_\,
            in2 => \N__50778\,
            in3 => \N__50555\,
            lcout => n8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_1101_i22_2_lut_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48700\,
            in2 => \_gnd_net_\,
            in3 => \N__50773\,
            lcout => n22_adj_740,
            ltout => \n22_adj_740_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2691_3_lut_4_lut_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__46722\,
            in1 => \N__46963\,
            in2 => \N__35475\,
            in3 => \N__46642\,
            lcout => n5907,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2936_3_lut_4_lut_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__46923\,
            in1 => \N__40397\,
            in2 => \N__49049\,
            in3 => \N__38910\,
            lcout => n6156,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i21_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__39072\,
            in1 => \N__39084\,
            in2 => \N__42899\,
            in3 => \N__46529\,
            lcout => pin_out_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48418\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2942_3_lut_4_lut_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__40443\,
            in1 => \N__50127\,
            in2 => \N__46958\,
            in3 => \N__40361\,
            lcout => n6162,
            ltout => \n6162_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_163_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000000"
        )
    port map (
            in0 => \N__43294\,
            in1 => \N__37480\,
            in2 => \N__35448\,
            in3 => \N__47497\,
            lcout => n7278,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000101010"
        )
    port map (
            in0 => \N__47422\,
            in1 => \N__42640\,
            in2 => \N__35982\,
            in3 => \N__37481\,
            lcout => OPEN,
            ltout => \n7266_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i4_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__35981\,
            in1 => \N__35947\,
            in2 => \N__35967\,
            in3 => \N__46528\,
            lcout => pin_out_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_751_i10_2_lut_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50730\,
            in2 => \_gnd_net_\,
            in3 => \N__50564\,
            lcout => n10_adj_736,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1764_3_lut_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37833\,
            in1 => \N__37892\,
            in2 => \_gnd_net_\,
            in3 => \N__39509\,
            lcout => \nx.n2609\,
            ltout => \nx.n2609_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6_3_lut_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35899\,
            in2 => \N__35853\,
            in3 => \N__37681\,
            lcout => OPEN,
            ltout => \nx.n28_adj_599_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i18_4_lut_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35821\,
            in1 => \N__37660\,
            in2 => \N__35850\,
            in3 => \N__35847\,
            lcout => \nx.n40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1753_3_lut_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__38034\,
            in1 => \_gnd_net_\,
            in2 => \N__38070\,
            in3 => \N__39517\,
            lcout => \nx.n2598\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1763_3_lut_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37788\,
            in2 => \N__39538\,
            in3 => \N__37821\,
            lcout => \nx.n2608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9530_3_lut_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37754\,
            in2 => \N__37725\,
            in3 => \N__39513\,
            lcout => \nx.n2604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9520_3_lut_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__39597\,
            in1 => \_gnd_net_\,
            in2 => \N__39539\,
            in3 => \N__38085\,
            lcout => \nx.n2599\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1751_3_lut_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37989\,
            in2 => \N__39537\,
            in3 => \N__38003\,
            lcout => \nx.n2596\,
            ltout => \nx.n2596_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37921\,
            in1 => \N__36361\,
            in2 => \N__36342\,
            in3 => \N__36331\,
            lcout => \nx.n37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i16_4_lut_adj_18_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36259\,
            in1 => \N__39412\,
            in2 => \N__36302\,
            in3 => \N__36236\,
            lcout => \nx.n38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9526_3_lut_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38142\,
            in2 => \N__39357\,
            in3 => \N__39503\,
            lcout => \nx.n2602\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1761_3_lut_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37773\,
            in2 => \N__39536\,
            in3 => \N__39637\,
            lcout => \nx.n2606\,
            ltout => \nx.n2606_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1828_3_lut_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36222\,
            in2 => \N__36213\,
            in3 => \N__36172\,
            lcout => \nx.n2705\,
            ltout => \nx.n2705_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1895_3_lut_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36060\,
            in2 => \N__36051\,
            in3 => \N__36586\,
            lcout => \nx.n2804\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1749_3_lut_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38328\,
            in2 => \N__39387\,
            in3 => \N__39499\,
            lcout => \nx.n2594\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9536_3_lut_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41061\,
            in2 => \N__41031\,
            in3 => \N__41600\,
            lcout => \nx.n2504\,
            ltout => \nx.n2504_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9528_3_lut_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37710\,
            in2 => \N__36690\,
            in3 => \N__39518\,
            lcout => \nx.n2603\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_i6_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010101000000"
        )
    port map (
            in0 => \N__49581\,
            in1 => \N__50034\,
            in2 => \N__49828\,
            in3 => \N__40746\,
            lcout => neopxl_color_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48422\,
            ce => 'H',
            sr => \N__40719\
        );

    \nx.mod_5_i1744_3_lut_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39685\,
            in2 => \N__38187\,
            in3 => \N__39523\,
            lcout => \nx.n2589\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1878_3_lut_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36629\,
            in2 => \N__36609\,
            in3 => \N__36477\,
            lcout => \nx.n2787\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1745_3_lut_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38213\,
            in2 => \N__39540\,
            in3 => \N__38199\,
            lcout => \nx.n2590\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1746_3_lut_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38232\,
            in1 => \N__38252\,
            in2 => \_gnd_net_\,
            in3 => \N__39519\,
            lcout => \nx.n2591\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_i5_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001000100010"
        )
    port map (
            in0 => \N__39777\,
            in1 => \N__49580\,
            in2 => \N__50066\,
            in3 => \N__49818\,
            lcout => neopxl_color_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48425\,
            ce => 'H',
            sr => \N__39744\
        );

    \nx.mod_5_i1547_3_lut_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__40228\,
            in1 => \_gnd_net_\,
            in2 => \N__41988\,
            in3 => \N__40206\,
            lcout => \nx.n2296\,
            ltout => \nx.n2296_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1614_3_lut_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__45960\,
            in1 => \_gnd_net_\,
            in2 => \N__36723\,
            in3 => \N__44127\,
            lcout => \nx.n2395\,
            ltout => \nx.n2395_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1681_3_lut_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41826\,
            in2 => \N__36720\,
            in3 => \N__41598\,
            lcout => \nx.n2494\,
            ltout => \nx.n2494_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1748_3_lut_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38304\,
            in2 => \N__36717\,
            in3 => \N__39526\,
            lcout => \nx.n2593\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9542_3_lut_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41442\,
            in2 => \N__43626\,
            in3 => \N__41599\,
            lcout => \nx.n2501\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9529_3_lut_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__41076\,
            in1 => \_gnd_net_\,
            in2 => \N__41631\,
            in3 => \N__43599\,
            lcout => \nx.n2505\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i3_2_lut_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40230\,
            in3 => \N__40189\,
            lcout => \nx.n21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1694_3_lut_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41124\,
            in2 => \N__41154\,
            in3 => \N__41594\,
            lcout => \nx.n2507\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1545_3_lut_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40151\,
            in2 => \N__40125\,
            in3 => \N__41948\,
            lcout => \nx.n2294\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1544_3_lut_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40077\,
            in2 => \N__40106\,
            in3 => \N__41949\,
            lcout => \nx.n2293\,
            ltout => \nx.n2293_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i11_4_lut_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45934\,
            in1 => \N__45886\,
            in2 => \N__36921\,
            in3 => \N__45971\,
            lcout => \nx.n30_adj_640\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1546_3_lut_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40190\,
            in2 => \N__41974\,
            in3 => \N__40167\,
            lcout => \nx.n2295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_2_lut_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__36918\,
            in1 => \N__36917\,
            in2 => \N__36848\,
            in3 => \N__36876\,
            lcout => \nx.n2209\,
            ltout => OPEN,
            carryin => \bfn_11_23_0_\,
            carryout => \nx.n10673\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_3_lut_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__36869\,
            in1 => \N__36868\,
            in2 => \N__36849\,
            in3 => \N__36831\,
            lcout => \nx.n2208\,
            ltout => OPEN,
            carryin => \nx.n10673\,
            carryout => \nx.n10674\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_4_lut_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__36828\,
            in1 => \N__36827\,
            in2 => \N__37242\,
            in3 => \N__36810\,
            lcout => \nx.n2207\,
            ltout => OPEN,
            carryin => \nx.n10674\,
            carryout => \nx.n10675\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_5_lut_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__36807\,
            in1 => \N__36806\,
            in2 => \N__37245\,
            in3 => \N__36795\,
            lcout => \nx.n2206\,
            ltout => OPEN,
            carryin => \nx.n10675\,
            carryout => \nx.n10676\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_6_lut_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__36792\,
            in1 => \N__36791\,
            in2 => \N__37243\,
            in3 => \N__36774\,
            lcout => \nx.n2205\,
            ltout => OPEN,
            carryin => \nx.n10676\,
            carryout => \nx.n10677\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_7_lut_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__36771\,
            in1 => \N__36770\,
            in2 => \N__37246\,
            in3 => \N__36753\,
            lcout => \nx.n2204\,
            ltout => OPEN,
            carryin => \nx.n10677\,
            carryout => \nx.n10678\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_8_lut_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__36750\,
            in1 => \N__36749\,
            in2 => \N__37244\,
            in3 => \N__36726\,
            lcout => \nx.n2203\,
            ltout => OPEN,
            carryin => \nx.n10678\,
            carryout => \nx.n10679\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_9_lut_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__37110\,
            in1 => \N__37109\,
            in2 => \N__37247\,
            in3 => \N__37086\,
            lcout => \nx.n2202\,
            ltout => OPEN,
            carryin => \nx.n10679\,
            carryout => \nx.n10680\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_10_lut_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__37083\,
            in1 => \N__37082\,
            in2 => \N__37248\,
            in3 => \N__37065\,
            lcout => \nx.n2201\,
            ltout => OPEN,
            carryin => \bfn_11_24_0_\,
            carryout => \nx.n10681\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_11_lut_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__37062\,
            in1 => \N__37061\,
            in2 => \N__37252\,
            in3 => \N__37044\,
            lcout => \nx.n2200\,
            ltout => OPEN,
            carryin => \nx.n10681\,
            carryout => \nx.n10682\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_12_lut_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__37041\,
            in1 => \N__37040\,
            in2 => \N__37249\,
            in3 => \N__37014\,
            lcout => \nx.n2199\,
            ltout => OPEN,
            carryin => \nx.n10682\,
            carryout => \nx.n10683\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_13_lut_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__37011\,
            in1 => \N__37010\,
            in2 => \N__37253\,
            in3 => \N__36993\,
            lcout => \nx.n2198\,
            ltout => OPEN,
            carryin => \nx.n10683\,
            carryout => \nx.n10684\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_14_lut_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__36990\,
            in1 => \N__36989\,
            in2 => \N__37250\,
            in3 => \N__36963\,
            lcout => \nx.n2197\,
            ltout => OPEN,
            carryin => \nx.n10684\,
            carryout => \nx.n10685\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_15_lut_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__36960\,
            in1 => \N__36956\,
            in2 => \N__37254\,
            in3 => \N__36945\,
            lcout => \nx.n2196\,
            ltout => OPEN,
            carryin => \nx.n10685\,
            carryout => \nx.n10686\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_16_lut_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__36942\,
            in1 => \N__36941\,
            in2 => \N__37251\,
            in3 => \N__36924\,
            lcout => \nx.n2195\,
            ltout => OPEN,
            carryin => \nx.n10686\,
            carryout => \nx.n10687\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_17_lut_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__37329\,
            in1 => \N__37328\,
            in2 => \N__37255\,
            in3 => \N__37305\,
            lcout => \nx.n2194\,
            ltout => OPEN,
            carryin => \nx.n10687\,
            carryout => \nx.n10688\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_18_lut_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__37302\,
            in1 => \N__37301\,
            in2 => \N__37256\,
            in3 => \N__37281\,
            lcout => \nx.n2193\,
            ltout => OPEN,
            carryin => \bfn_11_25_0_\,
            carryout => \nx.n10689\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1473_19_lut_LC_11_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__37277\,
            in1 => \N__37278\,
            in2 => \N__37257\,
            in3 => \N__37137\,
            lcout => \nx.n2192\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7849_4_lut_LC_11_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__37347\,
            in1 => \N__38631\,
            in2 => \N__37134\,
            in3 => \N__38889\,
            lcout => n11612,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_adj_229_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38673\,
            in1 => \N__37125\,
            in2 => \N__38715\,
            in3 => \N__37443\,
            lcout => n12171,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_11_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__38691\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38652\,
            lcout => n6_adj_761,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_LC_11_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38378\,
            in1 => \N__38552\,
            in2 => \N__38397\,
            in3 => \N__38537\,
            lcout => OPEN,
            ltout => \n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_LC_11_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38567\,
            in1 => \N__38363\,
            in2 => \N__37119\,
            in3 => \N__37116\,
            lcout => n12091,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_3_lut_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__38597\,
            in1 => \N__38582\,
            in2 => \_gnd_net_\,
            in3 => \N__38612\,
            lcout => n14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1390_4_lut_LC_11_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__38504\,
            in1 => \N__37452\,
            in2 => \N__38523\,
            in3 => \N__38489\,
            lcout => OPEN,
            ltout => \n24_adj_720_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_226_LC_11_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__38744\,
            in1 => \N__38759\,
            in2 => \N__37446\,
            in3 => \N__38729\,
            lcout => n11898,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_adj_228_LC_11_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38792\,
            in1 => \N__39041\,
            in2 => \N__38856\,
            in3 => \N__38837\,
            lcout => n17_adj_765,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_195_LC_11_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__37416\,
            in1 => \N__50068\,
            in2 => \_gnd_net_\,
            in3 => \N__49834\,
            lcout => n22_adj_724,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_227_LC_11_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39011\,
            in1 => \N__38807\,
            in2 => \N__38778\,
            in3 => \N__39026\,
            lcout => OPEN,
            ltout => \n16_adj_764_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9_4_lut_LC_11_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38870\,
            in1 => \N__37356\,
            in2 => \N__37350\,
            in3 => \N__38822\,
            lcout => n10978,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_11_32_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_224_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000010"
        )
    port map (
            in0 => \N__50044\,
            in1 => \N__49830\,
            in2 => \N__49588\,
            in3 => \N__37461\,
            lcout => n36,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9315_3_lut_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37544\,
            in1 => \N__38926\,
            in2 => \_gnd_net_\,
            in3 => \N__49033\,
            lcout => n13162,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9564_2_lut_3_lut_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__47163\,
            in1 => \N__48133\,
            in2 => \_gnd_net_\,
            in3 => \N__47230\,
            lcout => \state_7_N_167_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_188_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47231\,
            in1 => \N__47164\,
            in2 => \N__48147\,
            in3 => \N__49032\,
            lcout => n7166,
            ltout => \n7166_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2932_3_lut_4_lut_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__40664\,
            in1 => \N__40442\,
            in2 => \N__37587\,
            in3 => \N__46944\,
            lcout => n6152,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_282_i8_2_lut_3_lut_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__48699\,
            in1 => \N__50777\,
            in2 => \_gnd_net_\,
            in3 => \N__50573\,
            lcout => n8_adj_751,
            ltout => \n8_adj_751_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_171_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101010"
        )
    port map (
            in0 => \N__47476\,
            in1 => \N__43295\,
            in2 => \N__37566\,
            in3 => \N__39062\,
            lcout => OPEN,
            ltout => \n7294_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i11_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__39063\,
            in1 => \N__37540\,
            in2 => \N__37563\,
            in3 => \N__46518\,
            lcout => pin_out_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48420\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2934_3_lut_4_lut_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__40334\,
            in1 => \N__40657\,
            in2 => \N__40448\,
            in3 => \N__46915\,
            lcout => n6154,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_284_i8_2_lut_3_lut_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__48698\,
            in1 => \N__50772\,
            in2 => \_gnd_net_\,
            in3 => \N__50534\,
            lcout => n8_adj_744,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9272_2_lut_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48482\,
            in2 => \_gnd_net_\,
            in3 => \N__48527\,
            lcout => OPEN,
            ltout => \n13048_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9443_4_lut_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__39053\,
            in1 => \N__47654\,
            in2 => \N__37464\,
            in3 => \N__48572\,
            lcout => n13264,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9434_3_lut_4_lut_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__48573\,
            in1 => \N__39054\,
            in2 => \N__48492\,
            in3 => \N__48534\,
            lcout => n13273,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__50007\,
            in1 => \N__49771\,
            in2 => \_gnd_net_\,
            in3 => \N__49510\,
            lcout => n7231,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1752_3_lut_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39729\,
            in2 => \N__38022\,
            in3 => \N__39525\,
            lcout => \nx.n2597\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9524_3_lut_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38133\,
            in2 => \N__39324\,
            in3 => \N__39524\,
            lcout => \nx.n2601\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1684_3_lut_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43233\,
            in2 => \N__41334\,
            in3 => \N__41660\,
            lcout => \nx.n2497\,
            ltout => \nx.n2497_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i5_3_lut_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37896\,
            in2 => \N__37641\,
            in3 => \N__37820\,
            lcout => OPEN,
            ltout => \nx.n26_adj_611_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i17_4_lut_adj_24_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37974\,
            in1 => \N__39376\,
            in2 => \N__37638\,
            in3 => \N__37635\,
            lcout => OPEN,
            ltout => \nx.n38_adj_612_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i20_4_lut_adj_48_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37902\,
            in1 => \N__39606\,
            in2 => \N__37623\,
            in3 => \N__39330\,
            lcout => \nx.n2522\,
            ltout => \nx.n2522_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9522_3_lut_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__38121\,
            in1 => \N__38097\,
            in2 => \N__37620\,
            in3 => \_gnd_net_\,
            lcout => \nx.n2600\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9532_3_lut_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37764\,
            in2 => \N__39273\,
            in3 => \N__39508\,
            lcout => \nx.n2605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i14_4_lut_adj_46_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38120\,
            in1 => \N__38065\,
            in2 => \N__37755\,
            in3 => \N__39724\,
            lcout => \nx.n35_adj_639\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_2_lut_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37891\,
            in2 => \_gnd_net_\,
            in3 => \N__37824\,
            lcout => \nx.n2577\,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => \nx.n10747\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_3_lut_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37819\,
            in3 => \N__37779\,
            lcout => \nx.n2576\,
            ltout => OPEN,
            carryin => \nx.n10747\,
            carryout => \nx.n10748\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_4_lut_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45450\,
            in2 => \N__39296\,
            in3 => \N__37776\,
            lcout => \nx.n2575\,
            ltout => OPEN,
            carryin => \nx.n10748\,
            carryout => \nx.n10749\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_5_lut_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45453\,
            in2 => \N__39638\,
            in3 => \N__37767\,
            lcout => \nx.n2574\,
            ltout => OPEN,
            carryin => \nx.n10749\,
            carryout => \nx.n10750\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_6_lut_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45451\,
            in2 => \N__39272\,
            in3 => \N__37758\,
            lcout => \nx.n2573\,
            ltout => OPEN,
            carryin => \nx.n10750\,
            carryout => \nx.n10751\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_7_lut_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45454\,
            in2 => \N__37744\,
            in3 => \N__37713\,
            lcout => \nx.n2572\,
            ltout => OPEN,
            carryin => \nx.n10751\,
            carryout => \nx.n10752\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_8_lut_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45452\,
            in2 => \N__39659\,
            in3 => \N__38145\,
            lcout => \nx.n2571\,
            ltout => OPEN,
            carryin => \nx.n10752\,
            carryout => \nx.n10753\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_9_lut_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45455\,
            in2 => \N__39350\,
            in3 => \N__38136\,
            lcout => \nx.n2570\,
            ltout => OPEN,
            carryin => \nx.n10753\,
            carryout => \nx.n10754\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_10_lut_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45440\,
            in2 => \N__39320\,
            in3 => \N__38124\,
            lcout => \nx.n2569\,
            ltout => OPEN,
            carryin => \bfn_12_21_0_\,
            carryout => \nx.n10755\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_11_lut_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45025\,
            in2 => \N__38114\,
            in3 => \N__38088\,
            lcout => \nx.n2568\,
            ltout => OPEN,
            carryin => \nx.n10755\,
            carryout => \nx.n10756\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_12_lut_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45441\,
            in2 => \N__39593\,
            in3 => \N__38073\,
            lcout => \nx.n2567\,
            ltout => OPEN,
            carryin => \nx.n10756\,
            carryout => \nx.n10757\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_13_lut_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45026\,
            in2 => \N__38066\,
            in3 => \N__38025\,
            lcout => \nx.n2566\,
            ltout => OPEN,
            carryin => \nx.n10757\,
            carryout => \nx.n10758\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_14_lut_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45442\,
            in2 => \N__39728\,
            in3 => \N__38010\,
            lcout => \nx.n2565\,
            ltout => OPEN,
            carryin => \nx.n10758\,
            carryout => \nx.n10759\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_15_lut_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45027\,
            in2 => \N__38007\,
            in3 => \N__37977\,
            lcout => \nx.n2564\,
            ltout => OPEN,
            carryin => \nx.n10759\,
            carryout => \nx.n10760\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_16_lut_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45443\,
            in2 => \N__37973\,
            in3 => \N__37935\,
            lcout => \nx.n2563\,
            ltout => OPEN,
            carryin => \nx.n10760\,
            carryout => \nx.n10761\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_17_lut_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45028\,
            in2 => \N__39380\,
            in3 => \N__38319\,
            lcout => \nx.n2562\,
            ltout => OPEN,
            carryin => \nx.n10761\,
            carryout => \nx.n10762\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_18_lut_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38316\,
            in2 => \N__45438\,
            in3 => \N__38298\,
            lcout => \nx.n2561\,
            ltout => OPEN,
            carryin => \bfn_12_22_0_\,
            carryout => \nx.n10763\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_19_lut_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38291\,
            in2 => \N__45437\,
            in3 => \N__38259\,
            lcout => \nx.n2560\,
            ltout => OPEN,
            carryin => \nx.n10763\,
            carryout => \nx.n10764\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_20_lut_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38256\,
            in2 => \N__45439\,
            in3 => \N__38223\,
            lcout => \nx.n2559\,
            ltout => OPEN,
            carryin => \nx.n10764\,
            carryout => \nx.n10765\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_21_lut_LC_12_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45036\,
            in2 => \N__38220\,
            in3 => \N__38190\,
            lcout => \nx.n2558\,
            ltout => OPEN,
            carryin => \nx.n10765\,
            carryout => \nx.n10766\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_22_lut_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45023\,
            in2 => \N__39693\,
            in3 => \N__38175\,
            lcout => \nx.n2557\,
            ltout => OPEN,
            carryin => \nx.n10766\,
            carryout => \nx.n10767\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1741_23_lut_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__45024\,
            in1 => \N__41538\,
            in2 => \N__39549\,
            in3 => \N__38172\,
            lcout => \nx.n2588\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i14_4_lut_adj_51_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43852\,
            in1 => \N__43936\,
            in2 => \N__43451\,
            in3 => \N__43399\,
            lcout => \nx.n33_adj_644\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_adj_47_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43899\,
            in1 => \N__44147\,
            in2 => \N__45810\,
            in3 => \N__38349\,
            lcout => \nx.n34_adj_641\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1559_3_lut_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40057\,
            in2 => \N__40035\,
            in3 => \N__41932\,
            lcout => \nx.n2308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i16_4_lut_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39949\,
            in1 => \N__42208\,
            in2 => \N__38475\,
            in3 => \N__38466\,
            lcout => OPEN,
            ltout => \nx.n34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i17_4_lut_LC_12_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38403\,
            in1 => \N__38409\,
            in2 => \N__38343\,
            in3 => \N__38340\,
            lcout => \nx.n2225\,
            ltout => \nx.n2225_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1556_3_lut_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39963\,
            in2 => \N__38331\,
            in3 => \N__39983\,
            lcout => \nx.n2305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1560_3_lut_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39804\,
            in1 => \N__39858\,
            in2 => \_gnd_net_\,
            in3 => \N__41928\,
            lcout => \nx.n2309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1558_3_lut_LC_12_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39999\,
            in2 => \N__41957\,
            in3 => \N__40022\,
            lcout => \nx.n2307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1555_3_lut_LC_12_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39950\,
            in2 => \N__39933\,
            in3 => \N__41933\,
            lcout => \nx.n2304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i6426_2_lut_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43567\,
            in2 => \_gnd_net_\,
            in3 => \N__43486\,
            lcout => \nx.n9650\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_4_lut_adj_78_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__41506\,
            in1 => \N__40018\,
            in2 => \N__42124\,
            in3 => \N__42076\,
            lcout => \nx.n31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i10_4_lut_adj_77_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40141\,
            in1 => \N__40090\,
            in2 => \N__42013\,
            in3 => \N__40376\,
            lcout => \nx.n28_adj_601\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_prev_i12_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38460\,
            lcout => neopxl_color_prev_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48439\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i12_4_lut_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40273\,
            in1 => \N__39910\,
            in2 => \N__42056\,
            in3 => \N__39982\,
            lcout => \nx.n30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i4_3_lut_adj_79_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__39857\,
            in1 => \_gnd_net_\,
            in2 => \N__40059\,
            in3 => \N__42169\,
            lcout => \nx.n22_adj_604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_adj_223_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__40806\,
            in1 => \N__47711\,
            in2 => \_gnd_net_\,
            in3 => \N__47678\,
            lcout => n7442,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_counter_1104__i0_LC_12_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38396\,
            in2 => \_gnd_net_\,
            in3 => \N__38382\,
            lcout => delay_counter_0,
            ltout => OPEN,
            carryin => \bfn_12_26_0_\,
            carryout => n10517,
            clk => \N__48445\,
            ce => \N__40812\,
            sr => \N__38976\
        );

    \delay_counter_1104__i1_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38379\,
            in2 => \_gnd_net_\,
            in3 => \N__38367\,
            lcout => delay_counter_1,
            ltout => OPEN,
            carryin => n10517,
            carryout => n10518,
            clk => \N__48445\,
            ce => \N__40812\,
            sr => \N__38976\
        );

    \delay_counter_1104__i2_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38364\,
            in2 => \_gnd_net_\,
            in3 => \N__38352\,
            lcout => delay_counter_2,
            ltout => OPEN,
            carryin => n10518,
            carryout => n10519,
            clk => \N__48445\,
            ce => \N__40812\,
            sr => \N__38976\
        );

    \delay_counter_1104__i3_LC_12_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38613\,
            in2 => \_gnd_net_\,
            in3 => \N__38601\,
            lcout => delay_counter_3,
            ltout => OPEN,
            carryin => n10519,
            carryout => n10520,
            clk => \N__48445\,
            ce => \N__40812\,
            sr => \N__38976\
        );

    \delay_counter_1104__i4_LC_12_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38598\,
            in2 => \_gnd_net_\,
            in3 => \N__38586\,
            lcout => delay_counter_4,
            ltout => OPEN,
            carryin => n10520,
            carryout => n10521,
            clk => \N__48445\,
            ce => \N__40812\,
            sr => \N__38976\
        );

    \delay_counter_1104__i5_LC_12_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38583\,
            in2 => \_gnd_net_\,
            in3 => \N__38571\,
            lcout => delay_counter_5,
            ltout => OPEN,
            carryin => n10521,
            carryout => n10522,
            clk => \N__48445\,
            ce => \N__40812\,
            sr => \N__38976\
        );

    \delay_counter_1104__i6_LC_12_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38568\,
            in2 => \_gnd_net_\,
            in3 => \N__38556\,
            lcout => delay_counter_6,
            ltout => OPEN,
            carryin => n10522,
            carryout => n10523,
            clk => \N__48445\,
            ce => \N__40812\,
            sr => \N__38976\
        );

    \delay_counter_1104__i7_LC_12_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38553\,
            in2 => \_gnd_net_\,
            in3 => \N__38541\,
            lcout => delay_counter_7,
            ltout => OPEN,
            carryin => n10523,
            carryout => n10524,
            clk => \N__48445\,
            ce => \N__40812\,
            sr => \N__38976\
        );

    \delay_counter_1104__i8_LC_12_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38538\,
            in2 => \_gnd_net_\,
            in3 => \N__38526\,
            lcout => delay_counter_8,
            ltout => OPEN,
            carryin => \bfn_12_27_0_\,
            carryout => n10525,
            clk => \N__48447\,
            ce => \N__40820\,
            sr => \N__38993\
        );

    \delay_counter_1104__i9_LC_12_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38522\,
            in2 => \_gnd_net_\,
            in3 => \N__38508\,
            lcout => delay_counter_9,
            ltout => OPEN,
            carryin => n10525,
            carryout => n10526,
            clk => \N__48447\,
            ce => \N__40820\,
            sr => \N__38993\
        );

    \delay_counter_1104__i10_LC_12_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38505\,
            in2 => \_gnd_net_\,
            in3 => \N__38493\,
            lcout => delay_counter_10,
            ltout => OPEN,
            carryin => n10526,
            carryout => n10527,
            clk => \N__48447\,
            ce => \N__40820\,
            sr => \N__38993\
        );

    \delay_counter_1104__i11_LC_12_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38490\,
            in2 => \_gnd_net_\,
            in3 => \N__38478\,
            lcout => delay_counter_11,
            ltout => OPEN,
            carryin => n10527,
            carryout => n10528,
            clk => \N__48447\,
            ce => \N__40820\,
            sr => \N__38993\
        );

    \delay_counter_1104__i12_LC_12_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38760\,
            in2 => \_gnd_net_\,
            in3 => \N__38748\,
            lcout => delay_counter_12,
            ltout => OPEN,
            carryin => n10528,
            carryout => n10529,
            clk => \N__48447\,
            ce => \N__40820\,
            sr => \N__38993\
        );

    \delay_counter_1104__i13_LC_12_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38745\,
            in2 => \_gnd_net_\,
            in3 => \N__38733\,
            lcout => delay_counter_13,
            ltout => OPEN,
            carryin => n10529,
            carryout => n10530,
            clk => \N__48447\,
            ce => \N__40820\,
            sr => \N__38993\
        );

    \delay_counter_1104__i14_LC_12_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38730\,
            in2 => \_gnd_net_\,
            in3 => \N__38718\,
            lcout => delay_counter_14,
            ltout => OPEN,
            carryin => n10530,
            carryout => n10531,
            clk => \N__48447\,
            ce => \N__40820\,
            sr => \N__38993\
        );

    \delay_counter_1104__i15_LC_12_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38708\,
            in2 => \_gnd_net_\,
            in3 => \N__38694\,
            lcout => delay_counter_15,
            ltout => OPEN,
            carryin => n10531,
            carryout => n10532,
            clk => \N__48447\,
            ce => \N__40820\,
            sr => \N__38993\
        );

    \delay_counter_1104__i16_LC_12_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38690\,
            in2 => \_gnd_net_\,
            in3 => \N__38676\,
            lcout => delay_counter_16,
            ltout => OPEN,
            carryin => \bfn_12_28_0_\,
            carryout => n10533,
            clk => \N__48448\,
            ce => \N__40813\,
            sr => \N__38989\
        );

    \delay_counter_1104__i17_LC_12_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38669\,
            in2 => \_gnd_net_\,
            in3 => \N__38655\,
            lcout => delay_counter_17,
            ltout => OPEN,
            carryin => n10533,
            carryout => n10534,
            clk => \N__48448\,
            ce => \N__40813\,
            sr => \N__38989\
        );

    \delay_counter_1104__i18_LC_12_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38648\,
            in2 => \_gnd_net_\,
            in3 => \N__38634\,
            lcout => delay_counter_18,
            ltout => OPEN,
            carryin => n10534,
            carryout => n10535,
            clk => \N__48448\,
            ce => \N__40813\,
            sr => \N__38989\
        );

    \delay_counter_1104__i19_LC_12_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38630\,
            in2 => \_gnd_net_\,
            in3 => \N__38616\,
            lcout => delay_counter_19,
            ltout => OPEN,
            carryin => n10535,
            carryout => n10536,
            clk => \N__48448\,
            ce => \N__40813\,
            sr => \N__38989\
        );

    \delay_counter_1104__i20_LC_12_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38888\,
            in2 => \_gnd_net_\,
            in3 => \N__38874\,
            lcout => delay_counter_20,
            ltout => OPEN,
            carryin => n10536,
            carryout => n10537,
            clk => \N__48448\,
            ce => \N__40813\,
            sr => \N__38989\
        );

    \delay_counter_1104__i21_LC_12_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38871\,
            in2 => \_gnd_net_\,
            in3 => \N__38859\,
            lcout => delay_counter_21,
            ltout => OPEN,
            carryin => n10537,
            carryout => n10538,
            clk => \N__48448\,
            ce => \N__40813\,
            sr => \N__38989\
        );

    \delay_counter_1104__i22_LC_12_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38855\,
            in2 => \_gnd_net_\,
            in3 => \N__38841\,
            lcout => delay_counter_22,
            ltout => OPEN,
            carryin => n10538,
            carryout => n10539,
            clk => \N__48448\,
            ce => \N__40813\,
            sr => \N__38989\
        );

    \delay_counter_1104__i23_LC_12_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38838\,
            in2 => \_gnd_net_\,
            in3 => \N__38826\,
            lcout => delay_counter_23,
            ltout => OPEN,
            carryin => n10539,
            carryout => n10540,
            clk => \N__48448\,
            ce => \N__40813\,
            sr => \N__38989\
        );

    \delay_counter_1104__i24_LC_12_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38823\,
            in2 => \_gnd_net_\,
            in3 => \N__38811\,
            lcout => delay_counter_24,
            ltout => OPEN,
            carryin => \bfn_12_29_0_\,
            carryout => n10541,
            clk => \N__48449\,
            ce => \N__40824\,
            sr => \N__38994\
        );

    \delay_counter_1104__i25_LC_12_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38808\,
            in2 => \_gnd_net_\,
            in3 => \N__38796\,
            lcout => delay_counter_25,
            ltout => OPEN,
            carryin => n10541,
            carryout => n10542,
            clk => \N__48449\,
            ce => \N__40824\,
            sr => \N__38994\
        );

    \delay_counter_1104__i26_LC_12_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38793\,
            in2 => \_gnd_net_\,
            in3 => \N__38781\,
            lcout => delay_counter_26,
            ltout => OPEN,
            carryin => n10542,
            carryout => n10543,
            clk => \N__48449\,
            ce => \N__40824\,
            sr => \N__38994\
        );

    \delay_counter_1104__i27_LC_12_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38777\,
            in2 => \_gnd_net_\,
            in3 => \N__38763\,
            lcout => delay_counter_27,
            ltout => OPEN,
            carryin => n10543,
            carryout => n10544,
            clk => \N__48449\,
            ce => \N__40824\,
            sr => \N__38994\
        );

    \delay_counter_1104__i28_LC_12_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39042\,
            in2 => \_gnd_net_\,
            in3 => \N__39030\,
            lcout => delay_counter_28,
            ltout => OPEN,
            carryin => n10544,
            carryout => n10545,
            clk => \N__48449\,
            ce => \N__40824\,
            sr => \N__38994\
        );

    \delay_counter_1104__i29_LC_12_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39027\,
            in2 => \_gnd_net_\,
            in3 => \N__39015\,
            lcout => delay_counter_29,
            ltout => OPEN,
            carryin => n10545,
            carryout => n10546,
            clk => \N__48449\,
            ce => \N__40824\,
            sr => \N__38994\
        );

    \delay_counter_1104__i30_LC_12_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39012\,
            in2 => \_gnd_net_\,
            in3 => \N__39000\,
            lcout => delay_counter_30,
            ltout => OPEN,
            carryin => n10546,
            carryout => n10547,
            clk => \N__48449\,
            ce => \N__40824\,
            sr => \N__38994\
        );

    \delay_counter_1104__i31_LC_12_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47707\,
            in2 => \_gnd_net_\,
            in3 => \N__38997\,
            lcout => delay_counter_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48449\,
            ce => \N__40824\,
            sr => \N__38994\
        );

    \i1_3_lut_4_lut_adj_245_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__42262\,
            in1 => \N__46980\,
            in2 => \N__40665\,
            in3 => \N__46657\,
            lcout => n10_adj_779,
            ltout => \n10_adj_779_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_169_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001001100"
        )
    port map (
            in0 => \N__42455\,
            in1 => \N__47505\,
            in2 => \N__38955\,
            in3 => \N__47994\,
            lcout => OPEN,
            ltout => \n7290_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i10_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__38952\,
            in1 => \N__38927\,
            in2 => \N__38946\,
            in3 => \N__46535\,
            lcout => pin_out_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48428\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_230_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47168\,
            in2 => \_gnd_net_\,
            in3 => \N__47236\,
            lcout => n7135,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_189_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__47235\,
            in1 => \N__48137\,
            in2 => \N__47176\,
            in3 => \N__49017\,
            lcout => n7155,
            ltout => \n7155_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2954_3_lut_4_lut_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__42252\,
            in1 => \N__42326\,
            in2 => \N__39087\,
            in3 => \N__46940\,
            lcout => n6174,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2970_3_lut_4_lut_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__42327\,
            in1 => \N__46970\,
            in2 => \N__40362\,
            in3 => \N__46776\,
            lcout => n6190,
            ltout => \n6190_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_197_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000101010"
        )
    port map (
            in0 => \N__47458\,
            in1 => \N__42715\,
            in2 => \N__39075\,
            in3 => \N__47290\,
            lcout => n7334,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2950_3_lut_4_lut_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__40351\,
            in1 => \N__42261\,
            in2 => \N__46979\,
            in3 => \N__40656\,
            lcout => n6170,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_217_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__47238\,
            in1 => \N__49803\,
            in2 => \N__47181\,
            in3 => \N__48149\,
            lcout => n11481,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6193_2_lut_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__50771\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48697\,
            lcout => n9415,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2966_3_lut_4_lut_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__46774\,
            in1 => \N__40648\,
            in2 => \N__46978\,
            in3 => \N__40354\,
            lcout => n6186,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i404_4_lut_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__40609\,
            in1 => \N__39248\,
            in2 => \N__50358\,
            in3 => \N__48920\,
            lcout => n2337,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2962_3_lut_4_lut_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__40353\,
            in1 => \N__46775\,
            in2 => \N__46745\,
            in3 => \N__46969\,
            lcout => n6182,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_270_i8_2_lut_3_lut_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__48696\,
            in1 => \N__50770\,
            in2 => \_gnd_net_\,
            in3 => \N__50533\,
            lcout => n8_adj_723,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_pin_0__bdd_4_lut_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__40703\,
            in1 => \N__50262\,
            in2 => \N__39194\,
            in3 => \N__48919\,
            lcout => OPEN,
            ltout => \n13480_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n13480_bdd_4_lut_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__39249\,
            in1 => \N__50348\,
            in2 => \N__39231\,
            in3 => \N__40583\,
            lcout => n13483,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__50005\,
            in1 => \N__49758\,
            in2 => \_gnd_net_\,
            in3 => \N__49508\,
            lcout => OPEN,
            ltout => \current_pin_7__N_157_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i16_4_lut_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47617\,
            in1 => \N__39093\,
            in2 => \N__39228\,
            in3 => \N__50006\,
            lcout => n45_adj_772,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i356_3_lut_4_lut_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__47797\,
            in1 => \N__39225\,
            in2 => \N__42626\,
            in3 => \N__42831\,
            lcout => OPEN,
            ltout => \n2289_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__47992\,
            in1 => \N__39195\,
            in2 => \N__39153\,
            in3 => \N__40610\,
            lcout => n39,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i392_4_lut_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__47991\,
            in1 => \N__50616\,
            in2 => \N__39150\,
            in3 => \N__47796\,
            lcout => n2325,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9515_3_lut_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50756\,
            in1 => \N__39108\,
            in2 => \_gnd_net_\,
            in3 => \N__39561\,
            lcout => OPEN,
            ltout => \n13364_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i37_4_lut_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000111100"
        )
    port map (
            in0 => \N__47808\,
            in1 => \N__46451\,
            in2 => \N__39096\,
            in3 => \N__48682\,
            lcout => n150,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6204_2_lut_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__50337\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49016\,
            lcout => n9426,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9511_3_lut_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50569\,
            in1 => \N__40959\,
            in2 => \_gnd_net_\,
            in3 => \N__39570\,
            lcout => n13360,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1762_3_lut_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39555\,
            in2 => \N__39297\,
            in3 => \N__39507\,
            lcout => \nx.n2607\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1682_3_lut_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41881\,
            in2 => \N__41301\,
            in3 => \N__41653\,
            lcout => \nx.n2495\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9538_3_lut_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40998\,
            in2 => \N__41663\,
            in3 => \N__41012\,
            lcout => \nx.n2503\,
            ltout => \nx.n2503_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_adj_44_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39268\,
            in1 => \N__39316\,
            in2 => \N__39333\,
            in3 => \N__39292\,
            lcout => \nx.n36_adj_636\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9540_3_lut_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43663\,
            in2 => \N__41664\,
            in3 => \N__41451\,
            lcout => \nx.n2502\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1695_rep_30_3_lut_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41163\,
            in2 => \N__41203\,
            in3 => \N__41640\,
            lcout => \nx.n2508\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9534_3_lut_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41085\,
            in2 => \N__41662\,
            in3 => \N__41109\,
            lcout => \nx.n2506\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_205_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__49753\,
            in1 => \N__39778\,
            in2 => \_gnd_net_\,
            in3 => \N__50001\,
            lcout => n22_adj_730,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1685_3_lut_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41366\,
            in2 => \N__41665\,
            in3 => \N__41346\,
            lcout => \nx.n2498\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1622_3_lut_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43941\,
            in2 => \N__43917\,
            in3 => \N__44081\,
            lcout => \nx.n2403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1623_3_lut_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43956\,
            in2 => \N__43986\,
            in3 => \N__44082\,
            lcout => \nx.n2404\,
            ltout => \nx.n2404_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i14_4_lut_adj_61_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43232\,
            in1 => \N__41104\,
            in2 => \N__39705\,
            in3 => \N__41362\,
            lcout => \nx.n34_adj_657\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i1_2_lut_adj_57_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41537\,
            in3 => \N__39686\,
            lcout => OPEN,
            ltout => \nx.n22_adj_637_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i16_4_lut_adj_45_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39663\,
            in1 => \N__39586\,
            in2 => \N__39642\,
            in3 => \N__39639\,
            lcout => \nx.n37_adj_638\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9544_3_lut_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__41669\,
            in1 => \N__41394\,
            in2 => \N__41423\,
            in3 => \_gnd_net_\,
            lcout => \nx.n2500\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1618_3_lut_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43752\,
            in2 => \N__44116\,
            in3 => \N__43766\,
            lcout => \nx.n2399\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1626_3_lut_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43425\,
            in2 => \N__44117\,
            in3 => \N__43447\,
            lcout => \nx.n2407\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1627_3_lut_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43490\,
            in2 => \N__43470\,
            in3 => \N__44086\,
            lcout => \nx.n2408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1553_3_lut_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39891\,
            in2 => \N__39918\,
            in3 => \N__41953\,
            lcout => \nx.n2302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1551_3_lut_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40278\,
            in2 => \N__41976\,
            in3 => \N__40251\,
            lcout => \nx.n2300\,
            ltout => \nx.n2300_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i13_4_lut_adj_50_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43810\,
            in1 => \N__43975\,
            in2 => \N__39879\,
            in3 => \N__43369\,
            lcout => OPEN,
            ltout => \nx.n32_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i18_4_lut_adj_53_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39876\,
            in1 => \N__39870\,
            in2 => \N__39864\,
            in3 => \N__42144\,
            lcout => \nx.n2324\,
            ltout => \nx.n2324_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9497_3_lut_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43353\,
            in2 => \N__39861\,
            in3 => \N__43370\,
            lcout => \nx.n2405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i9489_3_lut_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43853\,
            in2 => \N__43833\,
            in3 => \N__44090\,
            lcout => \nx.n2401\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_2_lut_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39856\,
            in2 => \_gnd_net_\,
            in3 => \N__39798\,
            lcout => \nx.n2277\,
            ltout => OPEN,
            carryin => \bfn_13_23_0_\,
            carryout => \nx.n10690\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_3_lut_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40058\,
            in2 => \_gnd_net_\,
            in3 => \N__40026\,
            lcout => \nx.n2276\,
            ltout => OPEN,
            carryin => \nx.n10690\,
            carryout => \nx.n10691\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_4_lut_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45571\,
            in2 => \N__40023\,
            in3 => \N__39993\,
            lcout => \nx.n2275\,
            ltout => OPEN,
            carryin => \nx.n10691\,
            carryout => \nx.n10692\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_5_lut_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44644\,
            in2 => \N__41513\,
            in3 => \N__39990\,
            lcout => \nx.n2274\,
            ltout => OPEN,
            carryin => \nx.n10692\,
            carryout => \nx.n10693\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_6_lut_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45572\,
            in2 => \N__39987\,
            in3 => \N__39957\,
            lcout => \nx.n2273\,
            ltout => OPEN,
            carryin => \nx.n10693\,
            carryout => \nx.n10694\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_7_lut_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44645\,
            in2 => \N__39954\,
            in3 => \N__39924\,
            lcout => \nx.n2272\,
            ltout => OPEN,
            carryin => \nx.n10694\,
            carryout => \nx.n10695\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_8_lut_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42209\,
            in2 => \N__45019\,
            in3 => \N__39921\,
            lcout => \nx.n2271\,
            ltout => OPEN,
            carryin => \nx.n10695\,
            carryout => \nx.n10696\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_9_lut_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39911\,
            in2 => \N__45731\,
            in3 => \N__39885\,
            lcout => \nx.n2270\,
            ltout => OPEN,
            carryin => \nx.n10696\,
            carryout => \nx.n10697\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_10_lut_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45218\,
            in2 => \N__42129\,
            in3 => \N__39882\,
            lcout => \nx.n2269\,
            ltout => OPEN,
            carryin => \bfn_13_24_0_\,
            carryout => \nx.n10698\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_11_lut_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45227\,
            in2 => \N__40277\,
            in3 => \N__40242\,
            lcout => \nx.n2268\,
            ltout => OPEN,
            carryin => \nx.n10698\,
            carryout => \nx.n10699\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_12_lut_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45219\,
            in2 => \N__42089\,
            in3 => \N__40239\,
            lcout => \nx.n2267\,
            ltout => OPEN,
            carryin => \nx.n10699\,
            carryout => \nx.n10700\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_13_lut_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42052\,
            in2 => \N__45568\,
            in3 => \N__40236\,
            lcout => \nx.n2266\,
            ltout => OPEN,
            carryin => \nx.n10700\,
            carryout => \nx.n10701\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_14_lut_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45223\,
            in2 => \N__42182\,
            in3 => \N__40233\,
            lcout => \nx.n2265\,
            ltout => OPEN,
            carryin => \nx.n10701\,
            carryout => \nx.n10702\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_15_lut_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40229\,
            in2 => \N__45569\,
            in3 => \N__40194\,
            lcout => \nx.n2264\,
            ltout => OPEN,
            carryin => \nx.n10702\,
            carryout => \nx.n10703\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_16_lut_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40191\,
            in2 => \N__45570\,
            in3 => \N__40155\,
            lcout => \nx.n2263\,
            ltout => OPEN,
            carryin => \nx.n10703\,
            carryout => \nx.n10704\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_17_lut_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45231\,
            in2 => \N__40152\,
            in3 => \N__40110\,
            lcout => \nx.n2262\,
            ltout => OPEN,
            carryin => \nx.n10704\,
            carryout => \nx.n10705\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_18_lut_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44859\,
            in2 => \N__40107\,
            in3 => \N__40065\,
            lcout => \nx.n2261\,
            ltout => OPEN,
            carryin => \bfn_13_25_0_\,
            carryout => \nx.n10706\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_19_lut_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44860\,
            in2 => \N__42020\,
            in3 => \N__40062\,
            lcout => \nx.n2260\,
            ltout => OPEN,
            carryin => \nx.n10706\,
            carryout => \nx.n10707\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1540_20_lut_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__44861\,
            in1 => \N__41975\,
            in2 => \N__40383\,
            in3 => \N__40365\,
            lcout => \nx.n2291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1628_3_lut_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43509\,
            in2 => \N__44123\,
            in3 => \N__43571\,
            lcout => \nx.n2409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2958_3_lut_4_lut_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__50128\,
            in1 => \N__46941\,
            in2 => \N__42264\,
            in3 => \N__40346\,
            lcout => n6178,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i9_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__40287\,
            in1 => \N__40296\,
            in2 => \N__42494\,
            in3 => \N__46517\,
            lcout => pin_out_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48429\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2946_3_lut_4_lut_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__42260\,
            in1 => \N__46942\,
            in2 => \N__46746\,
            in3 => \N__40347\,
            lcout => n6166,
            ltout => \n6166_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_167_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001001100"
        )
    port map (
            in0 => \N__42456\,
            in1 => \N__47526\,
            in2 => \N__40290\,
            in3 => \N__42726\,
            lcout => n7286,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_282_i7_2_lut_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48691\,
            in2 => \_gnd_net_\,
            in3 => \N__50758\,
            lcout => n7_adj_753,
            ltout => \n7_adj_753_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2944_3_lut_4_lut_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__46943\,
            in1 => \N__46743\,
            in2 => \N__40281\,
            in3 => \N__46677\,
            lcout => n6164,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i13_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__42270\,
            in1 => \N__42284\,
            in2 => \N__48073\,
            in3 => \N__46516\,
            lcout => pin_out_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48429\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2968_3_lut_4_lut_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__42324\,
            in1 => \N__46916\,
            in2 => \N__46688\,
            in3 => \N__46788\,
            lcout => n6188,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_1098_i21_2_lut_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__50354\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50557\,
            lcout => n21_adj_714,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12_4_lut_adj_238_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__40479\,
            in1 => \N__40671\,
            in2 => \N__49349\,
            in3 => \N__47795\,
            lcout => n41,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_1100_i21_2_lut_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__50355\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50558\,
            lcout => n21_adj_741,
            ltout => \n21_adj_741_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40449\,
            in2 => \N__40404\,
            in3 => \N__48148\,
            lcout => n7128,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_879_i9_2_lut_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50263\,
            in2 => \_gnd_net_\,
            in3 => \N__48921\,
            lcout => n9_adj_733,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_903_i11_2_lut_4_lut_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__50264\,
            in1 => \N__50722\,
            in2 => \N__48994\,
            in3 => \N__50544\,
            lcout => n11_adj_743,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_231_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__48666\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47263\,
            lcout => n14_adj_752,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_274_i8_2_lut_3_lut_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__50532\,
            in1 => \N__50726\,
            in2 => \_gnd_net_\,
            in3 => \N__48671\,
            lcout => n8_adj_746,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_215_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__50721\,
            in1 => \N__50531\,
            in2 => \N__48695\,
            in3 => \N__47264\,
            lcout => n7150,
            ltout => \n7150_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i422_4_lut_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100000000"
        )
    port map (
            in0 => \N__50265\,
            in1 => \N__49004\,
            in2 => \N__40710\,
            in3 => \N__40707\,
            lcout => n2355,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_273_i7_2_lut_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__48670\,
            in1 => \_gnd_net_\,
            in2 => \N__50757\,
            in3 => \_gnd_net_\,
            lcout => n7_adj_719,
            ltout => \n7_adj_719_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2964_3_lut_4_lut_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__40655\,
            in1 => \N__46977\,
            in2 => \N__40614\,
            in3 => \N__46687\,
            lcout => n6184,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i410_4_lut_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__40611\,
            in1 => \N__50353\,
            in2 => \N__40593\,
            in3 => \N__48985\,
            lcout => OPEN,
            ltout => \n2343_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40563\,
            in1 => \N__42918\,
            in2 => \N__40557\,
            in3 => \N__47034\,
            lcout => n53_adj_769,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_4_lut_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101010"
        )
    port map (
            in0 => \N__40554\,
            in1 => \N__40548\,
            in2 => \N__48197\,
            in3 => \N__47798\,
            lcout => n43,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_235_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__42765\,
            in1 => \N__50352\,
            in2 => \N__40986\,
            in3 => \N__48984\,
            lcout => n2361,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_adj_237_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__42927\,
            in1 => \N__47799\,
            in2 => \N__40518\,
            in3 => \N__40485\,
            lcout => n33,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_pin_0__bdd_4_lut_9624_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010110000"
        )
    port map (
            in0 => \N__40928\,
            in1 => \N__50333\,
            in2 => \N__49040\,
            in3 => \N__42807\,
            lcout => OPEN,
            ltout => \n13474_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n13474_bdd_4_lut_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__50334\,
            in1 => \N__40953\,
            in2 => \N__40989\,
            in3 => \N__40985\,
            lcout => n13477,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_236_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011001100"
        )
    port map (
            in0 => \N__50335\,
            in1 => \N__40952\,
            in2 => \N__42768\,
            in3 => \N__49014\,
            lcout => n2367,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i446_4_lut_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__42766\,
            in1 => \N__50336\,
            in2 => \N__40932\,
            in3 => \N__49015\,
            lcout => OPEN,
            ltout => \n2379_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i23_4_lut_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40911\,
            in1 => \N__40905\,
            in2 => \N__40899\,
            in3 => \N__40896\,
            lcout => n52_adj_770,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_209_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__49985\,
            in1 => \N__49775\,
            in2 => \_gnd_net_\,
            in3 => \N__40887\,
            lcout => n22_adj_732,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_219_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__49774\,
            in1 => \N__49984\,
            in2 => \_gnd_net_\,
            in3 => \N__49553\,
            lcout => n7232,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i26_4_lut_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47727\,
            in1 => \N__40773\,
            in2 => \N__43332\,
            in3 => \N__40764\,
            lcout => n55_adj_767,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_201_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010101000"
        )
    port map (
            in0 => \N__40755\,
            in1 => \N__49986\,
            in2 => \N__49811\,
            in3 => \_gnd_net_\,
            lcout => n22_adj_728,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_212_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__47265\,
            in1 => \N__50755\,
            in2 => \N__48702\,
            in3 => \N__50556\,
            lcout => n7145,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_2_lut_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41283\,
            in2 => \_gnd_net_\,
            in3 => \N__41211\,
            lcout => \nx.n2477\,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => \nx.n10727\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_3_lut_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__41204\,
            in3 => \N__41157\,
            lcout => \nx.n2476\,
            ltout => OPEN,
            carryin => \nx.n10727\,
            carryout => \nx.n10728\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_4_lut_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45444\,
            in2 => \N__41146\,
            in3 => \N__41112\,
            lcout => \nx.n2475\,
            ltout => OPEN,
            carryin => \nx.n10728\,
            carryout => \nx.n10729\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_5_lut_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45447\,
            in2 => \N__41108\,
            in3 => \N__41079\,
            lcout => \nx.n2474\,
            ltout => OPEN,
            carryin => \nx.n10729\,
            carryout => \nx.n10730\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_6_lut_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45445\,
            in2 => \N__43595\,
            in3 => \N__41064\,
            lcout => \nx.n2473\,
            ltout => OPEN,
            carryin => \nx.n10730\,
            carryout => \nx.n10731\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_7_lut_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45448\,
            in2 => \N__41059\,
            in3 => \N__41016\,
            lcout => \nx.n2472\,
            ltout => OPEN,
            carryin => \nx.n10731\,
            carryout => \nx.n10732\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_8_lut_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45446\,
            in2 => \N__41013\,
            in3 => \N__40992\,
            lcout => \nx.n2471\,
            ltout => OPEN,
            carryin => \nx.n10732\,
            carryout => \nx.n10733\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_9_lut_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45449\,
            in2 => \N__43667\,
            in3 => \N__41445\,
            lcout => \nx.n2470\,
            ltout => OPEN,
            carryin => \nx.n10733\,
            carryout => \nx.n10734\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_10_lut_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43616\,
            in2 => \N__45732\,
            in3 => \N__41430\,
            lcout => \nx.n2469\,
            ltout => OPEN,
            carryin => \bfn_14_22_0_\,
            carryout => \nx.n10735\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_11_lut_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45584\,
            in2 => \N__41422\,
            in3 => \N__41388\,
            lcout => \nx.n2468\,
            ltout => OPEN,
            carryin => \nx.n10735\,
            carryout => \nx.n10736\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_12_lut_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45588\,
            in2 => \N__43688\,
            in3 => \N__41370\,
            lcout => \nx.n2467\,
            ltout => OPEN,
            carryin => \nx.n10736\,
            carryout => \nx.n10737\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_13_lut_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45585\,
            in2 => \N__41367\,
            in3 => \N__41337\,
            lcout => \nx.n2466\,
            ltout => OPEN,
            carryin => \nx.n10737\,
            carryout => \nx.n10738\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_14_lut_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45589\,
            in2 => \N__43228\,
            in3 => \N__41319\,
            lcout => \nx.n2465\,
            ltout => OPEN,
            carryin => \nx.n10738\,
            carryout => \nx.n10739\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_15_lut_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45586\,
            in2 => \N__43198\,
            in3 => \N__41304\,
            lcout => \nx.n2464\,
            ltout => OPEN,
            carryin => \nx.n10739\,
            carryout => \nx.n10740\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_16_lut_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45590\,
            in2 => \N__41882\,
            in3 => \N__41286\,
            lcout => \nx.n2463\,
            ltout => OPEN,
            carryin => \nx.n10740\,
            carryout => \nx.n10741\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_17_lut_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45587\,
            in2 => \N__41847\,
            in3 => \N__41814\,
            lcout => \nx.n2462\,
            ltout => OPEN,
            carryin => \nx.n10741\,
            carryout => \nx.n10742\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_18_lut_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45576\,
            in2 => \N__41811\,
            in3 => \N__41775\,
            lcout => \nx.n2461\,
            ltout => OPEN,
            carryin => \bfn_14_23_0_\,
            carryout => \nx.n10743\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_19_lut_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45578\,
            in2 => \N__41772\,
            in3 => \N__41733\,
            lcout => \nx.n2460\,
            ltout => OPEN,
            carryin => \nx.n10743\,
            carryout => \nx.n10744\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_20_lut_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45577\,
            in2 => \N__41730\,
            in3 => \N__41688\,
            lcout => \nx.n2459\,
            ltout => OPEN,
            carryin => \nx.n10744\,
            carryout => \nx.n10745\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_21_lut_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45579\,
            in2 => \N__41473\,
            in3 => \N__41673\,
            lcout => \nx.n2458\,
            ltout => OPEN,
            carryin => \nx.n10745\,
            carryout => \nx.n10746\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1674_22_lut_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__45580\,
            in1 => \N__44006\,
            in2 => \N__41670\,
            in3 => \N__41541\,
            lcout => \nx.n2489\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1557_3_lut_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41514\,
            in2 => \N__41487\,
            in3 => \N__41973\,
            lcout => \nx.n2306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1610_3_lut_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45777\,
            in2 => \N__45806\,
            in3 => \N__44098\,
            lcout => \nx.n2391\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1554_3_lut_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42222\,
            in2 => \N__42213\,
            in3 => \N__41972\,
            lcout => \nx.n2303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1548_3_lut_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42189\,
            in2 => \N__41991\,
            in3 => \N__42183\,
            lcout => \nx.n2297\,
            ltout => \nx.n2297_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i12_4_lut_adj_52_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__46039\,
            in1 => \N__43726\,
            in2 => \N__42156\,
            in3 => \N__42153\,
            lcout => \nx.n31_adj_645\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1552_3_lut_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42135\,
            in2 => \N__41990\,
            in3 => \N__42128\,
            lcout => \nx.n2301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1550_3_lut_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42099\,
            in2 => \N__42093\,
            in3 => \N__41981\,
            lcout => \nx.n2299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1549_3_lut_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__42063\,
            in1 => \_gnd_net_\,
            in2 => \N__41989\,
            in3 => \N__42057\,
            lcout => \nx.n2298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1543_3_lut_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42030\,
            in2 => \N__42024\,
            in3 => \N__41977\,
            lcout => \nx.n2292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1615_3_lut_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45990\,
            in2 => \N__46008\,
            in3 => \N__44099\,
            lcout => \nx.n2396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9330_4_lut_LC_14_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011101100"
        )
    port map (
            in0 => \N__46218\,
            in1 => \N__46238\,
            in2 => \N__46278\,
            in3 => \N__46257\,
            lcout => OPEN,
            ltout => \n13177_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9331_3_lut_LC_14_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__42333\,
            in1 => \_gnd_net_\,
            in2 => \N__42354\,
            in3 => \N__46353\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9329_4_lut_LC_14_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100000"
        )
    port map (
            in0 => \N__46256\,
            in1 => \N__46217\,
            in2 => \N__46239\,
            in3 => \N__46274\,
            lcout => n13176,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_173_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101010"
        )
    port map (
            in0 => \N__47524\,
            in1 => \N__42303\,
            in2 => \N__42641\,
            in3 => \N__43319\,
            lcout => n7298,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2952_3_lut_4_lut_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__46669\,
            in1 => \N__42325\,
            in2 => \N__42263\,
            in3 => \N__46871\,
            lcout => n6172,
            ltout => \n6172_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i12_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__42297\,
            in1 => \N__48028\,
            in2 => \N__42291\,
            in3 => \N__46487\,
            lcout => pin_out_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_175_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000001010"
        )
    port map (
            in0 => \N__47525\,
            in1 => \N__50342\,
            in2 => \N__42288\,
            in3 => \N__48096\,
            lcout => n7302,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2956_3_lut_4_lut_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__50129\,
            in1 => \N__42256\,
            in2 => \N__46927\,
            in3 => \N__46670\,
            lcout => n6176,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_181_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101010"
        )
    port map (
            in0 => \N__47519\,
            in1 => \N__46592\,
            in2 => \N__42633\,
            in3 => \N__42974\,
            lcout => n7314,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_177_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011001100"
        )
    port map (
            in0 => \N__43318\,
            in1 => \N__47523\,
            in2 => \N__47997\,
            in3 => \N__42518\,
            lcout => OPEN,
            ltout => \n7306_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i14_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__42519\,
            in1 => \N__47839\,
            in2 => \N__42510\,
            in3 => \N__46482\,
            lcout => pin_out_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9314_3_lut_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42487\,
            in1 => \N__42400\,
            in2 => \_gnd_net_\,
            in3 => \N__48995\,
            lcout => OPEN,
            ltout => \n13161_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n13468_bdd_4_lut_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__50565\,
            in1 => \N__42471\,
            in2 => \N__42459\,
            in3 => \N__48006\,
            lcout => n13471,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_165_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110000"
        )
    port map (
            in0 => \N__42454\,
            in1 => \N__42425\,
            in2 => \N__47534\,
            in3 => \N__42625\,
            lcout => OPEN,
            ltout => \n7282_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i8_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__46481\,
            in1 => \N__42426\,
            in2 => \N__42414\,
            in3 => \N__42401\,
            lcout => pin_out_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_186_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000101010"
        )
    port map (
            in0 => \N__47506\,
            in1 => \N__47996\,
            in2 => \N__42387\,
            in3 => \N__42972\,
            lcout => OPEN,
            ltout => \n7322_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i18_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__42386\,
            in1 => \N__42538\,
            in2 => \N__42372\,
            in3 => \N__46483\,
            lcout => pin_out_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9513_3_lut_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42369\,
            in1 => \N__50713\,
            in2 => \_gnd_net_\,
            in3 => \N__42363\,
            lcout => n13362,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_276_i8_2_lut_3_lut_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__48680\,
            in1 => \N__50714\,
            in2 => \_gnd_net_\,
            in3 => \N__50535\,
            lcout => n8_adj_747,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__50130\,
            in1 => \N__47271\,
            in2 => \N__46692\,
            in3 => \N__46777\,
            lcout => n12135,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i20_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__42561\,
            in1 => \N__42575\,
            in2 => \N__42863\,
            in3 => \N__46450\,
            lcout => pin_out_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i452_3_lut_4_lut_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__42830\,
            in1 => \N__42609\,
            in2 => \N__49233\,
            in3 => \N__49123\,
            lcout => n2385,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i440_3_lut_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__47993\,
            in1 => \N__42800\,
            in2 => \_gnd_net_\,
            in3 => \N__42767\,
            lcout => n2373,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i16_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__42735\,
            in1 => \N__43085\,
            in2 => \N__46602\,
            in3 => \N__46448\,
            lcout => pin_out_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_184_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001001100"
        )
    port map (
            in0 => \N__42665\,
            in1 => \N__47494\,
            in2 => \N__42725\,
            in3 => \N__42973\,
            lcout => OPEN,
            ltout => \n7318_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i17_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__43048\,
            in1 => \N__42666\,
            in2 => \N__42648\,
            in3 => \N__46449\,
            lcout => pin_out_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_193_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100000000"
        )
    port map (
            in0 => \N__47298\,
            in1 => \N__42610\,
            in2 => \N__42576\,
            in3 => \N__47493\,
            lcout => n7330,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_pin_0__bdd_4_lut_9596_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__42542\,
            in1 => \N__49000\,
            in2 => \N__42998\,
            in3 => \N__50346\,
            lcout => OPEN,
            ltout => \n13438_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n13438_bdd_4_lut_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__50347\,
            in1 => \N__43084\,
            in2 => \N__43068\,
            in3 => \N__43052\,
            lcout => OPEN,
            ltout => \n13441_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9295_3_lut_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43338\,
            in2 => \N__43029\,
            in3 => \N__50536\,
            lcout => OPEN,
            ltout => \n13142_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9514_4_lut_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__48681\,
            in1 => \N__50759\,
            in2 => \N__43026\,
            in3 => \N__43023\,
            lcout => n149,
            ltout => \n149_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i19_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__42994\,
            in1 => \N__42948\,
            in2 => \N__43014\,
            in3 => \N__42933\,
            lcout => pin_out_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_190_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110000"
        )
    port map (
            in0 => \N__42978\,
            in1 => \N__43289\,
            in2 => \N__47527\,
            in3 => \N__42947\,
            lcout => n7326,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_887_i11_2_lut_4_lut_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__50345\,
            in1 => \N__48999\,
            in2 => \N__50567\,
            in3 => \N__50761\,
            lcout => n11_adj_734,
            ltout => \n11_adj_734_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_adj_241_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__49191\,
            in1 => \N__49141\,
            in2 => \N__42921\,
            in3 => \N__46992\,
            lcout => n36_adj_773,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Mux_35_i19_3_lut_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42898\,
            in1 => \N__42856\,
            in2 => \_gnd_net_\,
            in3 => \N__48996\,
            lcout => OPEN,
            ltout => \n19_adj_735_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9294_4_lut_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__48997\,
            in1 => \N__47323\,
            in2 => \N__43341\,
            in3 => \N__50343\,
            lcout => n13141,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_783_i11_2_lut_4_lut_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__50344\,
            in1 => \N__48998\,
            in2 => \N__50566\,
            in3 => \N__50760\,
            lcout => n11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_183_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__49923\,
            in1 => \N__49722\,
            in2 => \_gnd_net_\,
            in3 => \N__49516\,
            lcout => n1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_179_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010101010"
        )
    port map (
            in0 => \N__47518\,
            in1 => \N__43323\,
            in2 => \N__43299\,
            in3 => \N__43250\,
            lcout => OPEN,
            ltout => \n7310_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i15_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__43251\,
            in1 => \N__47869\,
            in2 => \N__43236\,
            in3 => \N__46488\,
            lcout => pin_out_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48440\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_i14_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111100000010"
        )
    port map (
            in0 => \N__49554\,
            in1 => \N__49956\,
            in2 => \N__49757\,
            in3 => \N__43149\,
            lcout => neopxl_color_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48440\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1617_3_lut_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__44113\,
            in1 => \_gnd_net_\,
            in2 => \N__43737\,
            in3 => \N__43710\,
            lcout => \nx.n2398\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1616_3_lut_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46047\,
            in2 => \N__46023\,
            in3 => \N__44109\,
            lcout => \nx.n2397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \neopxl_color_prev_i14_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43159\,
            lcout => neopxl_color_prev_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48444\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1619_3_lut_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43785\,
            in2 => \N__43815\,
            in3 => \N__44115\,
            lcout => \nx.n2400\,
            ltout => \nx.n2400_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.i15_4_lut_adj_62_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__43591\,
            in1 => \N__43615\,
            in2 => \N__43671\,
            in3 => \N__43668\,
            lcout => \nx.n35_adj_658\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1621_3_lut_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44114\,
            in2 => \N__43872\,
            in3 => \N__43894\,
            lcout => \nx.n2402\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_i1625_rep_47_3_lut_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43380\,
            in2 => \N__44128\,
            in3 => \N__43410\,
            lcout => \nx.n2406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_2_lut_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43572\,
            in2 => \_gnd_net_\,
            in3 => \N__43497\,
            lcout => \nx.n2377\,
            ltout => OPEN,
            carryin => \bfn_15_23_0_\,
            carryout => \nx.n10708\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_3_lut_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43494\,
            in3 => \N__43455\,
            lcout => \nx.n2376\,
            ltout => OPEN,
            carryin => \nx.n10708\,
            carryout => \nx.n10709\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_4_lut_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45677\,
            in2 => \N__43452\,
            in3 => \N__43413\,
            lcout => \nx.n2375\,
            ltout => OPEN,
            carryin => \nx.n10709\,
            carryout => \nx.n10710\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_5_lut_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45679\,
            in2 => \N__43409\,
            in3 => \N__43374\,
            lcout => \nx.n2374\,
            ltout => OPEN,
            carryin => \nx.n10710\,
            carryout => \nx.n10711\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_6_lut_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45678\,
            in2 => \N__43371\,
            in3 => \N__43989\,
            lcout => \nx.n2373\,
            ltout => OPEN,
            carryin => \nx.n10711\,
            carryout => \nx.n10712\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_7_lut_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45680\,
            in2 => \N__43985\,
            in3 => \N__43944\,
            lcout => \nx.n2372\,
            ltout => OPEN,
            carryin => \nx.n10712\,
            carryout => \nx.n10713\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_8_lut_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43940\,
            in2 => \N__45756\,
            in3 => \N__43902\,
            lcout => \nx.n2371\,
            ltout => OPEN,
            carryin => \nx.n10713\,
            carryout => \nx.n10714\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_9_lut_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45684\,
            in2 => \N__43898\,
            in3 => \N__43863\,
            lcout => \nx.n2370\,
            ltout => OPEN,
            carryin => \nx.n10714\,
            carryout => \nx.n10715\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_10_lut_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45414\,
            in2 => \N__43860\,
            in3 => \N__43818\,
            lcout => \nx.n2369\,
            ltout => OPEN,
            carryin => \bfn_15_24_0_\,
            carryout => \nx.n10716\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_11_lut_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45433\,
            in2 => \N__43811\,
            in3 => \N__43776\,
            lcout => \nx.n2368\,
            ltout => OPEN,
            carryin => \nx.n10716\,
            carryout => \nx.n10717\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_12_lut_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45415\,
            in2 => \N__43773\,
            in3 => \N__43740\,
            lcout => \nx.n2367\,
            ltout => OPEN,
            carryin => \nx.n10717\,
            carryout => \nx.n10718\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_13_lut_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45434\,
            in2 => \N__43733\,
            in3 => \N__43701\,
            lcout => \nx.n2366\,
            ltout => OPEN,
            carryin => \nx.n10718\,
            carryout => \nx.n10719\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_14_lut_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45416\,
            in2 => \N__46046\,
            in3 => \N__46011\,
            lcout => \nx.n2365\,
            ltout => OPEN,
            carryin => \nx.n10719\,
            carryout => \nx.n10720\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_15_lut_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45435\,
            in2 => \N__46007\,
            in3 => \N__45984\,
            lcout => \nx.n2364\,
            ltout => OPEN,
            carryin => \nx.n10720\,
            carryout => \nx.n10721\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_16_lut_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45417\,
            in2 => \N__45981\,
            in3 => \N__45948\,
            lcout => \nx.n2363\,
            ltout => OPEN,
            carryin => \nx.n10721\,
            carryout => \nx.n10722\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_17_lut_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45436\,
            in2 => \N__45945\,
            in3 => \N__45900\,
            lcout => \nx.n2362\,
            ltout => OPEN,
            carryin => \nx.n10722\,
            carryout => \nx.n10723\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_18_lut_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45411\,
            in2 => \N__45897\,
            in3 => \N__45855\,
            lcout => \nx.n2361\,
            ltout => OPEN,
            carryin => \bfn_15_25_0_\,
            carryout => \nx.n10724\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_19_lut_LC_15_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45432\,
            in2 => \N__45852\,
            in3 => \N__45813\,
            lcout => \nx.n2360\,
            ltout => OPEN,
            carryin => \nx.n10724\,
            carryout => \nx.n10725\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_20_lut_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45412\,
            in2 => \N__45805\,
            in3 => \N__45768\,
            lcout => \nx.n2359\,
            ltout => OPEN,
            carryin => \nx.n10725\,
            carryout => \nx.n10726\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nx.mod_5_add_1607_21_lut_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__45413\,
            in1 => \N__44148\,
            in2 => \N__44130\,
            in3 => \N__44013\,
            lcout => \nx.n2390\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i0_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46119\,
            in2 => \_gnd_net_\,
            in3 => \N__46113\,
            lcout => n26,
            ltout => OPEN,
            carryin => \bfn_15_26_0_\,
            carryout => n10548,
            clk => \N__48450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i1_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46110\,
            in2 => \_gnd_net_\,
            in3 => \N__46104\,
            lcout => n25,
            ltout => OPEN,
            carryin => n10548,
            carryout => n10549,
            clk => \N__48450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i2_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46101\,
            in2 => \_gnd_net_\,
            in3 => \N__46095\,
            lcout => n24,
            ltout => OPEN,
            carryin => n10549,
            carryout => n10550,
            clk => \N__48450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i3_LC_15_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46092\,
            in2 => \_gnd_net_\,
            in3 => \N__46086\,
            lcout => n23,
            ltout => OPEN,
            carryin => n10550,
            carryout => n10551,
            clk => \N__48450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i4_LC_15_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46083\,
            in2 => \_gnd_net_\,
            in3 => \N__46077\,
            lcout => n22,
            ltout => OPEN,
            carryin => n10551,
            carryout => n10552,
            clk => \N__48450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i5_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46074\,
            in2 => \_gnd_net_\,
            in3 => \N__46068\,
            lcout => n21_adj_737,
            ltout => OPEN,
            carryin => n10552,
            carryout => n10553,
            clk => \N__48450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i6_LC_15_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46065\,
            in2 => \_gnd_net_\,
            in3 => \N__46059\,
            lcout => n20,
            ltout => OPEN,
            carryin => n10553,
            carryout => n10554,
            clk => \N__48450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i7_LC_15_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46056\,
            in2 => \_gnd_net_\,
            in3 => \N__46050\,
            lcout => n19_adj_718,
            ltout => OPEN,
            carryin => n10554,
            carryout => n10555,
            clk => \N__48450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i8_LC_15_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46200\,
            in2 => \_gnd_net_\,
            in3 => \N__46194\,
            lcout => n18,
            ltout => OPEN,
            carryin => \bfn_15_27_0_\,
            carryout => n10556,
            clk => \N__48451\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i9_LC_15_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46191\,
            in2 => \_gnd_net_\,
            in3 => \N__46185\,
            lcout => n17,
            ltout => OPEN,
            carryin => n10556,
            carryout => n10557,
            clk => \N__48451\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i10_LC_15_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46182\,
            in2 => \_gnd_net_\,
            in3 => \N__46176\,
            lcout => n16,
            ltout => OPEN,
            carryin => n10557,
            carryout => n10558,
            clk => \N__48451\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i11_LC_15_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46173\,
            in2 => \_gnd_net_\,
            in3 => \N__46167\,
            lcout => n15_adj_759,
            ltout => OPEN,
            carryin => n10558,
            carryout => n10559,
            clk => \N__48451\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i12_LC_15_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46164\,
            in2 => \_gnd_net_\,
            in3 => \N__46158\,
            lcout => n14_adj_745,
            ltout => OPEN,
            carryin => n10559,
            carryout => n10560,
            clk => \N__48451\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i13_LC_15_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46155\,
            in2 => \_gnd_net_\,
            in3 => \N__46149\,
            lcout => n13,
            ltout => OPEN,
            carryin => n10560,
            carryout => n10561,
            clk => \N__48451\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i14_LC_15_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46146\,
            in2 => \_gnd_net_\,
            in3 => \N__46140\,
            lcout => n12,
            ltout => OPEN,
            carryin => n10561,
            carryout => n10562,
            clk => \N__48451\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i15_LC_15_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46137\,
            in2 => \_gnd_net_\,
            in3 => \N__46131\,
            lcout => n11_adj_758,
            ltout => OPEN,
            carryin => n10562,
            carryout => n10563,
            clk => \N__48451\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i16_LC_15_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46128\,
            in2 => \_gnd_net_\,
            in3 => \N__46122\,
            lcout => n10_adj_757,
            ltout => OPEN,
            carryin => \bfn_15_28_0_\,
            carryout => n10564,
            clk => \N__48452\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i17_LC_15_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46314\,
            in2 => \_gnd_net_\,
            in3 => \N__46308\,
            lcout => n9,
            ltout => OPEN,
            carryin => n10564,
            carryout => n10565,
            clk => \N__48452\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i18_LC_15_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46305\,
            in2 => \_gnd_net_\,
            in3 => \N__46299\,
            lcout => n8_adj_755,
            ltout => OPEN,
            carryin => n10565,
            carryout => n10566,
            clk => \N__48452\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i19_LC_15_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46296\,
            in2 => \_gnd_net_\,
            in3 => \N__46290\,
            lcout => n7,
            ltout => OPEN,
            carryin => n10566,
            carryout => n10567,
            clk => \N__48452\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i20_LC_15_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46287\,
            in2 => \_gnd_net_\,
            in3 => \N__46281\,
            lcout => n6_adj_756,
            ltout => OPEN,
            carryin => n10567,
            carryout => n10568,
            clk => \N__48452\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i21_LC_15_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46273\,
            in2 => \_gnd_net_\,
            in3 => \N__46260\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n10568,
            carryout => n10569,
            clk => \N__48452\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i22_LC_15_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46255\,
            in2 => \_gnd_net_\,
            in3 => \N__46242\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n10569,
            carryout => n10570,
            clk => \N__48452\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i23_LC_15_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46234\,
            in2 => \_gnd_net_\,
            in3 => \N__46221\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n10570,
            carryout => n10571,
            clk => \N__48452\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i24_LC_15_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46216\,
            in2 => \_gnd_net_\,
            in3 => \N__46203\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_15_29_0_\,
            carryout => n10572,
            clk => \N__48453\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_1105__i25_LC_15_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46352\,
            in2 => \_gnd_net_\,
            in3 => \N__46356\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48453\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1103__i0_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__46578\,
            in1 => \N__49412\,
            in2 => \_gnd_net_\,
            in3 => \N__46341\,
            lcout => counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48441\,
            ce => \N__47530\,
            sr => \_gnd_net_\
        );

    \counter_1103_add_4_2_lut_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47570\,
            in2 => \N__47630\,
            in3 => \N__46335\,
            lcout => n45,
            ltout => OPEN,
            carryin => \bfn_16_15_0_\,
            carryout => n10510,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1103__i1_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__46567\,
            in1 => \N__48177\,
            in2 => \N__46928\,
            in3 => \N__46332\,
            lcout => counter_1,
            ltout => OPEN,
            carryin => n10510,
            carryout => n10511,
            clk => \N__48438\,
            ce => \N__47538\,
            sr => \_gnd_net_\
        );

    \counter_1103__i2_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__46579\,
            in1 => \N__46878\,
            in2 => \N__47556\,
            in3 => \N__46329\,
            lcout => counter_2,
            ltout => OPEN,
            carryin => n10511,
            carryout => n10512,
            clk => \N__48438\,
            ce => \N__47538\,
            sr => \_gnd_net_\
        );

    \counter_1103__i3_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__46568\,
            in1 => \N__47598\,
            in2 => \N__46929\,
            in3 => \N__46326\,
            lcout => counter_3,
            ltout => OPEN,
            carryin => n10512,
            carryout => n10513,
            clk => \N__48438\,
            ce => \N__47538\,
            sr => \_gnd_net_\
        );

    \counter_1103__i4_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__46580\,
            in1 => \N__46882\,
            in2 => \N__47586\,
            in3 => \N__46323\,
            lcout => counter_4,
            ltout => OPEN,
            carryin => n10513,
            carryout => n10514,
            clk => \N__48438\,
            ce => \N__47538\,
            sr => \_gnd_net_\
        );

    \counter_1103__i5_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__46569\,
            in1 => \N__48162\,
            in2 => \N__46930\,
            in3 => \N__46320\,
            lcout => counter_5,
            ltout => OPEN,
            carryin => n10514,
            carryout => n10515,
            clk => \N__48438\,
            ce => \N__47538\,
            sr => \_gnd_net_\
        );

    \counter_1103__i6_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__46581\,
            in1 => \N__46886\,
            in2 => \N__47172\,
            in3 => \N__46317\,
            lcout => counter_6,
            ltout => OPEN,
            carryin => n10515,
            carryout => n10516,
            clk => \N__48438\,
            ce => \N__47538\,
            sr => \_gnd_net_\
        );

    \counter_1103__i7_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__46570\,
            in1 => \N__47229\,
            in2 => \N__46931\,
            in3 => \N__46986\,
            lcout => counter_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48438\,
            ce => \N__47538\,
            sr => \_gnd_net_\
        );

    \i3_3_lut_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__47156\,
            in1 => \N__49999\,
            in2 => \_gnd_net_\,
            in3 => \N__48132\,
            lcout => OPEN,
            ltout => \n8_adj_763_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9579_4_lut_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__47105\,
            in1 => \N__47225\,
            in2 => \N__46983\,
            in3 => \N__49526\,
            lcout => n7223,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_adj_199_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__46787\,
            in1 => \N__50125\,
            in2 => \_gnd_net_\,
            in3 => \N__46679\,
            lcout => n12208,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state_7__I_0_205_i16_1_lut_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49406\,
            lcout => \current_pin_7__N_155\,
            ltout => \current_pin_7__N_155_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2960_3_lut_4_lut_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__46786\,
            in1 => \N__46744\,
            in2 => \N__46695\,
            in3 => \N__46678\,
            lcout => n6180,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_adj_220_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__49527\,
            in1 => \N__50000\,
            in2 => \_gnd_net_\,
            in3 => \N__49807\,
            lcout => n6971,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4169_2_lut_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49410\,
            in2 => \_gnd_net_\,
            in3 => \N__48233\,
            lcout => n7401,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4263_4_lut_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011110100"
        )
    port map (
            in0 => \N__46542\,
            in1 => \N__47528\,
            in2 => \N__47324\,
            in3 => \N__46475\,
            lcout => OPEN,
            ltout => \n7500_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pin_output_i0_i22_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110000"
        )
    port map (
            in0 => \N__47529\,
            in1 => \N__47346\,
            in2 => \N__47340\,
            in3 => \N__49411\,
            lcout => pin_out_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48427\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_233_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001011"
        )
    port map (
            in0 => \N__47294\,
            in1 => \N__50315\,
            in2 => \N__49413\,
            in3 => \N__48955\,
            lcout => n4_adj_778,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_216_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__48474\,
            in1 => \N__48519\,
            in2 => \_gnd_net_\,
            in3 => \N__48553\,
            lcout => n7142,
            ltout => \n7142_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_234_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__47241\,
            in3 => \N__48645\,
            lcout => n14_adj_717,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state__i2_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__47237\,
            in1 => \N__50016\,
            in2 => \N__47180\,
            in3 => \N__48150\,
            lcout => state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48436\,
            ce => \N__50820\,
            sr => \N__48213\
        );

    \i9575_2_lut_3_lut_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__50015\,
            in1 => \N__49751\,
            in2 => \_gnd_net_\,
            in3 => \N__49489\,
            lcout => n73,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_239_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__49003\,
            in1 => \N__47780\,
            in2 => \N__50338\,
            in3 => \N__50611\,
            lcout => OPEN,
            ltout => \n12123_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19_4_lut_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__47088\,
            in1 => \N__47043\,
            in2 => \N__47037\,
            in3 => \N__49056\,
            lcout => n48_adj_771,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i380_3_lut_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__47022\,
            in1 => \N__47742\,
            in2 => \_gnd_net_\,
            in3 => \N__47779\,
            lcout => n2313,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9297_4_lut_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__48717\,
            in1 => \N__50287\,
            in2 => \N__47927\,
            in3 => \N__49001\,
            lcout => OPEN,
            ltout => \n13144_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9442_4_lut_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__50752\,
            in1 => \N__49152\,
            in2 => \N__47811\,
            in3 => \N__50537\,
            lcout => n13279,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_791_i15_4_lut_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__47778\,
            in1 => \N__50288\,
            in2 => \N__50615\,
            in3 => \N__49002\,
            lcout => n15_adj_750,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_243_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110001111"
        )
    port map (
            in0 => \N__47741\,
            in1 => \N__48747\,
            in2 => \N__49772\,
            in3 => \N__49143\,
            lcout => n30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_adj_242_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__47718\,
            in1 => \N__49517\,
            in2 => \_gnd_net_\,
            in3 => \N__47685\,
            lcout => n6_adj_766,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \state__i1_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010001000100"
        )
    port map (
            in0 => \N__49749\,
            in1 => \N__49955\,
            in2 => \N__47664\,
            in3 => \N__47643\,
            lcout => state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48442\,
            ce => \N__50816\,
            sr => \N__50787\
        );

    \state__i0_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__49954\,
            in1 => \N__49750\,
            in2 => \_gnd_net_\,
            in3 => \N__47631\,
            lcout => state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48442\,
            ce => \N__50816\,
            sr => \N__50787\
        );

    \i4_4_lut_adj_246_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47597\,
            in1 => \N__47582\,
            in2 => \N__47571\,
            in3 => \N__47549\,
            lcout => OPEN,
            ltout => \n10_adj_762_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_3_lut_adj_247_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48176\,
            in2 => \N__48165\,
            in3 => \N__48161\,
            lcout => n18_adj_742,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_895_i11_2_lut_4_lut_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__50499\,
            in1 => \N__48913\,
            in2 => \N__50332\,
            in3 => \N__50753\,
            lcout => n11_adj_739,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__50492\,
            in1 => \N__48845\,
            in2 => \N__50754\,
            in3 => \N__48646\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9317_3_lut_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48843\,
            in1 => \N__48077\,
            in2 => \_gnd_net_\,
            in3 => \N__48038\,
            lcout => OPEN,
            ltout => \n13164_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_pin_1__bdd_4_lut_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__50491\,
            in1 => \N__50204\,
            in2 => \N__48009\,
            in3 => \N__47820\,
            lcout => n13468,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_280_i6_2_lut_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50205\,
            in2 => \_gnd_net_\,
            in3 => \N__48844\,
            lcout => n6_adj_748,
            ltout => \n6_adj_748_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i488_4_lut_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__47928\,
            in1 => \N__50595\,
            in2 => \N__47886\,
            in3 => \N__49146\,
            lcout => n2421,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9318_3_lut_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48842\,
            in1 => \N__47883\,
            in2 => \_gnd_net_\,
            in3 => \N__47843\,
            lcout => n13165,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_pin_i0_i0_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48894\,
            in2 => \_gnd_net_\,
            in3 => \N__47814\,
            lcout => current_pin_0,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => n10384,
            clk => \N__48433\,
            ce => \N__48234\,
            sr => \N__48222\
        );

    \current_pin_i0_i1_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50316\,
            in2 => \_gnd_net_\,
            in3 => \N__48711\,
            lcout => current_pin_1,
            ltout => OPEN,
            carryin => n10384,
            carryout => n10385,
            clk => \N__48433\,
            ce => \N__48234\,
            sr => \N__48222\
        );

    \current_pin_i0_i2_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50490\,
            in2 => \_gnd_net_\,
            in3 => \N__48708\,
            lcout => current_pin_2,
            ltout => OPEN,
            carryin => n10385,
            carryout => n10386,
            clk => \N__48433\,
            ce => \N__48234\,
            sr => \N__48222\
        );

    \current_pin_i0_i3_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50712\,
            in2 => \_gnd_net_\,
            in3 => \N__48705\,
            lcout => current_pin_3,
            ltout => OPEN,
            carryin => n10386,
            carryout => n10387,
            clk => \N__48433\,
            ce => \N__48234\,
            sr => \N__48222\
        );

    \current_pin_i0_i4_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48647\,
            in2 => \_gnd_net_\,
            in3 => \N__48576\,
            lcout => current_pin_4,
            ltout => OPEN,
            carryin => n10387,
            carryout => n10388,
            clk => \N__48433\,
            ce => \N__48234\,
            sr => \N__48222\
        );

    \current_pin_i0_i5_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48559\,
            in2 => \_gnd_net_\,
            in3 => \N__48537\,
            lcout => current_pin_5,
            ltout => OPEN,
            carryin => n10388,
            carryout => n10389,
            clk => \N__48433\,
            ce => \N__48234\,
            sr => \N__48222\
        );

    \current_pin_i0_i6_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48526\,
            in2 => \_gnd_net_\,
            in3 => \N__48498\,
            lcout => current_pin_6,
            ltout => OPEN,
            carryin => n10389,
            carryout => n10390,
            clk => \N__48433\,
            ce => \N__48234\,
            sr => \N__48222\
        );

    \current_pin_i0_i7_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48481\,
            in2 => \_gnd_net_\,
            in3 => \N__48495\,
            lcout => current_pin_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48433\,
            ce => \N__48234\,
            sr => \N__48222\
        );

    \i4172_2_lut_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__49752\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50815\,
            lcout => n7409,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13_4_lut_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001000"
        )
    port map (
            in0 => \N__49145\,
            in1 => \N__49290\,
            in2 => \N__48201\,
            in3 => \N__49368\,
            lcout => n42,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_4_lut_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__49263\,
            in1 => \N__49359\,
            in2 => \N__49350\,
            in3 => \N__49144\,
            lcout => OPEN,
            ltout => \n40_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i25_4_lut_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__49323\,
            in1 => \N__49311\,
            in2 => \N__49305\,
            in3 => \N__49302\,
            lcout => n54_adj_768,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_pin_0__bdd_4_lut_9619_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__49283\,
            in1 => \N__50284\,
            in2 => \N__49259\,
            in3 => \N__48968\,
            lcout => OPEN,
            ltout => \n13444_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n13444_bdd_4_lut_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__50285\,
            in1 => \N__49226\,
            in2 => \N__49194\,
            in3 => \N__49187\,
            lcout => n13447,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_919_i15_4_lut_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__49142\,
            in1 => \N__50286\,
            in2 => \N__50607\,
            in3 => \N__48969\,
            lcout => OPEN,
            ltout => \n15_adj_749_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_adj_240_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__48774\,
            in1 => \N__49095\,
            in2 => \N__49065\,
            in3 => \N__49062\,
            lcout => n37,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Mux_34_i19_3_lut_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48967\,
            in1 => \N__48773\,
            in2 => \_gnd_net_\,
            in3 => \N__48746\,
            lcout => n19_adj_715,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9261_4_lut_4_lut_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100010101000"
        )
    port map (
            in0 => \N__49524\,
            in1 => \N__49941\,
            in2 => \N__49796\,
            in3 => \N__50859\,
            lcout => OPEN,
            ltout => \n13037_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_244_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__50853\,
            in1 => \N__50844\,
            in2 => \N__50832\,
            in3 => \N__50829\,
            lcout => n7249,
            ltout => \n7249_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4158_2_lut_4_lut_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__49525\,
            in1 => \N__49942\,
            in2 => \N__50790\,
            in3 => \N__49697\,
            lcout => n7395,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_927_i10_2_lut_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50687\,
            in2 => \_gnd_net_\,
            in3 => \N__50444\,
            lcout => n10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6234_2_lut_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__50445\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50256\,
            lcout => n9456,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_218_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__50014\,
            in1 => \N__49773\,
            in2 => \_gnd_net_\,
            in3 => \N__49509\,
            lcout => n15_adj_721,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
