// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Wed Apr  7 16:39:04 2021
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(41[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(41[16:24])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, 
        INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(54[12:14])
    
    wire reset;
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(57[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, GHB, GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(103[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(104[21:25])
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(139[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(140[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(149[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(246[21:45])
    
    wire n1761;
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(248[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(249[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(250[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(251[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(252[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(254[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(255[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(256[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(257[22:30])
    wire [15:0]current;   // verilog/TinyFPGA_B.v(258[22:29])
    wire [15:0]current_limit;   // verilog/TinyFPGA_B.v(259[22:35])
    wire [31:0]baudrate;   // verilog/TinyFPGA_B.v(261[15:23])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(290[22:33])
    
    wire data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(360[11:24])
    
    wire n55388;
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(368[15:20])
    
    wire pwm_setpoint_23__N_207, n11590, n11592, n11594, n11596, n11598, 
        n11600, n11602, n11604, n11606, n11608, n11610, n11612, 
        n11614, n11616, n11618, n11620, n55296, n260, n11628, 
        n11626, n294, n298, n299, n300, n301, n302, n303, n304, 
        n305, n306, n307, n308, n309;
    wire [23:0]pwm_setpoint_23__N_3;
    wire [7:0]commutation_state_7__N_208;
    
    wire commutation_state_7__N_216;
    wire [7:0]commutation_state_7__N_27;
    
    wire n29437, n1763, n1765, n1767, n1769;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(245[11:28])
    
    wire GHA_N_355, GLA_N_372, GHB_N_377, GLB_N_386, GHC_N_391, GLC_N_400, 
        dti_N_404, n38194, n29434, n38221, n29431, RX_N_2, n1759, 
        n1757, n1755, n1753, n1751, n1749;
    wire [31:0]motor_state_23__N_91;
    wire [38:0]encoder1_position_scaled_23__N_43;
    wire [23:0]displacement_23__N_67;
    
    wire n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, 
        n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, 
        n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, 
        n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, 
        read_N_409, n1325, n62, n25, n23, n21, n1800;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(247[11:28])
    wire [10:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [10:0]t0;   // verilog/neopixel.v(10[12:14])
    wire [1:0]state;   // verilog/neopixel.v(19[11:16])
    wire [4:0]bit_ctr;   // verilog/neopixel.v(20[11:18])
    
    wire n55412, n8, n25_adj_5690, n24, n23_adj_5691, n22, n21_adj_5692, 
        n20, n19, n29428, n29424, n29421, n19_adj_5693, n17, n16, 
        n15, n13, n12, n11, n10, n9, n17_adj_5694, n2829, n16_adj_5695, 
        n38223, n15_adj_5696, n14, n13_adj_5697, n2, n14_adj_5698, 
        n15_adj_5699, n16_adj_5700, n17_adj_5701, n18, n19_adj_5702, 
        n20_adj_5703, n21_adj_5704, n22_adj_5705, n23_adj_5706, n24_adj_5707, 
        n25_adj_5708, n24_adj_5709, n33791, n29418, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(94[13:20])
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(99[12:25])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[3] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[1] ;   // verilog/coms.v(100[12:26])
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(100[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(105[12:33])
    
    wire tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(115[11:16])
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire \FRAME_MATCHER.rx_data_ready_prev , n4938, n4937, n4936, n4916, 
        n4915, n4917, n4918, n4919, n4920, n4921, n4922, n4923, 
        n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, 
        n4932, n4933, n4934, n4935, n55391, n3484, n2882, n25141, 
        n3, n38279, n38316, n29415, n39972, n31, n55533, n39937, 
        n9_adj_5710, n39919, n38386, n53, n55681, n55624, n57036, 
        n49097, n49096, n49095, n48277, n48276, n49094, n49093, 
        n49092, n49091, n48275, n48274, n48583, n48582, n48260, 
        n48581, n48580, n48259, n48579, n48273, n48578, n48577, 
        n48576, n32987, n55390, n55295, n48575, n48574, n48573, 
        n48572, n48571, n48570, n48569, n48568, n48567, n48566, 
        n48565, n25895, n48564, n48563, n48562, n48561, n48560, 
        n48258, n48559, n48558, n66702, n48557, n48556, n48555, 
        n48554, n48553, n48552, n48551, n48550, n48549, n48548, 
        n48272, n48547, n48546, n48271, n28910, n8_adj_5711, Kp_23__N_748, 
        n48545, n48544, Kp_23__N_875, n48270, n15_adj_5712, n8_adj_5713, 
        n48269, n65098, n29409, n38638, n29406, n29403, n29400, 
        \FRAME_MATCHER.i_31__N_2509 , n73, n29397, n20722, n29394, 
        n29392, n29389, n29384, n29381, n29378, n29374, n29371, 
        n29368, n29365, n29362, n29359, n29356, n29353, n29349, 
        n29346, n29343, n29316, n29313, n29309, n29306, n29303, 
        n29300, n29297, n29294, n29291, n29288, n29285, n66244, 
        n29282, n29278, n29275, n29272, n29269, n29266, n29263, 
        n29258, n29255, n29252, n29249, n29246, n29243, n15553, 
        n29176, n48257, n29156, n29155, n29154, n29153, n29152, 
        n29151, n29150, n29149, n29148, n29147, n29146, n29145, 
        n29144, n29143, n29142, n29141, n29140, n29139, n29138, 
        n29137, n29136, n29135, n29134, n29133, n29132, n29131, 
        n29130, n29129, n29128, n29127, n29126, n29125, n29124, 
        n29123, n29114, n29113, n29112, n29111, n29110, n29109, 
        n29108, n29107, n29106, n29105, n29104, n29103, n29102, 
        n29101, n29100, n29099, n29098, n29097, n29096, n29064, 
        n29063, n29062, n29061, n29060, n29051, n29048, n29045, 
        n65449, n29042, n29033, n29030, n29024, n29015, n29012, 
        n29009, n29006, n29003, n29000, n28997, n28994, n28991, 
        n7, n6, n5, n4, n24_adj_5714, n19_adj_5715, n17_adj_5716, 
        n16_adj_5717, n15_adj_5718, n13_adj_5719, n11_adj_5720, n9_adj_5721, 
        n8_adj_5722, n7_adj_5723, n6_adj_5724, n5_adj_5725, n4_adj_5726, 
        n30, n65225, n23_adj_5727, n21_adj_5728, n19_adj_5729, n17_adj_5730, 
        n16_adj_5731, n15_adj_5732, n13_adj_5733, n11_adj_5734, n10_adj_5735, 
        n9_adj_5736, n8_adj_5737, n7_adj_5738, n6_adj_5739, n4_adj_5740, 
        n48256, n66231, n55294, n55293, n55292, n55291, n55290, 
        n55243, n55385, n55289, n55386, n15_adj_5741, n55288, n55287, 
        n55286, n55285, n55284, n55283, n4_adj_5742, n4_adj_5743, 
        n66201, n4_adj_5744, n24971, n10_adj_5745, n28988, control_update;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(36[23:31])
    
    wire n105, n11588, n55282, n336, n337, n338, n339, n340, 
        n341, n342, n343, n344, n345, n346, n347, n348, n349, 
        n350, n351, n352, n353, n354, n355, n356, n357, n358, 
        n359, n24981, n7064, n5228, n5225, n3173, n22318, n5_adj_5746, 
        n11_adj_5747, n28982;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev, b_prev, debounce_cnt_N_3833, position_31__N_3836, n65457, 
        n22471, n15_adj_5748;
    wire [1:0]a_new_adj_5885;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [1:0]b_new_adj_5886;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire a_prev_adj_5751, b_prev_adj_5752, debounce_cnt_N_3833_adj_5753, 
        position_31__N_3836_adj_5754, n60219, n12_adj_5755, n11_adj_5756, 
        n10_adj_5757, n4_adj_5758, n3_adj_5759, n2_adj_5760;
    wire [7:0]data_adj_5899;   // verilog/eeprom.v(23[12:16])
    wire [7:0]state_7__N_3918;
    
    wire n66672, n66669, n28976, n5_adj_5761, n55281, n6911, n29826, 
        n29825, n29824, n29823, n24969, n66010, n29822, n29821, 
        n29820, n29819, n29818, n29817, n29816;
    wire [15:0]data_adj_5906;   // verilog/tli4970.v(27[14:18])
    
    wire n29815, n66002, n49510, n29814, n29812, n29811, n29810, 
        n29809, n29808, n49509, n49508, n29806, n49507, n49506, 
        n49505, n15_adj_5770, n29778, n29777, n55985, n49504, n5_adj_5771, 
        n29776, n29775, n29774, n29773, n29772, n29771, n49503, 
        n11622, n11624, n49502, n29770, n29769, n29768, n29767, 
        state_7__N_4319, n29766, n49501, n28967, n9_adj_5772, n8_adj_5773, 
        n49500, n7_adj_5774, n6_adj_5775, n5_adj_5776, n29765, n29764, 
        n29763, n29762, n29761, n29760, n29759, n29758, n29757, 
        n29754, n24966, n49499, r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(33[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(37[17:26])
    
    wire n49498, n57520, n49497, n49496;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n66654, n49495, n28964;
    wire [2:0]r_SM_Main_2__N_3446;
    wire [2:0]r_SM_Main_adj_5922;   // verilog/uart_tx.v(32[16:25])
    wire [8:0]r_Clock_Count_adj_5923;   // verilog/uart_tx.v(33[16:29])
    wire [2:0]r_Bit_Index_adj_5924;   // verilog/uart_tx.v(34[16:27])
    wire [2:0]r_SM_Main_2__N_3545;
    
    wire o_Tx_Serial_N_3598, n49494, n48268, n48267, n49493;
    wire [7:0]state_adj_5935;   // verilog/i2c_controller.v(33[12:17])
    
    wire n48511, enable_slow_N_4213, n29677, n29676, n29674, n28961, 
        n29673, n48510, n48509, n29671, n8_adj_5789, n29670;
    wire [7:0]state_7__N_4110;
    
    wire n29669, n29668, n29667, n29666, n29665, n29664, n29662, 
        n29661, n6715, n29660, n29659, n29658, n29657, n29656, 
        n48508, n29655, n29654, n48507, n48506, n29650, n29649;
    wire [7:0]state_7__N_4126;
    
    wire n29648, n29647, n29646, n29645, n29644, n29643, n29642, 
        n29640, n29638, n29637, n29636, n29635, n29634, n29633, 
        n29632, n48505, n48504, n58374, n48503, n48502, n28958, 
        n28952, n48501, n48500, n48499, n55280, n55279, n55403, 
        n55278, n55277, n27460, n38711, n55401, n55276, n28729, 
        n55400, n13260, n55381, n55275, n55402, n27441, n55274, 
        n55273, n29600, n55272, n55271, n55270, n21_adj_5790, n25_adj_5791, 
        n36, n40, n48266, n55380, n55398, n67455, n55269, n28721, 
        n55268, n55382, n55242, n55396, n29596, n55383, n55267, 
        n55394, n55266, n55265, n55264, n55263, n55393, n28713, 
        n55410, n55262, n13254, n48265, n65917, n38266, n38659, 
        n48264, n48255, n1, n28711, n57999, n48263, n29592, n55297, 
        n13241, n24804, n65484, n55411, n55261, n13255, n48254, 
        n66651, n15543, n55298, n38328, n64560, n13242, n13256, 
        n65816, n65815, n66101, n9_adj_5792, n13243, n13249, n20_adj_5793, 
        n65672, n18_adj_5794, n16_adj_5795, n65671, n13257, n48429, 
        n48428, n24633, n48427, n48426, n15542, n15544, n15551, 
        n48425, n48424, n29589, n48423, n48422, n13244, n13250, 
        n48421, n48420, n25095, n13258, n55260, n29586, n55153, 
        n7_adj_5796, n13245, n13251, n15552, n65522, n13259, n26439, 
        n51433, n65526, n15541, n15545, n25100, n55259, n55258, 
        n55408, n22369, n28706, n55257, n55392, n55407, n27321, 
        n4_adj_5797, n6_adj_5798, n8_adj_5799, n9_adj_5800, n11_adj_5801, 
        n13_adj_5802, n14_adj_5803, n15_adj_5804, n4_adj_5805, n6_adj_5806, 
        n8_adj_5807, n9_adj_5808, n27315, n35729, n27312, n54695, 
        n27308, n48419, n48418, n29582, n55409, n6_adj_5809, n27290, 
        n29581, n38, n39, n40_adj_5810, n41, n42, n43, n44, 
        n45, n28949, n28946, n55406, n13247, n13253, n55256, n28703, 
        n55405, n29580, n15546, n15540, n66009, n27260, n29578, 
        n55302, n29577, n29576, n55255, n29575, n29574, n55254, 
        n55253, n55252, n55251, n27236, n55397, n28696, n55300, 
        n55399, n55250, n55249, n55299, n51161, n51197, n55419, 
        n55418, n55417, n55416, n55415, n55414, n55248, n55379, 
        n55247, n55303, n55246, n55378, n28689, n55304, n28688, 
        n55377, n55245, n55376, n55244, n55375, n55455, n55374, 
        n55454, n55373, n55453, n55372, n55452, n55371, n55451, 
        n55370, n28680, n55369, n55456, n55368, n55446, n55367, 
        n55447, n55366, n55448, n55365, n55449, n55364, n55450, 
        n55363, n55444, n55362, n28672, n55361, n55360, n55445, 
        n55359, n55358, n55357, n55356, n55355, n55354, n55353, 
        n55352, n55351, n55350, n55349, n55348, n55989, n55347, 
        n55346, n55345, n55344, n55343, n55342, n55341, n55340, 
        n55339, n55338, n55337, n55336, n55335, n55334, n55333, 
        n55332, n28642, n55331, n55330, n51296, n55329, n55328, 
        n56165, n55327, n55306, n55326, n55325, n55324, n55323, 
        n55322, n55321, n55320, n55319, n55305, n55318, n28611, 
        n55317, n55316, n55315, n55314, n55648, n55313, n55312, 
        n55311, n65523, n55310, n55309, n55308, n27939, n27934, 
        n27932, n27929, n27926, n55151, n55184, n55152, n55149, 
        n27906, n27904, n27902, n27900, n27898, n28348, n25803, 
        n48417, n48416, n48415, n35156, n55413, n55301, n15554, 
        n55307, n55395, n15547, n15539, n65123, n15555, n15548, 
        n48414, n15538, n48413, n48412, n9941, n9939, n48411, 
        n54697, n27212, n48410, n66618, n66615, n3_adj_5811, n48409, 
        n48408, n48407, n65222, n33833, n65221, n29558, n29555, 
        n29552, n29549, n29546, n25941, n25933, n48262, n28940, 
        n28939, n28938, n28937, n63538, n29512, n29509, n51232, 
        n29506, n29499, n29496, n28927, n29493, n29487, n37097, 
        n25133, n37113, n29484, n29481, n29477, n29468, n76, n15549, 
        n28925, n28923, n28922, n28921, n29440, n25110, n25494, 
        n13252, n15550, n13246, n15537, n59906, n21266, n21262, 
        n58172, n55404, n10_adj_5812, n55775, n55387, n50377, n50591, 
        n50927, n51425, n48375, n63490, n48374, n48373, n57982, 
        n48372, n48371, n55884, n65851, n50264, n55181, n50260, 
        n67005, n48261, n66999, n64508, n66993, n66987, n66981, 
        n66975, n11586, n48370, n48369, n48368, n48367, n48366, 
        n48365, n48364, n48363, n48362, n48361, n48360, n48359, 
        n48358, n48357, n48356, n48355, n50946, n48354, n25490, 
        n48353, n25130, n25705, n25108, n55389, n48283, n48282, 
        n50183, n55384, n66969, n13248, n63461, n64582, n27513, 
        n63426, n48281, n66963, n63399, n37128, n63397, n60054, 
        n63392, n64439, n55526, n78, n63388, n67, n28912, n48280, 
        n48253, n38695, n48279, n48278, n66957, n66951, n64425, 
        n66945, n64415, n66939, n64310, n64308, n14_adj_5813, n10_adj_5814, 
        n64298, n66933, n65151, n58982, n56368, n56366, n65159, 
        n58976, n65167, n58970, n58964, n58958, n66927, n58952, 
        n6_adj_5815, n18_adj_5816, n17_adj_5817, n16_adj_5818, n14_adj_5819, 
        n12_adj_5820, n58946, n58940, n66200, n58934, n56301, n15_adj_5821, 
        n14_adj_5822, n58932, n66921, n58928, n56281, n58922, n8_adj_5823, 
        n7_adj_5824, n6_adj_5825, n58916, n17_adj_5826, n25_adj_5827, 
        n53719, n24_adj_5828, n58910, n58904, n29, n66915, n27, 
        n4_adj_5829, n58898, n23_adj_5830, n58896, n14_adj_5831, n58892, 
        n10_adj_5832, n53805, n58886, n64008, n58880, n58874, n58868, 
        n4_adj_5833, n58862, n58312, n58856, n58850, n63988, n63986, 
        n58844, n65778, n66909, n56024, n55587, n55655, n55668, 
        n56050, n66903, n66102, n55766, n60056, n60055, n55241, 
        n56109, n6_adj_5834, n63151, n56183, n55443, n55524, n56059, 
        n56201, n63134, n66897, n56062, n58029, n58026, n63131, 
        n63124, n63121, n56162, n66891, n57376, n57716, n56231, 
        n4_adj_5835, n4_adj_5836, n10_adj_5837, n6_adj_5838, n4_adj_5839, 
        n66714, n12_adj_5840, n5_adj_5841, n56120, n66253, n58618, 
        n58612, n58606, n58600, n55952, n58594, n63020, n65756, 
        n6_adj_5842, n57943, n54733, n60225, n60222, n60220, n58502, 
        n58462, n62960, n23_adj_5843, n66864, n58452, n56216, n58202, 
        n62948, n66861, n66097, n14_adj_5844, n13_adj_5845, n62934, 
        n7_adj_5846;
    
    VCC i2 (.Y(VCC_net));
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1 */ ;   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1 */ ;   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(clk16MHz), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(151[9] 230[5])
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(current[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_5707));   // verilog/TinyFPGA_B.v(129[16:24])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_DFF dir_183 (.Q(dir), .C(clk16MHz), .D(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFFE dti_185 (.Q(dti), .C(clk16MHz), .E(n27212), .D(dti_N_404));   // verilog/TinyFPGA_B.v(151[9] 230[5])
    SB_LUT4 i13298_3_lut (.I0(ID[3]), .I1(data_adj_5899[3]), .I2(n55524), 
            .I3(GND_net), .O(n29143));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13298_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[2]), .C(clk16MHz), 
           .D(encoder0_position[0]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(clk16MHz), 
           .D(encoder1_position[0]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4126[3])) /* synthesis syn_instantiated=1 */ ;   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk16MHz), .D(displacement_23__N_67[0]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1 */ ;   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.clk16MHz(clk16MHz), .bit_ctr({Open_0, 
            Open_1, Open_2, bit_ctr[1:0]}), .GND_net(GND_net), .state({state}), 
            .n3173(n3173), .neopxl_color({neopxl_color}), .t0({t0}), .n23(n23_adj_5843), 
            .n38711(n38711), .timer({timer}), .n35156(n35156), .n27441(n27441), 
            .VCC_net(VCC_net), .n29176(n29176), .n5(n5_adj_5841), .n29155(n29155), 
            .n29154(n29154), .n29151(n29151), .n29150(n29150), .n29149(n29149), 
            .n29148(n29148), .n29147(n29147), .n29146(n29146), .n29145(n29145), 
            .n29144(n29144), .NEOPXL_c(NEOPXL_c), .n28939(n28939), .\data_in_frame[4][2] (\data_in_frame[4] [2]), 
            .\data_in_frame[4][3] (\data_in_frame[4] [3]), .n56059(n56059), 
            .\data_in_frame[1][6] (\data_in_frame[1] [6]), .\data_in_frame[1][7] (\data_in_frame[1] [7]), 
            .n55668(n55668), .n56216(n56216), .n25933(n25933), .Kp_23__N_875(Kp_23__N_875), 
            .\data_out_frame[23][2] (\data_out_frame[23] [2]), .\data_out_frame[23][3] (\data_out_frame[23] [3]), 
            .n55952(n55952), .\data_out_frame[24][7] (\data_out_frame[24] [7]), 
            .n50377(n50377), .n56165(n56165), .\rx_data[3] (rx_data[3]), 
            .n27900(n27900), .n28964(n28964), .n22369(n22369), .n29658(n29658), 
            .n29659(n29659), .LED_c(LED_c), .n24633(n24633), .\data_out_frame[21][0] (\data_out_frame[21] [0]), 
            .n56162(n56162), .\data_in_frame[2][0] (\data_in_frame[2] [0])) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(59[24] 65[2])
    SB_LUT4 i13299_3_lut (.I0(t0[10]), .I1(timer[10]), .I2(n3173), .I3(GND_net), 
            .O(n29144));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13300_3_lut (.I0(t0[9]), .I1(timer[9]), .I2(n3173), .I3(GND_net), 
            .O(n29145));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13301_3_lut (.I0(t0[8]), .I1(timer[8]), .I2(n3173), .I3(GND_net), 
            .O(n29146));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13302_3_lut (.I0(t0[7]), .I1(timer[7]), .I2(n3173), .I3(GND_net), 
            .O(n29147));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13303_3_lut (.I0(t0[6]), .I1(timer[6]), .I2(n3173), .I3(GND_net), 
            .O(n29148));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13303_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n48408), .I0(encoder0_position_scaled[2]), 
            .I1(n23_adj_5691), .CO(n48409));
    SB_LUT4 i13304_3_lut (.I0(t0[5]), .I1(timer[5]), .I2(n3173), .I3(GND_net), 
            .O(n29149));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24), .I3(n48407), .O(displacement_23__N_67[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13305_3_lut (.I0(t0[4]), .I1(timer[4]), .I2(n3173), .I3(GND_net), 
            .O(n29150));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13667_3_lut (.I0(\data_in_frame[21] [5]), .I1(rx_data[5]), 
            .I2(n27934), .I3(GND_net), .O(n29512));   // verilog/coms.v(130[12] 305[6])
    defparam i13667_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13664_3_lut (.I0(\data_in_frame[21] [4]), .I1(rx_data[4]), 
            .I2(n27934), .I3(GND_net), .O(n29509));   // verilog/coms.v(130[12] 305[6])
    defparam i13664_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13661_3_lut (.I0(\data_in_frame[21] [3]), .I1(rx_data[3]), 
            .I2(n27934), .I3(GND_net), .O(n29506));   // verilog/coms.v(130[12] 305[6])
    defparam i13661_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13654_3_lut (.I0(\data_in_frame[21] [2]), .I1(rx_data[2]), 
            .I2(n27934), .I3(GND_net), .O(n29499));   // verilog/coms.v(130[12] 305[6])
    defparam i13654_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13651_3_lut (.I0(\data_in_frame[21] [1]), .I1(rx_data[1]), 
            .I2(n27934), .I3(GND_net), .O(n29496));   // verilog/coms.v(130[12] 305[6])
    defparam i13651_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13648_3_lut (.I0(\data_in_frame[21] [0]), .I1(rx_data[0]), 
            .I2(n27934), .I3(GND_net), .O(n29493));   // verilog/coms.v(130[12] 305[6])
    defparam i13648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13306_3_lut (.I0(t0[3]), .I1(timer[3]), .I2(n3173), .I3(GND_net), 
            .O(n29151));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13642_3_lut (.I0(\data_in_frame[20] [6]), .I1(rx_data[6]), 
            .I2(n27932), .I3(GND_net), .O(n29487));   // verilog/coms.v(130[12] 305[6])
    defparam i13642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13639_3_lut (.I0(\data_in_frame[20] [5]), .I1(rx_data[5]), 
            .I2(n27932), .I3(GND_net), .O(n29484));   // verilog/coms.v(130[12] 305[6])
    defparam i13639_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1677_i23_3_lut (.I0(duty[23]), .I1(duty[22]), .I2(n260), 
            .I3(GND_net), .O(n11586));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13636_3_lut (.I0(\data_in_frame[20] [4]), .I1(rx_data[4]), 
            .I2(n27932), .I3(GND_net), .O(n29481));   // verilog/coms.v(130[12] 305[6])
    defparam i13636_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13307_3_lut (.I0(ID[2]), .I1(data_adj_5899[2]), .I2(n55524), 
            .I3(GND_net), .O(n29152));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13632_3_lut (.I0(\data_in_frame[20] [3]), .I1(rx_data[3]), 
            .I2(n27932), .I3(GND_net), .O(n29477));   // verilog/coms.v(130[12] 305[6])
    defparam i13632_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13308_3_lut (.I0(ID[1]), .I1(data_adj_5899[1]), .I2(n55524), 
            .I3(GND_net), .O(n29153));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13309_3_lut (.I0(t0[2]), .I1(timer[2]), .I2(n3173), .I3(GND_net), 
            .O(n29154));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43163_3_lut (.I0(n4918), .I1(duty[20]), .I2(n9941), .I3(GND_net), 
            .O(n60225));
    defparam i43163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43165_3_lut (.I0(n60225), .I1(n60220), .I2(n9939), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[20]));
    defparam i43165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43160_3_lut (.I0(n4917), .I1(duty[21]), .I2(n9941), .I3(GND_net), 
            .O(n60222));
    defparam i43160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43162_3_lut (.I0(n60222), .I1(n60220), .I2(n9939), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[21]));
    defparam i43162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13623_3_lut (.I0(\data_in_frame[20] [0]), .I1(rx_data[0]), 
            .I2(n27932), .I3(GND_net), .O(n29468));   // verilog/coms.v(130[12] 305[6])
    defparam i13623_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i47114_2_lut (.I0(displacement[0]), .I1(n15_adj_5770), .I2(GND_net), 
            .I3(GND_net), .O(n62934));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam i47114_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i43158_3_lut (.I0(current[15]), .I1(duty[23]), .I2(n9941), 
            .I3(GND_net), .O(n60220));
    defparam i43158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43157_3_lut (.I0(n4916), .I1(duty[22]), .I2(n9941), .I3(GND_net), 
            .O(n60219));
    defparam i43157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43159_3_lut (.I0(n60219), .I1(n60220), .I2(n9939), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[22]));
    defparam i43159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5768_3_lut (.I0(n4915), .I1(current[15]), .I2(n9939), .I3(GND_net), 
            .O(n21266));
    defparam i5768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46251_2_lut (.I0(displacement[1]), .I1(n15_adj_5770), .I2(GND_net), 
            .I3(GND_net), .O(n62948));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam i46251_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5769_3_lut (.I0(n21266), .I1(duty[23]), .I2(n9941), .I3(GND_net), 
            .O(pwm_setpoint_23__N_3[23]));
    defparam i5769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21821_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(n1));
    defparam i21821_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i21822_3_lut (.I0(encoder0_position_scaled[2]), .I1(n1), .I2(n15_adj_5748), 
            .I3(GND_net), .O(n3_adj_5811));
    defparam i21822_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13498_3_lut (.I0(\data_in_frame[15] [0]), .I1(rx_data[0]), 
            .I2(n55152), .I3(GND_net), .O(n29343));   // verilog/coms.v(130[12] 305[6])
    defparam i13498_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13501_3_lut (.I0(\data_in_frame[15] [1]), .I1(rx_data[1]), 
            .I2(n55152), .I3(GND_net), .O(n29346));   // verilog/coms.v(130[12] 305[6])
    defparam i13501_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_245_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[3]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i4_3_lut (.I0(encoder0_position_scaled[3]), .I1(motor_state_23__N_91[3]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[10]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i11_3_lut (.I0(encoder0_position_scaled[10]), .I1(motor_state_23__N_91[10]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13310_3_lut (.I0(t0[1]), .I1(timer[1]), .I2(n3173), .I3(GND_net), 
            .O(n29155));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13504_3_lut (.I0(\data_in_frame[15] [2]), .I1(rx_data[2]), 
            .I2(n55152), .I3(GND_net), .O(n29349));   // verilog/coms.v(130[12] 305[6])
    defparam i13504_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13170_3_lut (.I0(\data_in_frame[6] [4]), .I1(rx_data[4]), .I2(n27904), 
            .I3(GND_net), .O(n29015));   // verilog/coms.v(130[12] 305[6])
    defparam i13170_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13508_3_lut (.I0(\data_in_frame[15] [3]), .I1(rx_data[3]), 
            .I2(n55152), .I3(GND_net), .O(n29353));   // verilog/coms.v(130[12] 305[6])
    defparam i13508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13511_3_lut (.I0(\data_in_frame[15] [4]), .I1(rx_data[4]), 
            .I2(n55152), .I3(GND_net), .O(n29356));   // verilog/coms.v(130[12] 305[6])
    defparam i13511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13514_3_lut (.I0(\data_in_frame[15] [5]), .I1(rx_data[5]), 
            .I2(n55152), .I3(GND_net), .O(n29359));   // verilog/coms.v(130[12] 305[6])
    defparam i13514_3_lut.LUT_INIT = 16'hacac;
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i13311_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5899[7]), 
            .I2(n38386), .I3(n25095), .O(n29156));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13311_4_lut.LUT_INIT = 16'hccac;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(clk16MHz));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFF reset_198 (.Q(reset), .C(clk16MHz), .D(n53805));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk16MHz), .D(displacement_23__N_67[2]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_LUT4 i13067_3_lut (.I0(\data_in_frame[3] [0]), .I1(rx_data[0]), .I2(n27898), 
            .I3(GND_net), .O(n28912));   // verilog/coms.v(130[12] 305[6])
    defparam i13067_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13517_3_lut (.I0(\data_in_frame[15] [6]), .I1(rx_data[6]), 
            .I2(n55152), .I3(GND_net), .O(n29362));   // verilog/coms.v(130[12] 305[6])
    defparam i13517_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[3]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[2]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[1]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[23]), 
           .C(clk16MHz), .D(encoder0_position[21]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_LUT4 i13595_3_lut (.I0(\data_in_frame[18] [7]), .I1(rx_data[7]), 
            .I2(n27929), .I3(GND_net), .O(n29440));   // verilog/coms.v(130[12] 305[6])
    defparam i13595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i589_2_lut (.I0(n1325), .I1(n38194), .I2(GND_net), .I3(GND_net), 
            .O(n2829));   // verilog/TinyFPGA_B.v(392[18] 394[12])
    defparam i589_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_151_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n48255), .O(n1242)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[22]), 
           .C(clk16MHz), .D(encoder0_position[20]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[21]), 
           .C(clk16MHz), .D(encoder0_position[19]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[20]), 
           .C(clk16MHz), .D(encoder0_position[18]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[19]), 
           .C(clk16MHz), .D(encoder0_position[17]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[18]), 
           .C(clk16MHz), .D(encoder0_position[16]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[17]), 
           .C(clk16MHz), .D(encoder0_position[15]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_CARRY add_151_14 (.CI(n48264), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n48265));
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(current[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5706));   // verilog/TinyFPGA_B.v(129[16:24])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[16]), 
           .C(clk16MHz), .D(encoder0_position[14]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_LUT4 i42853_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n59906));
    defparam i42853_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49434_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n6911), .I2(n59906), 
            .I3(n25_adj_5827), .O(n17_adj_5826));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i49434_4_lut.LUT_INIT = 16'h88ba;
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[15]), 
           .C(clk16MHz), .D(encoder0_position[13]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(current[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_5705));   // verilog/TinyFPGA_B.v(129[16:24])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[14]), 
           .C(clk16MHz), .D(encoder0_position[12]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n48407), .I0(GND_net), 
            .I1(n24), .CO(n48408));
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[13]), 
           .C(clk16MHz), .D(encoder0_position[11]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[12]), 
           .C(clk16MHz), .D(encoder0_position[10]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[11]), 
           .C(clk16MHz), .D(encoder0_position[9]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[10]), 
           .C(clk16MHz), .D(encoder0_position[8]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[9]), .C(clk16MHz), 
           .D(encoder0_position[7]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[8]), .C(clk16MHz), 
           .D(encoder0_position[6]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_LUT4 mux_245_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[4]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i5_3_lut (.I0(encoder0_position_scaled[4]), .I1(motor_state_23__N_91[4]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(current[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5704));   // verilog/TinyFPGA_B.v(129[16:24])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[7]), .C(clk16MHz), 
           .D(encoder0_position[5]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_LUT4 i22441_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(100[16:31])
    defparam i22441_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22440_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(98[16:31])
    defparam i22440_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(current[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_5703));   // verilog/TinyFPGA_B.v(129[16:24])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22551_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(96[16:31])
    defparam i22551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13592_3_lut (.I0(\data_in_frame[18] [6]), .I1(rx_data[6]), 
            .I2(n27929), .I3(GND_net), .O(n29437));   // verilog/coms.v(130[12] 305[6])
    defparam i13592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(current[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5702));   // verilog/TinyFPGA_B.v(129[16:24])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_5690), .I3(VCC_net), .O(displacement_23__N_67[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(n25_adj_5690), .CO(n48407));
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(current[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(129[16:24])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[6]), .C(clk16MHz), 
           .D(encoder0_position[4]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[5]), .C(clk16MHz), 
           .D(encoder0_position[3]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[4]), .C(clk16MHz), 
           .D(encoder0_position[2]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[3]), .C(clk16MHz), 
           .D(encoder0_position[1]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_LUT4 mux_245_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[5]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i6_3_lut (.I0(encoder0_position_scaled[5]), .I1(motor_state_23__N_91[5]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(current[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5701));   // verilog/TinyFPGA_B.v(129[16:24])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(current[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5700));   // verilog/TinyFPGA_B.v(129[16:24])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13520_3_lut (.I0(\data_in_frame[15] [7]), .I1(rx_data[7]), 
            .I2(n55152), .I3(GND_net), .O(n29365));   // verilog/coms.v(130[12] 305[6])
    defparam i13520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(current[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5699));   // verilog/TinyFPGA_B.v(129[16:24])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(current[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5698));   // verilog/TinyFPGA_B.v(129[16:24])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(current[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(129[16:24])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_151_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n48263), .O(n1234)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_245_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[6]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i7_3_lut (.I0(encoder0_position_scaled[6]), .I1(motor_state_23__N_91[6]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i3_4_lut (.I0(byte_transmit_counter[5]), .I1(byte_transmit_counter[6]), 
            .I2(n58202), .I3(byte_transmit_counter[7]), .O(n53));   // verilog/coms.v(105[12:33])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk16MHz), .D(displacement_23__N_67[1]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[23]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[22]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[21]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_LUT4 i18720_3_lut (.I0(duty[3]), .I1(duty[0]), .I2(n260), .I3(GND_net), 
            .O(n3));
    defparam i18720_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i2_3_lut (.I0(duty[4]), .I1(duty[1]), .I2(n260), 
            .I3(GND_net), .O(n11628));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i3_3_lut (.I0(duty[5]), .I1(duty[2]), .I2(n260), 
            .I3(GND_net), .O(n11626));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i3_3_lut.LUT_INIT = 16'h3535;
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[20]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_CARRY add_151_13 (.CI(n48263), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n48264));
    SB_LUT4 add_151_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n48283), .O(n1214)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_5 (.CI(n48255), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n48256));
    SB_LUT4 add_151_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n48262), .O(n1235)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[19]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_LUT4 add_151_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n48282), .O(n1215)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1677_i4_3_lut (.I0(duty[6]), .I1(duty[3]), .I2(n260), 
            .I3(GND_net), .O(n11624));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i4_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_151_32 (.CI(n48282), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n48283));
    SB_LUT4 mux_1677_i5_3_lut (.I0(duty[7]), .I1(duty[4]), .I2(n260), 
            .I3(GND_net), .O(n11622));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i5_3_lut.LUT_INIT = 16'h3535;
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[18]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_LUT4 mux_1677_i6_3_lut (.I0(duty[8]), .I1(duty[5]), .I2(n260), 
            .I3(GND_net), .O(n11620));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i7_3_lut (.I0(duty[9]), .I1(duty[6]), .I2(n260), 
            .I3(GND_net), .O(n11618));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 n9941_bdd_4_lut (.I0(n9941), .I1(current[15]), .I2(duty[22]), 
            .I3(n9939), .O(n67005));
    defparam n9941_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n67005_bdd_4_lut (.I0(n67005), .I1(duty[19]), .I2(n4919), 
            .I3(n9939), .O(pwm_setpoint_23__N_3[19]));
    defparam n67005_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9941_bdd_4_lut_49860 (.I0(n9941), .I1(current[15]), .I2(duty[21]), 
            .I3(n9939), .O(n66999));
    defparam n9941_bdd_4_lut_49860.LUT_INIT = 16'he4aa;
    SB_LUT4 n66999_bdd_4_lut (.I0(n66999), .I1(duty[18]), .I2(n4920), 
            .I3(n9939), .O(pwm_setpoint_23__N_3[18]));
    defparam n66999_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9941_bdd_4_lut_49855 (.I0(n9941), .I1(current[15]), .I2(duty[20]), 
            .I3(n9939), .O(n66993));
    defparam n9941_bdd_4_lut_49855.LUT_INIT = 16'he4aa;
    SB_LUT4 n66993_bdd_4_lut (.I0(n66993), .I1(duty[17]), .I2(n4921), 
            .I3(n9939), .O(pwm_setpoint_23__N_3[17]));
    defparam n66993_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9941_bdd_4_lut_49850 (.I0(n9941), .I1(current[15]), .I2(duty[19]), 
            .I3(n9939), .O(n66987));
    defparam n9941_bdd_4_lut_49850.LUT_INIT = 16'he4aa;
    SB_LUT4 n66987_bdd_4_lut (.I0(n66987), .I1(duty[16]), .I2(n4922), 
            .I3(n9939), .O(pwm_setpoint_23__N_3[16]));
    defparam n66987_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9941_bdd_4_lut_49845 (.I0(n9941), .I1(current[15]), .I2(duty[18]), 
            .I3(n9939), .O(n66981));
    defparam n9941_bdd_4_lut_49845.LUT_INIT = 16'he4aa;
    SB_LUT4 n66981_bdd_4_lut (.I0(n66981), .I1(duty[15]), .I2(n4923), 
            .I3(n9939), .O(pwm_setpoint_23__N_3[15]));
    defparam n66981_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9941_bdd_4_lut_49840 (.I0(n9941), .I1(current[15]), .I2(duty[17]), 
            .I3(n9939), .O(n66975));
    defparam n9941_bdd_4_lut_49840.LUT_INIT = 16'he4aa;
    SB_LUT4 n66975_bdd_4_lut (.I0(n66975), .I1(duty[14]), .I2(n4924), 
            .I3(n9939), .O(pwm_setpoint_23__N_3[14]));
    defparam n66975_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9941_bdd_4_lut_49835 (.I0(n9941), .I1(current[15]), .I2(duty[16]), 
            .I3(n9939), .O(n66969));
    defparam n9941_bdd_4_lut_49835.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_1677_i8_3_lut (.I0(duty[10]), .I1(duty[7]), .I2(n260), 
            .I3(GND_net), .O(n11616));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5690));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19933_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[7]));
    defparam i19933_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i8_3_lut (.I0(encoder0_position_scaled[7]), .I1(motor_state_23__N_91[7]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_1677_i9_3_lut (.I0(duty[11]), .I1(duty[8]), .I2(n260), 
            .I3(GND_net), .O(n11614));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut (.I0(state[0]), .I1(n23_adj_5843), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5839));
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13_4_lut (.I0(n35156), .I1(n38711), .I2(state[1]), .I3(n4_adj_5839), 
            .O(n5_adj_5841));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13_4_lut.LUT_INIT = 16'hcafa;
    SB_LUT4 add_151_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n48281), .O(n1216)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_31 (.CI(n48281), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n48282));
    SB_CARRY add_151_12 (.CI(n48262), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n48263));
    SB_LUT4 add_151_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n48280), .O(n1217)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_30 (.CI(n48280), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n48281));
    SB_LUT4 mux_1677_i10_3_lut (.I0(duty[12]), .I1(duty[9]), .I2(n260), 
            .I3(GND_net), .O(n11612));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 add_151_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n48254), .O(n1243)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_4_lut.LUT_INIT = 16'hC33C;
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_151_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n48261), .O(n1236)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_11_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[17]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[16]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[15]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[14]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[13]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[12]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[11]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(clk16MHz), .D(encoder1_position_scaled_23__N_43[10]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[9]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[8]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[7]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[6]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[5]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[4]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[3]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(clk16MHz), 
           .D(encoder1_position_scaled_23__N_43[2]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(clk16MHz), 
           .D(encoder1_position[1]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_LUT4 n66969_bdd_4_lut (.I0(n66969), .I1(duty[13]), .I2(n4925), 
            .I3(n9939), .O(pwm_setpoint_23__N_3[13]));
    defparam n66969_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_151_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n48279), .O(n1218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_29 (.CI(n48279), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n48280));
    SB_LUT4 mux_1677_i11_3_lut (.I0(duty[13]), .I1(duty[10]), .I2(n260), 
            .I3(GND_net), .O(n11610));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 add_151_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n48278), .O(n1219)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9941_bdd_4_lut_49830 (.I0(n9941), .I1(current[15]), .I2(duty[15]), 
            .I3(n9939), .O(n66963));
    defparam n9941_bdd_4_lut_49830.LUT_INIT = 16'he4aa;
    SB_CARRY add_151_11 (.CI(n48261), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n48262));
    SB_LUT4 n66963_bdd_4_lut (.I0(n66963), .I1(duty[12]), .I2(n4926), 
            .I3(n9939), .O(pwm_setpoint_23__N_3[12]));
    defparam n66963_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13206_3_lut (.I0(\data_in_frame[7] [7]), .I1(rx_data[7]), .I2(n27906), 
            .I3(GND_net), .O(n29051));   // verilog/coms.v(130[12] 305[6])
    defparam i13206_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n9941_bdd_4_lut_49825 (.I0(n9941), .I1(current[11]), .I2(duty[14]), 
            .I3(n9939), .O(n66957));
    defparam n9941_bdd_4_lut_49825.LUT_INIT = 16'he4aa;
    SB_LUT4 dti_counter_2038_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[7]), 
            .I3(n49097), .O(n38)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n66957_bdd_4_lut (.I0(n66957), .I1(duty[11]), .I2(n4927), 
            .I3(n9939), .O(pwm_setpoint_23__N_3[11]));
    defparam n66957_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 dti_counter_2038_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[6]), 
            .I3(n49096), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_28 (.CI(n48278), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n48279));
    SB_LUT4 mux_1677_i12_3_lut (.I0(duty[14]), .I1(duty[11]), .I2(n260), 
            .I3(GND_net), .O(n11608));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i12_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_151_4 (.CI(n48254), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n48255));
    SB_CARRY dti_counter_2038_add_4_8 (.CI(n49096), .I0(VCC_net), .I1(dti_counter[6]), 
            .CO(n49097));
    SB_LUT4 dti_counter_2038_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[5]), 
            .I3(n49095), .O(n40_adj_5810)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR dti_counter_2038__i0 (.Q(dti_counter[0]), .C(clk16MHz), .E(n27460), 
            .D(n45), .R(n28642));   // verilog/TinyFPGA_B.v(182[23:37])
    SB_CARRY dti_counter_2038_add_4_7 (.CI(n49095), .I0(VCC_net), .I1(dti_counter[5]), 
            .CO(n49096));
    SB_LUT4 dti_counter_2038_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[4]), 
            .I3(n49094), .O(n41)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2038_add_4_6 (.CI(n49094), .I0(VCC_net), .I1(dti_counter[4]), 
            .CO(n49095));
    SB_LUT4 dti_counter_2038_add_4_5_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[3]), 
            .I3(n49093), .O(n42)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n48277), .O(n1220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2038_add_4_5 (.CI(n49093), .I0(VCC_net), .I1(dti_counter[3]), 
            .CO(n49094));
    SB_LUT4 dti_counter_2038_add_4_4_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[2]), 
            .I3(n49092), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2038_add_4_4 (.CI(n49092), .I0(VCC_net), .I1(dti_counter[2]), 
            .CO(n49093));
    SB_LUT4 dti_counter_2038_add_4_3_lut (.I0(GND_net), .I1(VCC_net), .I2(dti_counter[1]), 
            .I3(n49091), .O(n44)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2038_add_4_3 (.CI(n49091), .I0(VCC_net), .I1(dti_counter[1]), 
            .CO(n49092));
    SB_LUT4 dti_counter_2038_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2038_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2038_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(dti_counter[0]), 
            .CO(n49091));
    SB_CARRY add_151_27 (.CI(n48277), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n48278));
    SB_LUT4 add_151_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n48276), .O(n1221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_1677_i13_3_lut (.I0(duty[15]), .I1(duty[12]), .I2(n260), 
            .I3(GND_net), .O(n11606));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i13_3_lut.LUT_INIT = 16'h3535;
    SB_DFFESR delay_counter__i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n27321), 
            .D(n1244), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_LUT4 mux_1677_i14_3_lut (.I0(duty[16]), .I1(duty[13]), .I2(n260), 
            .I3(GND_net), .O(n11604));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 n9941_bdd_4_lut_49820 (.I0(n9941), .I1(current[10]), .I2(duty[13]), 
            .I3(n9939), .O(n66951));
    defparam n9941_bdd_4_lut_49820.LUT_INIT = 16'he4aa;
    SB_DFFESR delay_counter__i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n27321), 
            .D(n1243), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFFESR delay_counter__i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n27321), 
            .D(n1242), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFFESR delay_counter__i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n27321), 
            .D(n1241), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_LUT4 n66951_bdd_4_lut (.I0(n66951), .I1(duty[10]), .I2(n4928), 
            .I3(n9939), .O(pwm_setpoint_23__N_3[10]));
    defparam n66951_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_4757_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(encoder1_position[19]), 
            .I3(n49510), .O(n15537)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4757_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(encoder1_position[18]), 
            .I3(n49509), .O(n15538)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4757_19 (.CI(n49509), .I0(encoder1_position[17]), .I1(encoder1_position[18]), 
            .CO(n49510));
    SB_LUT4 add_4757_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(encoder1_position[17]), 
            .I3(n49508), .O(n15539)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4757_18 (.CI(n49508), .I0(encoder1_position[16]), .I1(encoder1_position[17]), 
            .CO(n49509));
    SB_LUT4 add_4757_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(encoder1_position[16]), 
            .I3(n49507), .O(n15540)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4757_17 (.CI(n49507), .I0(encoder1_position[15]), .I1(encoder1_position[16]), 
            .CO(n49508));
    SB_LUT4 add_4757_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(encoder1_position[15]), 
            .I3(n49506), .O(n15541)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4757_16 (.CI(n49506), .I0(encoder1_position[14]), .I1(encoder1_position[15]), 
            .CO(n49507));
    SB_LUT4 add_4757_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(encoder1_position[14]), 
            .I3(n49505), .O(n15542)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4757_15 (.CI(n49505), .I0(encoder1_position[13]), .I1(encoder1_position[14]), 
            .CO(n49506));
    SB_LUT4 add_4757_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(encoder1_position[13]), 
            .I3(n49504), .O(n15543)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4757_14 (.CI(n49504), .I0(encoder1_position[12]), .I1(encoder1_position[13]), 
            .CO(n49505));
    SB_LUT4 add_4757_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(encoder1_position[12]), 
            .I3(n49503), .O(n15544)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4757_13 (.CI(n49503), .I0(encoder1_position[11]), .I1(encoder1_position[12]), 
            .CO(n49504));
    SB_LUT4 add_4757_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(encoder1_position[11]), 
            .I3(n49502), .O(n15545)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13203_3_lut (.I0(\data_in_frame[7] [6]), .I1(rx_data[6]), .I2(n27906), 
            .I3(GND_net), .O(n29048));   // verilog/coms.v(130[12] 305[6])
    defparam i13203_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_4757_12 (.CI(n49502), .I0(encoder1_position[10]), .I1(encoder1_position[11]), 
            .CO(n49503));
    SB_LUT4 add_4757_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(encoder1_position[10]), 
            .I3(n49501), .O(n15546)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4757_11 (.CI(n49501), .I0(encoder1_position[9]), .I1(encoder1_position[10]), 
            .CO(n49502));
    SB_LUT4 n9941_bdd_4_lut_49815 (.I0(n9941), .I1(current[9]), .I2(duty[12]), 
            .I3(n9939), .O(n66945));
    defparam n9941_bdd_4_lut_49815.LUT_INIT = 16'he4aa;
    SB_LUT4 add_4757_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(encoder1_position[9]), 
            .I3(n49500), .O(n15547)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4757_10 (.CI(n49500), .I0(encoder1_position[8]), .I1(encoder1_position[9]), 
            .CO(n49501));
    SB_LUT4 add_4757_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(encoder1_position[8]), 
            .I3(n49499), .O(n15548)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13200_3_lut (.I0(\data_in_frame[7] [5]), .I1(rx_data[5]), .I2(n27906), 
            .I3(GND_net), .O(n29045));   // verilog/coms.v(130[12] 305[6])
    defparam i13200_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1677_i15_3_lut (.I0(duty[17]), .I1(duty[14]), .I2(n260), 
            .I3(GND_net), .O(n11602));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i15_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_4757_9 (.CI(n49499), .I0(encoder1_position[7]), .I1(encoder1_position[8]), 
            .CO(n49500));
    SB_LUT4 add_4757_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(encoder1_position[7]), 
            .I3(n49498), .O(n15549)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4757_8 (.CI(n49498), .I0(encoder1_position[6]), .I1(encoder1_position[7]), 
            .CO(n49499));
    SB_LUT4 add_4757_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(encoder1_position[6]), 
            .I3(n49497), .O(n15550)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4757_7 (.CI(n49497), .I0(encoder1_position[5]), .I1(encoder1_position[6]), 
            .CO(n49498));
    SB_LUT4 add_4757_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(encoder1_position[5]), 
            .I3(n49496), .O(n15551)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4757_6 (.CI(n49496), .I0(encoder1_position[4]), .I1(encoder1_position[5]), 
            .CO(n49497));
    SB_LUT4 add_4757_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(encoder1_position[4]), 
            .I3(n49495), .O(n15552)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4757_5 (.CI(n49495), .I0(encoder1_position[3]), .I1(encoder1_position[4]), 
            .CO(n49496));
    SB_DFFESR delay_counter__i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n27321), 
            .D(n1240), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_LUT4 add_4757_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(encoder1_position[3]), 
            .I3(n49494), .O(n15553)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4757_4 (.CI(n49494), .I0(encoder1_position[2]), .I1(encoder1_position[3]), 
            .CO(n49495));
    SB_LUT4 add_4757_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(encoder1_position[2]), 
            .I3(n49493), .O(n15554)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13197_3_lut (.I0(\data_in_frame[7] [4]), .I1(rx_data[4]), .I2(n27906), 
            .I3(GND_net), .O(n29042));   // verilog/coms.v(130[12] 305[6])
    defparam i13197_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_4757_3 (.CI(n49493), .I0(encoder1_position[1]), .I1(encoder1_position[2]), 
            .CO(n49494));
    SB_LUT4 add_4757_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(encoder1_position[1]), 
            .I3(GND_net), .O(n15555)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4757_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4757_2 (.CI(GND_net), .I0(encoder1_position[0]), .I1(encoder1_position[1]), 
            .CO(n49493));
    SB_LUT4 n66945_bdd_4_lut (.I0(n66945), .I1(duty[9]), .I2(n4929), .I3(n9939), 
            .O(pwm_setpoint_23__N_3[9]));
    defparam n66945_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1677_i16_3_lut (.I0(duty[18]), .I1(duty[15]), .I2(n260), 
            .I3(GND_net), .O(n11600));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 n9941_bdd_4_lut_49810 (.I0(n9941), .I1(current[8]), .I2(duty[11]), 
            .I3(n9939), .O(n66939));
    defparam n9941_bdd_4_lut_49810.LUT_INIT = 16'he4aa;
    SB_LUT4 n66939_bdd_4_lut (.I0(n66939), .I1(duty[8]), .I2(n4930), .I3(n9939), 
            .O(pwm_setpoint_23__N_3[8]));
    defparam n66939_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut (.I0(ID[4]), .I1(ID[7]), .I2(ID[6]), .I3(ID[5]), 
            .O(n14_adj_5844));   // verilog/TinyFPGA_B.v(386[12:17])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(ID[0]), .I1(ID[1]), .I2(ID[3]), .I3(ID[2]), 
            .O(n13_adj_5845));   // verilog/TinyFPGA_B.v(386[12:17])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22454_4_lut (.I0(n13_adj_5845), .I1(baudrate[0]), .I2(n14_adj_5844), 
            .I3(n25108), .O(n38194));
    defparam i22454_4_lut.LUT_INIT = 16'hc8fa;
    SB_LUT4 n9941_bdd_4_lut_49805 (.I0(n9941), .I1(current[7]), .I2(duty[10]), 
            .I3(n9939), .O(n66933));
    defparam n9941_bdd_4_lut_49805.LUT_INIT = 16'he4aa;
    SB_LUT4 n66933_bdd_4_lut (.I0(n66933), .I1(duty[7]), .I2(n4931), .I3(n9939), 
            .O(pwm_setpoint_23__N_3[7]));
    defparam n66933_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/luis/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFFE \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n17_adj_5826));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(clk16MHz), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(151[9] 230[5])
    SB_LUT4 add_151_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n48260), .O(n1237)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13188_3_lut (.I0(\data_in_frame[7] [2]), .I1(rx_data[2]), .I2(n27906), 
            .I3(GND_net), .O(n29033));   // verilog/coms.v(130[12] 305[6])
    defparam i13188_3_lut.LUT_INIT = 16'hacac;
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(clk16MHz), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(151[9] 230[5])
    SB_LUT4 add_1190_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_207), 
            .I3(n48375), .O(n4915)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_26 (.CI(n48276), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n48277));
    SB_LUT4 i13185_3_lut (.I0(\data_in_frame[7] [1]), .I1(rx_data[1]), .I2(n27906), 
            .I3(GND_net), .O(n29030));   // verilog/coms.v(130[12] 305[6])
    defparam i13185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_151_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n48253), .O(n1244)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[23]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_LUT4 n9941_bdd_4_lut_49800 (.I0(n9941), .I1(current[6]), .I2(duty[9]), 
            .I3(n9939), .O(n66927));
    defparam n9941_bdd_4_lut_49800.LUT_INIT = 16'he4aa;
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[22]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[21]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[20]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[19]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[18]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[17]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_LUT4 add_1190_24_lut (.I0(GND_net), .I1(GND_net), .I2(n11586), 
            .I3(n48374), .O(n4916)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_24 (.CI(n48374), .I0(GND_net), .I1(n11586), .CO(n48375));
    SB_CARRY add_151_10 (.CI(n48260), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n48261));
    SB_LUT4 add_151_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n48275), .O(n1222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n48259), .O(n1238)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_25 (.CI(n48275), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n48276));
    SB_LUT4 add_151_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n48274), .O(n1223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_3 (.CI(n48253), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n48254));
    SB_DFFESR dti_counter_2038__i7 (.Q(dti_counter[7]), .C(clk16MHz), .E(n27460), 
            .D(n38), .R(n28642));   // verilog/TinyFPGA_B.v(182[23:37])
    SB_DFFESR dti_counter_2038__i6 (.Q(dti_counter[6]), .C(clk16MHz), .E(n27460), 
            .D(n39), .R(n28642));   // verilog/TinyFPGA_B.v(182[23:37])
    SB_DFFESR dti_counter_2038__i5 (.Q(dti_counter[5]), .C(clk16MHz), .E(n27460), 
            .D(n40_adj_5810), .R(n28642));   // verilog/TinyFPGA_B.v(182[23:37])
    SB_DFFESR dti_counter_2038__i4 (.Q(dti_counter[4]), .C(clk16MHz), .E(n27460), 
            .D(n41), .R(n28642));   // verilog/TinyFPGA_B.v(182[23:37])
    SB_DFFESR dti_counter_2038__i3 (.Q(dti_counter[3]), .C(clk16MHz), .E(n27460), 
            .D(n42), .R(n28642));   // verilog/TinyFPGA_B.v(182[23:37])
    SB_DFFESR dti_counter_2038__i2 (.Q(dti_counter[2]), .C(clk16MHz), .E(n27460), 
            .D(n43), .R(n28642));   // verilog/TinyFPGA_B.v(182[23:37])
    SB_DFFESR dti_counter_2038__i1 (.Q(dti_counter[1]), .C(clk16MHz), .E(n27460), 
            .D(n44), .R(n28642));   // verilog/TinyFPGA_B.v(182[23:37])
    SB_LUT4 add_1190_23_lut (.I0(GND_net), .I1(GND_net), .I2(n11588), 
            .I3(n48373), .O(n4917)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_23_lut.LUT_INIT = 16'hC33C;
    SB_DFF read_197 (.Q(state_7__N_3918[0]), .C(clk16MHz), .D(n58312));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(clk16MHz), 
           .D(n56301));   // verilog/TinyFPGA_B.v(151[9] 230[5])
    SB_LUT4 add_4650_23_lut (.I0(GND_net), .I1(n13241), .I2(encoder1_position[23]), 
            .I3(n48583), .O(encoder1_position_scaled_23__N_43[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut (.I0(hall2), .I1(commutation_state_7__N_27[2]), .I2(GND_net), 
            .I3(GND_net), .O(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(174[7:32])
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_DFFESR delay_counter__i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n27321), 
            .D(n1239), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_LUT4 add_4650_22_lut (.I0(GND_net), .I1(n13242), .I2(encoder1_position[22]), 
            .I3(n48582), .O(encoder1_position_scaled_23__N_43[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4650_22 (.CI(n48582), .I0(n13242), .I1(encoder1_position[22]), 
            .CO(n48583));
    SB_LUT4 add_4650_21_lut (.I0(GND_net), .I1(n13243), .I2(encoder1_position[21]), 
            .I3(n48581), .O(encoder1_position_scaled_23__N_43[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4650_21 (.CI(n48581), .I0(n13243), .I1(encoder1_position[21]), 
            .CO(n48582));
    SB_LUT4 add_4650_20_lut (.I0(GND_net), .I1(n13244), .I2(encoder1_position[20]), 
            .I3(n48580), .O(encoder1_position_scaled_23__N_43[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4650_20 (.CI(n48580), .I0(n13244), .I1(encoder1_position[20]), 
            .CO(n48581));
    SB_CARRY add_1190_23 (.CI(n48373), .I0(GND_net), .I1(n11588), .CO(n48374));
    SB_LUT4 add_1190_22_lut (.I0(GND_net), .I1(GND_net), .I2(n11590), 
            .I3(n48372), .O(n4918)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n66927_bdd_4_lut (.I0(n66927), .I1(duty[6]), .I2(n4932), .I3(n9939), 
            .O(pwm_setpoint_23__N_3[6]));
    defparam n66927_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_4650_19_lut (.I0(GND_net), .I1(n13245), .I2(encoder1_position[19]), 
            .I3(n48579), .O(encoder1_position_scaled_23__N_43[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_19_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[16]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_CARRY add_151_9 (.CI(n48259), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n48260));
    SB_CARRY add_151_24 (.CI(n48274), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n48275));
    SB_CARRY add_4650_19 (.CI(n48579), .I0(n13245), .I1(encoder1_position[19]), 
            .CO(n48580));
    SB_LUT4 add_4650_18_lut (.I0(GND_net), .I1(n13246), .I2(encoder1_position[18]), 
            .I3(n48578), .O(encoder1_position_scaled_23__N_43[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_18_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[15]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[14]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[13]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[12]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[11]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[10]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[9]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[8]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[7]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[6]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[5]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[4]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_LUT4 i1_3_lut (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(commutation_state_7__N_208[0]));   // verilog/TinyFPGA_B.v(171[4] 173[7])
    defparam i1_3_lut.LUT_INIT = 16'h1414;
    SB_DFFESR delay_counter__i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n27321), 
            .D(n1238), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFFESR delay_counter__i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n27321), 
            .D(n1237), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFFESR delay_counter__i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n27321), 
            .D(n1236), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_CARRY add_4650_18 (.CI(n48578), .I0(n13246), .I1(encoder1_position[18]), 
            .CO(n48579));
    SB_LUT4 add_4650_17_lut (.I0(GND_net), .I1(n13247), .I2(encoder1_position[17]), 
            .I3(n48577), .O(encoder1_position_scaled_23__N_43[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4650_17 (.CI(n48577), .I0(n13247), .I1(encoder1_position[17]), 
            .CO(n48578));
    SB_CARRY add_1190_22 (.CI(n48372), .I0(GND_net), .I1(n11590), .CO(n48373));
    SB_LUT4 add_1190_21_lut (.I0(GND_net), .I1(GND_net), .I2(n11592), 
            .I3(n48371), .O(n4919)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9941_bdd_4_lut_49795 (.I0(n9941), .I1(current[5]), .I2(duty[8]), 
            .I3(n9939), .O(n66921));
    defparam n9941_bdd_4_lut_49795.LUT_INIT = 16'he4aa;
    SB_LUT4 add_4650_16_lut (.I0(GND_net), .I1(n13248), .I2(encoder1_position[16]), 
            .I3(n48576), .O(encoder1_position_scaled_23__N_43[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4650_16 (.CI(n48576), .I0(n13248), .I1(encoder1_position[16]), 
            .CO(n48577));
    SB_LUT4 add_4650_15_lut (.I0(GND_net), .I1(n13249), .I2(encoder1_position[15]), 
            .I3(n48575), .O(encoder1_position_scaled_23__N_43[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4650_15 (.CI(n48575), .I0(n13249), .I1(encoder1_position[15]), 
            .CO(n48576));
    SB_LUT4 add_4650_14_lut (.I0(GND_net), .I1(n13250), .I2(encoder1_position[14]), 
            .I3(n48574), .O(encoder1_position_scaled_23__N_43[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_14_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i10 (.Q(delay_counter[10]), .C(clk16MHz), .E(n27321), 
            .D(n1235), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_CARRY add_4650_14 (.CI(n48574), .I0(n13250), .I1(encoder1_position[14]), 
            .CO(n48575));
    SB_LUT4 add_4650_13_lut (.I0(GND_net), .I1(n13251), .I2(encoder1_position[13]), 
            .I3(n48573), .O(encoder1_position_scaled_23__N_43[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4650_13 (.CI(n48573), .I0(n13251), .I1(encoder1_position[13]), 
            .CO(n48574));
    SB_LUT4 add_4650_12_lut (.I0(GND_net), .I1(n13252), .I2(encoder1_position[12]), 
            .I3(n48572), .O(encoder1_position_scaled_23__N_43[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_21 (.CI(n48371), .I0(GND_net), .I1(n11592), .CO(n48372));
    SB_LUT4 add_1190_20_lut (.I0(GND_net), .I1(GND_net), .I2(n11594), 
            .I3(n48370), .O(n4920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4650_12 (.CI(n48572), .I0(n13252), .I1(encoder1_position[12]), 
            .CO(n48573));
    SB_LUT4 add_151_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n48273), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4650_11_lut (.I0(GND_net), .I1(n13253), .I2(encoder1_position[11]), 
            .I3(n48571), .O(encoder1_position_scaled_23__N_43[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4650_11 (.CI(n48571), .I0(n13253), .I1(encoder1_position[11]), 
            .CO(n48572));
    SB_LUT4 add_4650_10_lut (.I0(GND_net), .I1(n13254), .I2(encoder1_position[10]), 
            .I3(n48570), .O(encoder1_position_scaled_23__N_43[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4650_10 (.CI(n48570), .I0(n13254), .I1(encoder1_position[10]), 
            .CO(n48571));
    SB_LUT4 add_4650_9_lut (.I0(GND_net), .I1(n13255), .I2(encoder1_position[9]), 
            .I3(n48569), .O(encoder1_position_scaled_23__N_43[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4650_9 (.CI(n48569), .I0(n13255), .I1(encoder1_position[9]), 
            .CO(n48570));
    SB_LUT4 i2_3_lut (.I0(\data_in_frame[16] [2]), .I1(n50260), .I2(n25895), 
            .I3(GND_net), .O(n56120));
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1729 (.I0(n55775), .I1(\data_in_frame[20] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5814));
    defparam i2_2_lut_adj_1729.LUT_INIT = 16'h6666;
    SB_LUT4 add_4650_8_lut (.I0(GND_net), .I1(n13256), .I2(encoder1_position[8]), 
            .I3(n48568), .O(encoder1_position_scaled_23__N_43[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_20 (.CI(n48370), .I0(GND_net), .I1(n11594), .CO(n48371));
    SB_CARRY add_4650_8 (.CI(n48568), .I0(n13256), .I1(encoder1_position[8]), 
            .CO(n48569));
    SB_LUT4 add_1190_19_lut (.I0(GND_net), .I1(GND_net), .I2(n11596), 
            .I3(n48369), .O(n4921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_23 (.CI(n48273), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n48274));
    SB_LUT4 i6_4_lut_adj_1730 (.I0(n56120), .I1(\data_in_frame[18] [4]), 
            .I2(\data_in_frame[18] [5]), .I3(\data_in_frame[19] [0]), .O(n14_adj_5813));
    defparam i6_4_lut_adj_1730.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(\data_in_frame[21] [0]), .I1(n14_adj_5813), .I2(n10_adj_5814), 
            .I3(n24804), .O(n57376));
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4650_7_lut (.I0(GND_net), .I1(n13257), .I2(encoder1_position[7]), 
            .I3(n48567), .O(encoder1_position_scaled_23__N_43[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4650_7 (.CI(n48567), .I0(n13257), .I1(encoder1_position[7]), 
            .CO(n48568));
    SB_LUT4 add_4650_6_lut (.I0(GND_net), .I1(n13258), .I2(encoder1_position[6]), 
            .I3(n48566), .O(encoder1_position_scaled_23__N_43[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_19 (.CI(n48369), .I0(GND_net), .I1(n11596), .CO(n48370));
    SB_CARRY add_4650_6 (.CI(n48566), .I0(n13258), .I1(encoder1_position[6]), 
            .CO(n48567));
    SB_LUT4 add_1190_18_lut (.I0(GND_net), .I1(GND_net), .I2(n11598), 
            .I3(n48368), .O(n4922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n48272), .O(n1225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4650_5_lut (.I0(GND_net), .I1(n13259), .I2(encoder1_position[5]), 
            .I3(n48565), .O(encoder1_position_scaled_23__N_43[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4650_5 (.CI(n48565), .I0(n13259), .I1(encoder1_position[5]), 
            .CO(n48566));
    SB_LUT4 add_4650_4_lut (.I0(GND_net), .I1(n13260), .I2(encoder1_position[4]), 
            .I3(n48564), .O(encoder1_position_scaled_23__N_43[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4650_4 (.CI(n48564), .I0(n13260), .I1(encoder1_position[4]), 
            .CO(n48565));
    SB_LUT4 add_4650_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(encoder1_position[3]), 
            .I3(n48563), .O(encoder1_position_scaled_23__N_43[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_18 (.CI(n48368), .I0(GND_net), .I1(n11598), .CO(n48369));
    SB_CARRY add_4650_3 (.CI(n48563), .I0(encoder1_position[1]), .I1(encoder1_position[3]), 
            .CO(n48564));
    SB_LUT4 add_4650_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(encoder1_position[2]), 
            .I3(GND_net), .O(encoder1_position_scaled_23__N_43[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4650_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4650_2 (.CI(GND_net), .I0(encoder1_position[0]), .I1(encoder1_position[2]), 
            .CO(n48563));
    SB_LUT4 add_4762_21_lut (.I0(GND_net), .I1(n15537), .I2(encoder1_position[21]), 
            .I3(n48562), .O(n13241)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4762_20_lut (.I0(GND_net), .I1(n15538), .I2(encoder1_position[20]), 
            .I3(n48561), .O(n13242)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4762_20 (.CI(n48561), .I0(n15538), .I1(encoder1_position[20]), 
            .CO(n48562));
    SB_LUT4 add_4762_19_lut (.I0(GND_net), .I1(n15539), .I2(encoder1_position[19]), 
            .I3(n48560), .O(n13243)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4762_19 (.CI(n48560), .I0(n15539), .I1(encoder1_position[19]), 
            .CO(n48561));
    SB_LUT4 add_4762_18_lut (.I0(GND_net), .I1(n15540), .I2(encoder1_position[18]), 
            .I3(n48559), .O(n13244)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4762_18 (.CI(n48559), .I0(n15540), .I1(encoder1_position[18]), 
            .CO(n48560));
    SB_LUT4 n66921_bdd_4_lut (.I0(n66921), .I1(duty[5]), .I2(n4933), .I3(n9939), 
            .O(pwm_setpoint_23__N_3[5]));
    defparam n66921_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_4762_17_lut (.I0(GND_net), .I1(n15541), .I2(encoder1_position[17]), 
            .I3(n48558), .O(n13245)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4762_17 (.CI(n48558), .I0(n15541), .I1(encoder1_position[17]), 
            .CO(n48559));
    SB_LUT4 add_4762_16_lut (.I0(GND_net), .I1(n15542), .I2(encoder1_position[16]), 
            .I3(n48557), .O(n13246)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4762_16 (.CI(n48557), .I0(n15542), .I1(encoder1_position[16]), 
            .CO(n48558));
    SB_LUT4 add_4762_15_lut (.I0(GND_net), .I1(n15543), .I2(encoder1_position[15]), 
            .I3(n48556), .O(n13247)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4762_15 (.CI(n48556), .I0(n15543), .I1(encoder1_position[15]), 
            .CO(n48557));
    SB_LUT4 add_4762_14_lut (.I0(GND_net), .I1(n15544), .I2(encoder1_position[14]), 
            .I3(n48555), .O(n13248)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4762_14 (.CI(n48555), .I0(n15544), .I1(encoder1_position[14]), 
            .CO(n48556));
    SB_LUT4 add_4762_13_lut (.I0(GND_net), .I1(n15545), .I2(encoder1_position[13]), 
            .I3(n48554), .O(n13249)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4762_13 (.CI(n48554), .I0(n15545), .I1(encoder1_position[13]), 
            .CO(n48555));
    SB_LUT4 add_4762_12_lut (.I0(GND_net), .I1(n15546), .I2(encoder1_position[12]), 
            .I3(n48553), .O(n13250)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4762_12 (.CI(n48553), .I0(n15546), .I1(encoder1_position[12]), 
            .CO(n48554));
    SB_LUT4 add_4762_11_lut (.I0(GND_net), .I1(n15547), .I2(encoder1_position[11]), 
            .I3(n48552), .O(n13251)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4762_11 (.CI(n48552), .I0(n15547), .I1(encoder1_position[11]), 
            .CO(n48553));
    SB_LUT4 add_4762_10_lut (.I0(GND_net), .I1(n15548), .I2(encoder1_position[10]), 
            .I3(n48551), .O(n13252)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4762_10 (.CI(n48551), .I0(n15548), .I1(encoder1_position[10]), 
            .CO(n48552));
    SB_LUT4 add_4762_9_lut (.I0(GND_net), .I1(n15549), .I2(encoder1_position[9]), 
            .I3(n48550), .O(n13253)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n27321), 
            .D(n1245), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_CARRY add_4762_9 (.CI(n48550), .I0(n15549), .I1(encoder1_position[9]), 
            .CO(n48551));
    SB_LUT4 add_4762_8_lut (.I0(GND_net), .I1(n15550), .I2(encoder1_position[8]), 
            .I3(n48549), .O(n13254)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4762_8 (.CI(n48549), .I0(n15550), .I1(encoder1_position[8]), 
            .CO(n48550));
    SB_DFFESR GHC_192 (.Q(GHC), .C(clk16MHz), .E(n27236), .D(GHC_N_391), 
            .R(n28348));   // verilog/TinyFPGA_B.v(151[9] 230[5])
    SB_LUT4 add_4762_7_lut (.I0(GND_net), .I1(n15551), .I2(encoder1_position[7]), 
            .I3(n48548), .O(n13255)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR GHB_190 (.Q(GHB), .C(clk16MHz), .E(n27236), .D(GHB_N_377), 
            .R(n28348));   // verilog/TinyFPGA_B.v(151[9] 230[5])
    SB_CARRY add_4762_7 (.CI(n48548), .I0(n15551), .I1(encoder1_position[7]), 
            .CO(n48549));
    SB_DFFESR GHA_188 (.Q(GHA), .C(clk16MHz), .E(n27236), .D(GHA_N_355), 
            .R(n28348));   // verilog/TinyFPGA_B.v(151[9] 230[5])
    SB_LUT4 add_4762_6_lut (.I0(GND_net), .I1(n15552), .I2(encoder1_position[6]), 
            .I3(n48547), .O(n13256)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(clk16MHz), 
            .E(n7_adj_5846), .D(commutation_state_7__N_208[0]), .S(commutation_state_7__N_216));   // verilog/TinyFPGA_B.v(151[9] 230[5])
    SB_CARRY add_4762_6 (.CI(n48547), .I0(n15552), .I1(encoder1_position[6]), 
            .CO(n48548));
    SB_DFFESR GLA_189 (.Q(INLA_c_0), .C(clk16MHz), .E(n27236), .D(GLA_N_372), 
            .R(n28348));   // verilog/TinyFPGA_B.v(151[9] 230[5])
    SB_DFFESR GLB_191 (.Q(INLB_c_0), .C(clk16MHz), .E(n27236), .D(GLB_N_386), 
            .R(n28348));   // verilog/TinyFPGA_B.v(151[9] 230[5])
    SB_LUT4 add_4762_5_lut (.I0(GND_net), .I1(n15553), .I2(encoder1_position[5]), 
            .I3(n48546), .O(n13257)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4762_5 (.CI(n48546), .I0(n15553), .I1(encoder1_position[5]), 
            .CO(n48547));
    SB_DFFESR GLC_193 (.Q(INLC_c_0), .C(clk16MHz), .E(n27236), .D(GLC_N_400), 
            .R(n28348));   // verilog/TinyFPGA_B.v(151[9] 230[5])
    SB_LUT4 add_1190_17_lut (.I0(GND_net), .I1(GND_net), .I2(n11600), 
            .I3(n48367), .O(n4923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_17_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i11 (.Q(delay_counter[11]), .C(clk16MHz), .E(n27321), 
            .D(n1234), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_LUT4 add_4762_4_lut (.I0(GND_net), .I1(n15554), .I2(encoder1_position[4]), 
            .I3(n48545), .O(n13258)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4762_4 (.CI(n48545), .I0(n15554), .I1(encoder1_position[4]), 
            .CO(n48546));
    SB_CARRY add_1190_17 (.CI(n48367), .I0(GND_net), .I1(n11600), .CO(n48368));
    SB_LUT4 add_4762_3_lut (.I0(GND_net), .I1(n15555), .I2(encoder1_position[3]), 
            .I3(n48544), .O(n13259)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4762_3 (.CI(n48544), .I0(n15555), .I1(encoder1_position[3]), 
            .CO(n48545));
    SB_LUT4 add_1190_16_lut (.I0(GND_net), .I1(GND_net), .I2(n11602), 
            .I3(n48366), .O(n4924)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4762_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(encoder1_position[2]), 
            .I3(GND_net), .O(n13260)) /* synthesis syn_instantiated=1 */ ;
    defparam add_4762_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4762_2 (.CI(GND_net), .I0(encoder1_position[0]), .I1(encoder1_position[2]), 
            .CO(n48544));
    GND i1 (.Y(GND_net));
    SB_CARRY add_151_22 (.CI(n48272), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n48273));
    SB_LUT4 add_151_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n48258), .O(n1239)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_16 (.CI(n48366), .I0(GND_net), .I1(n11602), .CO(n48367));
    SB_LUT4 LessThan_1181_i15_2_lut (.I0(r_Clock_Count_adj_5923[7]), .I1(o_Rx_DV_N_3488[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5804));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1181_i9_2_lut (.I0(r_Clock_Count_adj_5923[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5800));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_1190_15_lut (.I0(GND_net), .I1(GND_net), .I2(n11604), 
            .I3(n48365), .O(n4925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_15 (.CI(n48365), .I0(GND_net), .I1(n11604), .CO(n48366));
    SB_LUT4 LessThan_1181_i13_2_lut (.I0(r_Clock_Count_adj_5923[6]), .I1(o_Rx_DV_N_3488[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5802));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_1181_i11_2_lut (.I0(r_Clock_Count_adj_5923[5]), .I1(o_Rx_DV_N_3488[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5801));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_1190_14_lut (.I0(GND_net), .I1(GND_net), .I2(n11606), 
            .I3(n48364), .O(n4926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_14_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i12 (.Q(delay_counter[12]), .C(clk16MHz), .E(n27321), 
            .D(n1233), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_CARRY add_1190_14 (.CI(n48364), .I0(GND_net), .I1(n11606), .CO(n48365));
    SB_LUT4 add_1190_13_lut (.I0(GND_net), .I1(GND_net), .I2(n11608), 
            .I3(n48363), .O(n4927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_13 (.CI(n48363), .I0(GND_net), .I1(n11608), .CO(n48364));
    SB_LUT4 LessThan_1181_i4_4_lut (.I0(r_Clock_Count_adj_5923[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count_adj_5923[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5797));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i1_2_lut_adj_1731 (.I0(\data_in_frame[16] [6]), .I1(n25941), 
            .I2(GND_net), .I3(GND_net), .O(n56183));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1731.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1732 (.I0(\data_in_frame[19] [2]), .I1(n56183), 
            .I2(n55985), .I3(n55655), .O(n32987));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1732.LUT_INIT = 16'h6996;
    SB_LUT4 add_1190_12_lut (.I0(GND_net), .I1(GND_net), .I2(n11610), 
            .I3(n48362), .O(n4928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_12 (.CI(n48362), .I0(GND_net), .I1(n11610), .CO(n48363));
    SB_LUT4 add_1190_11_lut (.I0(GND_net), .I1(GND_net), .I2(n11612), 
            .I3(n48361), .O(n4929)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_11 (.CI(n48361), .I0(GND_net), .I1(n11612), .CO(n48362));
    SB_LUT4 i48753_3_lut (.I0(n4_adj_5797), .I1(o_Rx_DV_N_3488[5]), .I2(n11_adj_5801), 
            .I3(GND_net), .O(n65815));   // verilog/uart_tx.v(117[17:57])
    defparam i48753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48754_3_lut (.I0(n65815), .I1(o_Rx_DV_N_3488[6]), .I2(n13_adj_5802), 
            .I3(GND_net), .O(n65816));   // verilog/uart_tx.v(117[17:57])
    defparam i48754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1733 (.I0(\data_in_frame[16] [7]), .I1(n57943), 
            .I2(\data_in_frame[14] [6]), .I3(\data_in_frame[17] [0]), .O(n55655));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1733.LUT_INIT = 16'h9669;
    SB_LUT4 add_1190_10_lut (.I0(GND_net), .I1(GND_net), .I2(n11614), 
            .I3(n48360), .O(n4930)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_10 (.CI(n48360), .I0(GND_net), .I1(n11614), .CO(n48361));
    SB_LUT4 add_1190_9_lut (.I0(GND_net), .I1(GND_net), .I2(n11616), .I3(n48359), 
            .O(n4931)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_1734 (.I0(\data_in_frame[19] [1]), .I1(n55655), 
            .I2(n50264), .I3(GND_net), .O(n56050));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1734.LUT_INIT = 16'h9696;
    SB_LUT4 i47353_4_lut (.I0(n13_adj_5802), .I1(n11_adj_5801), .I2(n9_adj_5800), 
            .I3(n63461), .O(n64415));
    defparam i47353_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_1181_i8_3_lut (.I0(n6_adj_5798), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5800), .I3(GND_net), .O(n8_adj_5799));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1735 (.I0(\data_in_frame[18] [7]), .I1(n56050), 
            .I2(n55648), .I3(n55624), .O(n25705));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1735.LUT_INIT = 16'h6996;
    SB_LUT4 i48443_3_lut (.I0(n65816), .I1(o_Rx_DV_N_3488[7]), .I2(n15_adj_5804), 
            .I3(GND_net), .O(n14_adj_5803));   // verilog/uart_tx.v(117[17:57])
    defparam i48443_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1190_9 (.CI(n48359), .I0(GND_net), .I1(n11616), .CO(n48360));
    SB_LUT4 add_1190_8_lut (.I0(GND_net), .I1(GND_net), .I2(n11618), .I3(n48358), 
            .O(n4932)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_8 (.CI(n48358), .I0(GND_net), .I1(n11618), .CO(n48359));
    SB_LUT4 n9941_bdd_4_lut_49790 (.I0(n9941), .I1(current[4]), .I2(duty[7]), 
            .I3(n9939), .O(n66915));
    defparam n9941_bdd_4_lut_49790.LUT_INIT = 16'he4aa;
    SB_LUT4 i48061_4_lut (.I0(n14_adj_5803), .I1(n8_adj_5799), .I2(n15_adj_5804), 
            .I3(n64415), .O(n65123));   // verilog/uart_tx.v(117[17:57])
    defparam i48061_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48062_3_lut (.I0(n65123), .I1(o_Rx_DV_N_3488[8]), .I2(r_Clock_Count_adj_5923[8]), 
            .I3(GND_net), .O(n5228));   // verilog/uart_tx.v(117[17:57])
    defparam i48062_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_1190_7_lut (.I0(GND_net), .I1(GND_net), .I2(n11620), .I3(n48357), 
            .O(n4933)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_7 (.CI(n48357), .I0(GND_net), .I1(n11620), .CO(n48358));
    SB_LUT4 add_1190_6_lut (.I0(GND_net), .I1(GND_net), .I2(n11622), .I3(n48356), 
            .O(n4934)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n66915_bdd_4_lut (.I0(n66915), .I1(duty[4]), .I2(n4934), .I3(n9939), 
            .O(pwm_setpoint_23__N_3[4]));
    defparam n66915_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_1190_6 (.CI(n48356), .I0(GND_net), .I1(n11622), .CO(n48357));
    SB_LUT4 add_1190_5_lut (.I0(GND_net), .I1(GND_net), .I2(n11624), .I3(n48355), 
            .O(n4935)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_5 (.CI(n48355), .I0(GND_net), .I1(n11624), .CO(n48356));
    SB_LUT4 add_1190_4_lut (.I0(GND_net), .I1(GND_net), .I2(n11626), .I3(n48354), 
            .O(n4936)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_4 (.CI(n48354), .I0(GND_net), .I1(n11626), .CO(n48355));
    SB_LUT4 add_1190_3_lut (.I0(GND_net), .I1(GND_net), .I2(n11628), .I3(n48353), 
            .O(n4937)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12497_2_lut (.I0(n27236), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n28348));   // verilog/TinyFPGA_B.v(151[9] 230[5])
    defparam i12497_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_1190_3 (.CI(n48353), .I0(GND_net), .I1(n11628), .CO(n48354));
    SB_LUT4 add_1190_2_lut (.I0(GND_net), .I1(GND_net), .I2(n3), .I3(VCC_net), 
            .O(n4938)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1190_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n48271), .O(n1226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1190_2 (.CI(VCC_net), .I0(GND_net), .I1(n3), .CO(n48353));
    SB_CARRY add_151_21 (.CI(n48271), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n48272));
    SB_LUT4 n9941_bdd_4_lut_49785 (.I0(n9941), .I1(current[3]), .I2(duty[6]), 
            .I3(n9939), .O(n66909));
    defparam n9941_bdd_4_lut_49785.LUT_INIT = 16'he4aa;
    SB_LUT4 n66909_bdd_4_lut (.I0(n66909), .I1(duty[3]), .I2(n4935), .I3(n9939), 
            .O(pwm_setpoint_23__N_3[3]));
    defparam n66909_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9941_bdd_4_lut_49780 (.I0(n9941), .I1(current[2]), .I2(duty[5]), 
            .I3(n9939), .O(n66903));
    defparam n9941_bdd_4_lut_49780.LUT_INIT = 16'he4aa;
    SB_LUT4 n66903_bdd_4_lut (.I0(n66903), .I1(duty[2]), .I2(n4936), .I3(n9939), 
            .O(pwm_setpoint_23__N_3[2]));
    defparam n66903_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9941_bdd_4_lut_49775 (.I0(n9941), .I1(current[1]), .I2(duty[4]), 
            .I3(n9939), .O(n66897));
    defparam n9941_bdd_4_lut_49775.LUT_INIT = 16'he4aa;
    SB_LUT4 n66897_bdd_4_lut (.I0(n66897), .I1(duty[1]), .I2(n4937), .I3(n9939), 
            .O(pwm_setpoint_23__N_3[1]));
    defparam n66897_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9941_bdd_4_lut_49770 (.I0(n9941), .I1(current[0]), .I2(duty[3]), 
            .I3(n9939), .O(n66891));
    defparam n9941_bdd_4_lut_49770.LUT_INIT = 16'he4aa;
    SB_LUT4 n66891_bdd_4_lut (.I0(n66891), .I1(duty[0]), .I2(n4938), .I3(n9939), 
            .O(pwm_setpoint_23__N_3[0]));
    defparam n66891_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i49193_4_lut (.I0(commutation_state[1]), .I1(n22471), .I2(dti), 
            .I3(commutation_state[2]), .O(n27236));
    defparam i49193_4_lut.LUT_INIT = 16'hc5cf;
    SB_DFFESR delay_counter__i13 (.Q(delay_counter[13]), .C(clk16MHz), .E(n27321), 
            .D(n1232), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n48511), .O(n294)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter__i14 (.Q(delay_counter[14]), .C(clk16MHz), .E(n27321), 
            .D(n1231), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFFESR delay_counter__i15 (.Q(delay_counter[15]), .C(clk16MHz), .E(n27321), 
            .D(n1230), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n2), 
            .I3(n48510), .O(n298)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n48510), .I0(GND_net), .I1(n2), 
            .CO(n48511));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14_adj_5698), 
            .I3(n48509), .O(n299)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n48509), .I0(GND_net), .I1(n14_adj_5698), 
            .CO(n48510));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5699), 
            .I3(n48508), .O(n300)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n48508), .I0(GND_net), .I1(n15_adj_5699), 
            .CO(n48509));
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk16MHz), .D(displacement_23__N_67[23]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk16MHz), .D(displacement_23__N_67[22]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_LUT4 i13398_3_lut (.I0(\data_in_frame[11] [0]), .I1(rx_data[0]), 
            .I2(n55149), .I3(GND_net), .O(n29243));   // verilog/coms.v(130[12] 305[6])
    defparam i13398_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16_adj_5700), 
            .I3(n48507), .O(n301)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n48507), .I0(GND_net), .I1(n16_adj_5700), 
            .CO(n48508));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5701), 
            .I3(n48506), .O(n302)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n48506), .I0(GND_net), .I1(n17_adj_5701), 
            .CO(n48507));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18), 
            .I3(n48505), .O(n303)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n48505), .I0(GND_net), .I1(n18), 
            .CO(n48506));
    SB_LUT4 add_151_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n48270), .O(n1227)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5702), 
            .I3(n48504), .O(n304)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n48504), .I0(GND_net), .I1(n19_adj_5702), 
            .CO(n48505));
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk16MHz), .D(displacement_23__N_67[21]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk16MHz), .D(displacement_23__N_67[20]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk16MHz), .D(displacement_23__N_67[19]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk16MHz), .D(displacement_23__N_67[18]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk16MHz), .D(displacement_23__N_67[17]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk16MHz), .D(displacement_23__N_67[16]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk16MHz), .D(displacement_23__N_67[15]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk16MHz), .D(displacement_23__N_67[14]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk16MHz), .D(displacement_23__N_67[13]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk16MHz), .D(displacement_23__N_67[12]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk16MHz), .D(displacement_23__N_67[11]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk16MHz), .D(displacement_23__N_67[10]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk16MHz), .D(displacement_23__N_67[9]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk16MHz), .D(displacement_23__N_67[8]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk16MHz), .D(displacement_23__N_67[7]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk16MHz), .D(displacement_23__N_67[6]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk16MHz), .D(displacement_23__N_67[5]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk16MHz), .D(displacement_23__N_67[4]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk16MHz), .D(displacement_23__N_67[3]));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    SB_DFFESR delay_counter__i16 (.Q(delay_counter[16]), .C(clk16MHz), .E(n27321), 
            .D(n1229), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_CARRY add_151_20 (.CI(n48270), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n48271));
    SB_LUT4 i13401_3_lut (.I0(\data_in_frame[11] [1]), .I1(rx_data[1]), 
            .I2(n55149), .I3(GND_net), .O(n29246));   // verilog/coms.v(130[12] 305[6])
    defparam i13401_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20_adj_5703), 
            .I3(n48503), .O(n305)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n48503), .I0(GND_net), .I1(n20_adj_5703), 
            .CO(n48504));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21_adj_5704), 
            .I3(n48502), .O(n306)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n48502), .I0(GND_net), .I1(n21_adj_5704), 
            .CO(n48503));
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22_adj_5705), 
            .I3(n48501), .O(n307)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n48501), .I0(GND_net), .I1(n22_adj_5705), 
            .CO(n48502));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5706), 
            .I3(n48500), .O(n308)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13404_3_lut (.I0(\data_in_frame[11] [2]), .I1(rx_data[2]), 
            .I2(n55149), .I3(GND_net), .O(n29249));   // verilog/coms.v(130[12] 305[6])
    defparam i13404_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13407_3_lut (.I0(\data_in_frame[11] [3]), .I1(rx_data[3]), 
            .I2(n55149), .I3(GND_net), .O(n29252));   // verilog/coms.v(130[12] 305[6])
    defparam i13407_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13410_3_lut (.I0(\data_in_frame[11] [4]), .I1(rx_data[4]), 
            .I2(n55149), .I3(GND_net), .O(n29255));   // verilog/coms.v(130[12] 305[6])
    defparam i13410_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i17 (.Q(delay_counter[17]), .C(clk16MHz), .E(n27321), 
            .D(n1228), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFFESR delay_counter__i18 (.Q(delay_counter[18]), .C(clk16MHz), .E(n27321), 
            .D(n1227), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_CARRY unary_minus_16_add_3_4 (.CI(n48500), .I0(GND_net), .I1(n23_adj_5706), 
            .CO(n48501));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5707), 
            .I3(n48499), .O(n309)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF commutation_state_i1 (.Q(commutation_state[1]), .C(clk16MHz), 
           .D(n29574));   // verilog/TinyFPGA_B.v(151[9] 230[5])
    SB_DFF \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(clk16MHz), 
           .D(n53719));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFFESR delay_counter__i19 (.Q(delay_counter[19]), .C(clk16MHz), .E(n27321), 
            .D(n1226), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_CARRY unary_minus_16_add_3_3 (.CI(n48499), .I0(GND_net), .I1(n24_adj_5707), 
            .CO(n48500));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n38659), .I1(GND_net), .I2(n25_adj_5708), 
            .I3(VCC_net), .O(n62960)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_5708), 
            .CO(n48499));
    SB_LUT4 add_151_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n48269), .O(n1228)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13413_3_lut (.I0(\data_in_frame[11] [5]), .I1(rx_data[5]), 
            .I2(n55149), .I3(GND_net), .O(n29258));   // verilog/coms.v(130[12] 305[6])
    defparam i13413_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter__i20 (.Q(delay_counter[20]), .C(clk16MHz), .E(n27321), 
            .D(n1225), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFFESR delay_counter__i21 (.Q(delay_counter[21]), .C(clk16MHz), .E(n27321), 
            .D(n1224), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFFESR delay_counter__i22 (.Q(delay_counter[22]), .C(clk16MHz), .E(n27321), 
            .D(n1223), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFFESR delay_counter__i23 (.Q(delay_counter[23]), .C(clk16MHz), .E(n27321), 
            .D(n1222), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFFESR delay_counter__i24 (.Q(delay_counter[24]), .C(clk16MHz), .E(n27321), 
            .D(n1221), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFFESR delay_counter__i25 (.Q(delay_counter[25]), .C(clk16MHz), .E(n27321), 
            .D(n1220), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFFESR delay_counter__i26 (.Q(delay_counter[26]), .C(clk16MHz), .E(n27321), 
            .D(n1219), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFFESR delay_counter__i27 (.Q(delay_counter[27]), .C(clk16MHz), .E(n27321), 
            .D(n1218), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFFESR delay_counter__i28 (.Q(delay_counter[28]), .C(clk16MHz), .E(n27321), 
            .D(n1217), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFFESR delay_counter__i29 (.Q(delay_counter[29]), .C(clk16MHz), .E(n27321), 
            .D(n1216), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFFESR delay_counter__i30 (.Q(delay_counter[30]), .C(clk16MHz), .E(n27321), 
            .D(n1215), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_DFFESR delay_counter__i31 (.Q(delay_counter[31]), .C(clk16MHz), .E(n27321), 
            .D(n1214), .R(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    SB_LUT4 i13179_3_lut (.I0(\data_in_frame[6] [7]), .I1(rx_data[7]), .I2(n27904), 
            .I3(GND_net), .O(n29024));   // verilog/coms.v(130[12] 305[6])
    defparam i13179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13418_3_lut (.I0(\data_in_frame[11] [6]), .I1(rx_data[6]), 
            .I2(n55149), .I3(GND_net), .O(n29263));   // verilog/coms.v(130[12] 305[6])
    defparam i13418_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk16MHz), .D(pwm_setpoint_23__N_3[0]));   // verilog/TinyFPGA_B.v(112[9] 137[5])
    SB_LUT4 i13421_3_lut (.I0(\data_in_frame[11] [7]), .I1(rx_data[7]), 
            .I2(n55149), .I3(GND_net), .O(n29266));   // verilog/coms.v(130[12] 305[6])
    defparam i13421_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13424_3_lut (.I0(\data_in_frame[12] [0]), .I1(rx_data[0]), 
            .I2(n55151), .I3(GND_net), .O(n29269));   // verilog/coms.v(130[12] 305[6])
    defparam i13424_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13427_3_lut (.I0(\data_in_frame[12] [1]), .I1(rx_data[1]), 
            .I2(n55151), .I3(GND_net), .O(n29272));   // verilog/coms.v(130[12] 305[6])
    defparam i13427_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13430_3_lut (.I0(\data_in_frame[12] [2]), .I1(rx_data[2]), 
            .I2(n55151), .I3(GND_net), .O(n29275));   // verilog/coms.v(130[12] 305[6])
    defparam i13430_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_151_19 (.CI(n48269), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n48270));
    SB_CARRY add_151_8 (.CI(n48258), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n48259));
    SB_LUT4 i13433_3_lut (.I0(\data_in_frame[12] [3]), .I1(rx_data[3]), 
            .I2(n55151), .I3(GND_net), .O(n29278));   // verilog/coms.v(130[12] 305[6])
    defparam i13433_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_151_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n48268), .O(n1229)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2_adj_5760), .I3(n48429), .O(displacement_23__N_67[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_5759), .I3(n48428), .O(displacement_23__N_67[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n48428), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_5759), .CO(n48429));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5758), .I3(n48427), .O(displacement_23__N_67[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n48427), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5758), .CO(n48428));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5776), .I3(n48426), .O(displacement_23__N_67[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n48426), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5776), .CO(n48427));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5775), .I3(n48425), .O(displacement_23__N_67[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n48425), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5775), .CO(n48426));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5774), .I3(n48424), .O(displacement_23__N_67[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n48424), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5774), .CO(n48425));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5773), .I3(n48423), .O(displacement_23__N_67[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_18 (.CI(n48268), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n48269));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n48423), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5773), .CO(n48424));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5772), .I3(n48422), .O(displacement_23__N_67[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n48422), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5772), .CO(n48423));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5757), .I3(n48421), .O(displacement_23__N_67[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n48421), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5757), .CO(n48422));
    SB_LUT4 add_151_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n48267), .O(n1230)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5756), .I3(n48420), .O(displacement_23__N_67[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n48420), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5756), .CO(n48421));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5755), .I3(n48419), .O(displacement_23__N_67[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n48419), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5755), .CO(n48420));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5697), .I3(n48418), .O(displacement_23__N_67[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n48418), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5697), .CO(n48419));
    SB_LUT4 add_151_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n48257), .O(n1240)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_17 (.CI(n48267), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n48268));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14), .I3(n48417), .O(displacement_23__N_67[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n48417), .I0(encoder0_position_scaled[11]), 
            .I1(n14), .CO(n48418));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5696), .I3(n48416), .O(displacement_23__N_67[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n48416), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5696), .CO(n48417));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5695), .I3(n48415), .O(displacement_23__N_67[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n48415), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5695), .CO(n48416));
    SB_CARRY add_151_7 (.CI(n48257), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n48258));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5694), .I3(n48414), .O(displacement_23__N_67[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n48414), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5694), .CO(n48415));
    SB_LUT4 add_151_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n48266), .O(n1231)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1245)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n35729), .I3(n48413), .O(displacement_23__N_67[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n48256), .O(n1241)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_16 (.CI(n48266), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n48267));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n48413), .I0(encoder0_position_scaled[7]), 
            .I1(n35729), .CO(n48414));
    SB_LUT4 add_151_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n48265), .O(n1232)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19), .I3(n48412), .O(displacement_23__N_67[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_15 (.CI(n48265), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n48266));
    SB_CARRY add_151_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n48253));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n48412), .I0(encoder0_position_scaled[6]), 
            .I1(n19), .CO(n48413));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20), .I3(n48411), .O(displacement_23__N_67[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n48411), .I0(encoder0_position_scaled[5]), 
            .I1(n20), .CO(n48412));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21_adj_5692), .I3(n48410), .O(displacement_23__N_67[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_151_6 (.CI(n48256), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n48257));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n48410), .I0(encoder0_position_scaled[4]), 
            .I1(n21_adj_5692), .CO(n48411));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22), .I3(n48409), .O(displacement_23__N_67[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_151_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n48264), .O(n1233)) /* synthesis syn_instantiated=1 */ ;
    defparam add_151_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n48409), .I0(encoder0_position_scaled[3]), 
            .I1(n22), .CO(n48410));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23_adj_5691), .I3(n48408), .O(displacement_23__N_67[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49751 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(byte_transmit_counter[1]), .O(n66861));
    defparam byte_transmit_counter_0__bdd_4_lut_49751.LUT_INIT = 16'he4aa;
    SB_LUT4 n66861_bdd_4_lut (.I0(n66861), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(byte_transmit_counter[1]), 
            .O(n66864));
    defparam n66861_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13437_3_lut (.I0(\data_in_frame[12] [4]), .I1(rx_data[4]), 
            .I2(n55151), .I3(GND_net), .O(n29282));   // verilog/coms.v(130[12] 305[6])
    defparam i13437_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13440_3_lut (.I0(\data_in_frame[12] [5]), .I1(rx_data[5]), 
            .I2(n55151), .I3(GND_net), .O(n29285));   // verilog/coms.v(130[12] 305[6])
    defparam i13440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13443_3_lut (.I0(\data_in_frame[12] [6]), .I1(rx_data[6]), 
            .I2(n55151), .I3(GND_net), .O(n29288));   // verilog/coms.v(130[12] 305[6])
    defparam i13443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11_2_lut (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[3] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n25490));   // verilog/coms.v(99[12:25])
    defparam i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13446_3_lut (.I0(\data_in_frame[12] [7]), .I1(rx_data[7]), 
            .I2(n55151), .I3(GND_net), .O(n29291));   // verilog/coms.v(130[12] 305[6])
    defparam i13446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_1736 (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[1] [4]), 
            .I2(n56216), .I3(n56062), .O(n55681));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1736.LUT_INIT = 16'h6996;
    SB_LUT4 i13449_3_lut (.I0(\data_in_frame[13] [0]), .I1(rx_data[0]), 
            .I2(n55153), .I3(GND_net), .O(n29294));   // verilog/coms.v(130[12] 305[6])
    defparam i13449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13452_3_lut (.I0(\data_in_frame[13] [1]), .I1(rx_data[1]), 
            .I2(n55153), .I3(GND_net), .O(n29297));   // verilog/coms.v(130[12] 305[6])
    defparam i13452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1737 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5829));
    defparam i1_2_lut_adj_1737.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut (.I0(delay_counter[9]), .I1(n4_adj_5829), .I2(delay_counter[10]), 
            .I3(n24969), .O(n58172));
    defparam i2_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1738 (.I0(n58172), .I1(n24966), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n57520));
    defparam i2_4_lut_adj_1738.LUT_INIT = 16'hffec;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_5823));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut_adj_1739 (.I0(delay_counter[22]), .I1(n57520), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5824));
    defparam i2_4_lut_adj_1739.LUT_INIT = 16'ha8a0;
    SB_LUT4 i22486_4_lut (.I0(n7_adj_5824), .I1(delay_counter[31]), .I2(n24971), 
            .I3(n8_adj_5823), .O(n1325));   // verilog/TinyFPGA_B.v(388[14:38])
    defparam i22486_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i5_4_lut_adj_1740 (.I0(delay_counter[27]), .I1(delay_counter[29]), 
            .I2(delay_counter[24]), .I3(delay_counter[26]), .O(n12_adj_5840));
    defparam i5_4_lut_adj_1740.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1741 (.I0(delay_counter[28]), .I1(n12_adj_5840), 
            .I2(delay_counter[25]), .I3(delay_counter[30]), .O(n24971));
    defparam i6_4_lut_adj_1741.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1742 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n24966));
    defparam i2_3_lut_adj_1742.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_3_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n14_adj_5822));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1743 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15_adj_5821));
    defparam i6_4_lut_adj_1743.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5821), .I1(delay_counter[2]), .I2(n14_adj_5822), 
            .I3(delay_counter[6]), .O(n24969));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4290_4_lut (.I0(n24969), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5709));
    defparam i4290_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut_adj_1744 (.I0(n24_adj_5709), .I1(delay_counter[14]), 
            .I2(delay_counter[12]), .I3(delay_counter[13]), .O(n57982));
    defparam i2_4_lut_adj_1744.LUT_INIT = 16'hc800;
    SB_LUT4 i2_3_lut_adj_1745 (.I0(n57982), .I1(delay_counter[18]), .I2(n24966), 
            .I3(GND_net), .O(n57716));
    defparam i2_3_lut_adj_1745.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_1746 (.I0(delay_counter[23]), .I1(n57716), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7_adj_5796));
    defparam i2_4_lut_adj_1746.LUT_INIT = 16'heaaa;
    SB_LUT4 i4_4_lut (.I0(n7_adj_5796), .I1(delay_counter[21]), .I2(delay_counter[22]), 
            .I3(n24971), .O(n62));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22538_2_lut (.I0(n62), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_409));   // verilog/TinyFPGA_B.v(374[12:35])
    defparam i22538_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12795_4_lut (.I0(n27321), .I1(n1325), .I2(n63020), .I3(n38279), 
            .O(n28611));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i12795_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i13455_3_lut (.I0(\data_in_frame[13] [2]), .I1(rx_data[2]), 
            .I2(n55153), .I3(GND_net), .O(n29300));   // verilog/coms.v(130[12] 305[6])
    defparam i13455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13458_3_lut (.I0(\data_in_frame[13] [3]), .I1(rx_data[3]), 
            .I2(n55153), .I3(GND_net), .O(n29303));   // verilog/coms.v(130[12] 305[6])
    defparam i13458_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13461_3_lut (.I0(\data_in_frame[13] [4]), .I1(rx_data[4]), 
            .I2(n55153), .I3(GND_net), .O(n29306));   // verilog/coms.v(130[12] 305[6])
    defparam i13461_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13464_3_lut (.I0(\data_in_frame[13] [5]), .I1(rx_data[5]), 
            .I2(n55153), .I3(GND_net), .O(n29309));   // verilog/coms.v(130[12] 305[6])
    defparam i13464_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13468_3_lut (.I0(\data_in_frame[13] [6]), .I1(rx_data[6]), 
            .I2(n55153), .I3(GND_net), .O(n29313));   // verilog/coms.v(130[12] 305[6])
    defparam i13468_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i42993_3_lut (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[7] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60055));
    defparam i42993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42994_4_lut (.I0(n60055), .I1(n27513), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n60056));
    defparam i42994_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i42992_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60054));
    defparam i42992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46320_2_lut (.I0(n66702), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n63131));
    defparam i46320_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13471_3_lut (.I0(\data_in_frame[13] [7]), .I1(rx_data[7]), 
            .I2(n55153), .I3(GND_net), .O(n29316));   // verilog/coms.v(130[12] 305[6])
    defparam i13471_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13167_3_lut (.I0(\data_in_frame[6] [3]), .I1(rx_data[3]), .I2(n27904), 
            .I3(GND_net), .O(n29012));   // verilog/coms.v(130[12] 305[6])
    defparam i13167_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5692));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1747 (.I0(n23_adj_5830), .I1(o_Rx_DV_N_3488[12]), 
            .I2(n5228), .I3(GND_net), .O(n58452));
    defparam i1_3_lut_adj_1747.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut (.I0(o_Rx_DV_N_3488[24]), .I1(n27), .I2(n29), .I3(n58452), 
            .O(n39937));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1748 (.I0(o_Rx_DV_N_3488[12]), .I1(n5228), .I2(n31), 
            .I3(GND_net), .O(n58600));
    defparam i1_3_lut_adj_1748.LUT_INIT = 16'hefef;
    SB_LUT4 i1_4_lut_adj_1749 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5830), 
            .I3(n58600), .O(n58606));
    defparam i1_4_lut_adj_1749.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1750 (.I0(r_SM_Main_2__N_3545[0]), .I1(n58606), 
            .I2(r_SM_Main_adj_5922[1]), .I3(n27), .O(n9_adj_5710));   // verilog/uart_tx.v(32[16:25])
    defparam i13_4_lut_adj_1750.LUT_INIT = 16'h0a3a;
    SB_LUT4 i14_3_lut (.I0(n9_adj_5710), .I1(n39937), .I2(r_SM_Main_adj_5922[0]), 
            .I3(GND_net), .O(n20722));   // verilog/uart_tx.v(32[16:25])
    defparam i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24232_3_lut (.I0(r_SM_Main_adj_5922[0]), .I1(o_Tx_Serial_N_3598), 
            .I2(r_SM_Main_adj_5922[1]), .I3(GND_net), .O(n39972));   // verilog/uart_tx.v(32[16:25])
    defparam i24232_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i19941_1_lut (.I0(encoder1_position_scaled[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n35729));   // verilog/TinyFPGA_B.v(329[10] 333[6])
    defparam i19941_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5694));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5695));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[11]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i12_3_lut (.I0(encoder0_position_scaled[11]), .I1(motor_state_23__N_91[11]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5696));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[12]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i13_3_lut (.I0(encoder0_position_scaled[12]), .I1(motor_state_23__N_91[12]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[13]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i14_3_lut (.I0(encoder0_position_scaled[13]), .I1(motor_state_23__N_91[13]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5697));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(n8));
    defparam i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i10_3_lut (.I0(encoder0_position_scaled[14]), .I1(n8), .I2(n15_adj_5748), 
            .I3(GND_net), .O(n9_adj_5792));
    defparam i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5755));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_4_lut_adj_1751 (.I0(n51197), .I1(n50927), .I2(n56024), 
            .I3(n51232), .O(n18_adj_5794));
    defparam i7_4_lut_adj_1751.LUT_INIT = 16'h6996;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5756));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[15]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i5_2_lut (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[21] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_5795));
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_243_i16_3_lut (.I0(encoder0_position_scaled[15]), .I1(motor_state_23__N_91[15]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5757));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9_4_lut_adj_1752 (.I0(\data_out_frame[23] [2]), .I1(n18_adj_5794), 
            .I2(n50183), .I3(n56231), .O(n20_adj_5793));
    defparam i9_4_lut_adj_1752.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut (.I0(n56201), .I1(n20_adj_5793), .I2(n16_adj_5795), 
            .I3(n55989), .O(n50946));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mux_245_i17_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[16]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i17_3_lut (.I0(encoder0_position_scaled[16]), .I1(motor_state_23__N_91[16]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5772));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[17]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i18_3_lut (.I0(encoder0_position_scaled[17]), .I1(motor_state_23__N_91[17]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_245_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[18]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i19_3_lut (.I0(encoder0_position_scaled[18]), .I1(motor_state_23__N_91[18]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5773));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_2));   // verilog/TinyFPGA_B.v(270[11:14])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5774));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[19]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i20_3_lut (.I0(encoder0_position_scaled[19]), .I1(motor_state_23__N_91[19]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5775));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[20]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i21_3_lut (.I0(encoder0_position_scaled[20]), .I1(motor_state_23__N_91[20]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49606 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[20] [7]), .I2(\data_out_frame[21] [7]), 
            .I3(byte_transmit_counter[2]), .O(n66669));
    defparam byte_transmit_counter_0__bdd_4_lut_49606.LUT_INIT = 16'he4aa;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5776));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_245_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[21]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i22_3_lut (.I0(encoder0_position_scaled[21]), .I1(motor_state_23__N_91[21]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5758));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1753 (.I0(n23_adj_5830), .I1(o_Rx_DV_N_3488[12]), 
            .I2(n5225), .I3(o_Rx_DV_N_3488[8]), .O(n58462));
    defparam i1_4_lut_adj_1753.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_245_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[22]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i23_3_lut (.I0(encoder0_position_scaled[22]), .I1(motor_state_23__N_91[22]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_4_lut_adj_1754 (.I0(o_Rx_DV_N_3488[24]), .I1(n27), .I2(n29), 
            .I3(n58462), .O(r_SM_Main_2__N_3446[1]));
    defparam i1_4_lut_adj_1754.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_245_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[23]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i24_3_lut (.I0(encoder0_position_scaled[23]), .I1(motor_state_23__N_91[23]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i24_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5759));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5760));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_1178_i9_2_lut (.I0(r_Clock_Count[4]), .I1(o_Rx_DV_N_3488[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5808));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5123_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_400));   // verilog/TinyFPGA_B.v(208[7] 227[14])
    defparam i5123_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 i5121_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_391));   // verilog/TinyFPGA_B.v(208[7] 227[14])
    defparam i5121_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 LessThan_1178_i4_4_lut (.I0(r_Clock_Count[0]), .I1(o_Rx_DV_N_3488[1]), 
            .I2(r_Clock_Count[1]), .I3(o_Rx_DV_N_3488[0]), .O(n4_adj_5805));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 LessThan_1178_i8_3_lut (.I0(n6_adj_5806), .I1(o_Rx_DV_N_3488[4]), 
            .I2(n9_adj_5808), .I3(GND_net), .O(n8_adj_5807));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49039_4_lut (.I0(n8_adj_5807), .I1(n4_adj_5805), .I2(n9_adj_5808), 
            .I3(n63426), .O(n66101));   // verilog/uart_rx.v(119[17:57])
    defparam i49039_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47092_2_lut (.I0(n66714), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n63134));
    defparam i47092_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49040_3_lut (.I0(n66101), .I1(o_Rx_DV_N_3488[5]), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n66102));   // verilog/uart_rx.v(119[17:57])
    defparam i49040_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48940_3_lut (.I0(n66102), .I1(o_Rx_DV_N_3488[6]), .I2(r_Clock_Count[6]), 
            .I3(GND_net), .O(n66002));   // verilog/uart_rx.v(119[17:57])
    defparam i48940_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48760_3_lut (.I0(n66002), .I1(o_Rx_DV_N_3488[7]), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(n5225));   // verilog/uart_rx.v(119[17:57])
    defparam i48760_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_4_lut_adj_1755 (.I0(o_Rx_DV_N_3488[12]), .I1(n5225), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n55184), .O(n58612));
    defparam i1_4_lut_adj_1755.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_1756 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5830), 
            .I3(n58612), .O(n58618));
    defparam i1_4_lut_adj_1756.LUT_INIT = 16'hfffe;
    SB_LUT4 i46399_3_lut_4_lut (.I0(r_Clock_Count_adj_5923[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count_adj_5923[2]), .O(n63461));   // verilog/uart_tx.v(117[17:57])
    defparam i46399_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_1181_i6_3_lut_3_lut (.I0(r_Clock_Count_adj_5923[3]), 
            .I1(o_Rx_DV_N_3488[3]), .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), 
            .O(n6_adj_5798));   // verilog/uart_tx.v(117[17:57])
    defparam LessThan_1181_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i39361_2_lut_3_lut (.I0(n3484), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n56368));
    defparam i39361_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 mux_245_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[8]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i9_3_lut (.I0(encoder0_position_scaled[8]), .I1(motor_state_23__N_91[8]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13065_3_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(n359), 
            .I2(n27260), .I3(GND_net), .O(n28910));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13158_3_lut (.I0(\data_in_frame[6] [0]), .I1(rx_data[0]), .I2(n27904), 
            .I3(GND_net), .O(n29003));   // verilog/coms.v(130[12] 305[6])
    defparam i13158_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13155_3_lut (.I0(\data_in_frame[5] [7]), .I1(rx_data[7]), .I2(n27902), 
            .I3(GND_net), .O(n29000));   // verilog/coms.v(130[12] 305[6])
    defparam i13155_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut (.I0(n15_adj_5741), .I1(n22471), .I2(dti), 
            .I3(GND_net), .O(n27212));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hbaba;
    SB_LUT4 i13076_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n22369), .I3(GND_net), .O(n28921));   // verilog/coms.v(130[12] 305[6])
    defparam i13076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13077_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n22318), .I3(GND_net), .O(n28922));   // verilog/coms.v(130[12] 305[6])
    defparam i13077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13078_3_lut (.I0(current_limit[0]), .I1(\data_in_frame[21] [0]), 
            .I2(n22318), .I3(GND_net), .O(n28923));   // verilog/coms.v(130[12] 305[6])
    defparam i13078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13152_3_lut (.I0(\data_in_frame[5] [6]), .I1(rx_data[6]), .I2(n27902), 
            .I3(GND_net), .O(n28997));   // verilog/coms.v(130[12] 305[6])
    defparam i13152_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13149_3_lut (.I0(\data_in_frame[5] [5]), .I1(rx_data[5]), .I2(n27902), 
            .I3(GND_net), .O(n28994));   // verilog/coms.v(130[12] 305[6])
    defparam i13149_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13080_3_lut (.I0(ID[0]), .I1(data_adj_5899[0]), .I2(n55524), 
            .I3(GND_net), .O(n28925));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13080_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13146_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n27902), 
            .I3(GND_net), .O(n28991));   // verilog/coms.v(130[12] 305[6])
    defparam i13146_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13143_3_lut (.I0(\data_in_frame[5] [3]), .I1(rx_data[3]), .I2(n27902), 
            .I3(GND_net), .O(n28988));   // verilog/coms.v(130[12] 305[6])
    defparam i13143_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13082_3_lut (.I0(current[0]), .I1(data_adj_5906[0]), .I2(n27290), 
            .I3(GND_net), .O(n28927));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1757 (.I0(n4_adj_5836), .I1(\data_out_frame[16] [4]), 
            .I2(n26439), .I3(n25803), .O(n10_adj_5837));
    defparam i4_4_lut_adj_1757.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5922[1]), .I2(n58502), 
            .I3(n39919), .O(n51433));   // verilog/uart_tx.v(32[16:25])
    defparam i12_4_lut.LUT_INIT = 16'h3aba;
    SB_LUT4 i13137_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n27902), 
            .I3(GND_net), .O(n28982));   // verilog/coms.v(130[12] 305[6])
    defparam i13137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1758 (.I0(r_SM_Main[1]), .I1(n6_adj_5838), .I2(r_Bit_Index[0]), 
            .I3(n4_adj_5744), .O(n58862));
    defparam i1_4_lut_adj_1758.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_4_lut_adj_1759 (.I0(o_Rx_DV_N_3488[12]), .I1(n5225), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n58862), .O(n58868));
    defparam i1_4_lut_adj_1759.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1760 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5830), 
            .I3(n58868), .O(n58874));
    defparam i1_4_lut_adj_1760.LUT_INIT = 16'hfffe;
    SB_LUT4 i13730_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n58874), 
            .I3(n27), .O(n29575));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13730_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1761 (.I0(o_Rx_DV_N_3488[12]), .I1(n5225), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n58880), .O(n58886));
    defparam i1_4_lut_adj_1761.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1762 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5830), 
            .I3(n58886), .O(n58892));
    defparam i1_4_lut_adj_1762.LUT_INIT = 16'hfffe;
    SB_LUT4 i13731_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n58892), 
            .I3(n27), .O(n29576));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13731_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_1677_i17_3_lut (.I0(duty[19]), .I1(duty[16]), .I2(n260), 
            .I3(GND_net), .O(n11598));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_4_lut_adj_1763 (.I0(o_Rx_DV_N_3488[12]), .I1(n5225), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n58952), .O(n58958));
    defparam i1_4_lut_adj_1763.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1764 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5830), 
            .I3(n58958), .O(n58964));
    defparam i1_4_lut_adj_1764.LUT_INIT = 16'hfffe;
    SB_LUT4 i13732_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n58964), 
            .I3(n27), .O(n29577));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13732_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1765 (.I0(o_Rx_DV_N_3488[12]), .I1(n5225), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n58970), .O(n58976));
    defparam i1_4_lut_adj_1765.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1766 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5830), 
            .I3(n58976), .O(n58982));
    defparam i1_4_lut_adj_1766.LUT_INIT = 16'hfffe;
    SB_LUT4 i13733_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n58982), 
            .I3(n27), .O(n29578));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13733_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i2_3_lut_4_lut (.I0(n3484), .I1(\FRAME_MATCHER.i [5]), .I2(n8_adj_5711), 
            .I3(n73), .O(n67));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i1_4_lut_adj_1767 (.I0(o_Rx_DV_N_3488[12]), .I1(n5225), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n58934), .O(n58940));
    defparam i1_4_lut_adj_1767.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1768 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5830), 
            .I3(n58940), .O(n58946));
    defparam i1_4_lut_adj_1768.LUT_INIT = 16'hfffe;
    SB_LUT4 i13735_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n58946), 
            .I3(n27), .O(n29580));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13735_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_1677_i18_3_lut (.I0(duty[20]), .I1(duty[17]), .I2(n260), 
            .I3(GND_net), .O(n11596));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_4_lut_adj_1769 (.I0(o_Rx_DV_N_3488[12]), .I1(n5225), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n58898), .O(n58904));
    defparam i1_4_lut_adj_1769.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1770 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5830), 
            .I3(n58904), .O(n58910));
    defparam i1_4_lut_adj_1770.LUT_INIT = 16'hfffe;
    SB_LUT4 i13736_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n58910), 
            .I3(n27), .O(n29581));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13736_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1771 (.I0(o_Rx_DV_N_3488[12]), .I1(n5225), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n58844), .O(n58850));
    defparam i1_4_lut_adj_1771.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1772 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5830), 
            .I3(n58850), .O(n58856));
    defparam i1_4_lut_adj_1772.LUT_INIT = 16'hfffe;
    SB_LUT4 i13737_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n58856), 
            .I3(n27), .O(n29582));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13737_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13093_3_lut (.I0(b_prev_adj_5752), .I1(b_new_adj_5886[1]), 
            .I2(debounce_cnt_N_3833_adj_5753), .I3(GND_net), .O(n28938));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13093_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13094_3_lut (.I0(t0[0]), .I1(timer[0]), .I2(n3173), .I3(GND_net), 
            .O(n28939));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13094_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46404_3_lut (.I0(state_7__N_4110[0]), .I1(n38221), .I2(enable_slow_N_4213), 
            .I3(GND_net), .O(n63151));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i46404_3_lut.LUT_INIT = 16'h4c4c;
    SB_LUT4 i14_4_lut (.I0(n63151), .I1(state_adj_5935[0]), .I2(n6715), 
            .I3(n38223), .O(n6_adj_5842));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14_4_lut.LUT_INIT = 16'h5cfc;
    SB_LUT4 i13131_3_lut (.I0(\data_in_frame[4] [7]), .I1(rx_data[7]), .I2(n27900), 
            .I3(GND_net), .O(n28976));   // verilog/coms.v(130[12] 305[6])
    defparam i13131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13741_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5899[0]), 
            .I2(n10_adj_5812), .I3(n25100), .O(n29586));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13741_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_1677_i19_3_lut (.I0(duty[21]), .I1(duty[18]), .I2(n260), 
            .I3(GND_net), .O(n11594));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_4_lut_adj_1773 (.I0(n4_adj_5744), .I1(r_SM_Main[1]), .I2(n6_adj_5838), 
            .I3(r_Bit_Index[0]), .O(n58916));
    defparam i1_4_lut_adj_1773.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_4_lut_adj_1774 (.I0(o_Rx_DV_N_3488[12]), .I1(n5225), .I2(o_Rx_DV_N_3488[8]), 
            .I3(n58916), .O(n58922));
    defparam i1_4_lut_adj_1774.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1775 (.I0(o_Rx_DV_N_3488[24]), .I1(n29), .I2(n23_adj_5830), 
            .I3(n58922), .O(n58928));
    defparam i1_4_lut_adj_1775.LUT_INIT = 16'hfffe;
    SB_LUT4 i13751_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n58928), 
            .I3(n27), .O(n29596));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13751_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13755_4_lut (.I0(CS_MISO_c), .I1(data_adj_5906[0]), .I2(n11_adj_5747), 
            .I3(state_7__N_4319), .O(n29600));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13755_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13122_3_lut (.I0(\data_in_frame[4] [4]), .I1(rx_data[4]), .I2(n27900), 
            .I3(GND_net), .O(n28967));   // verilog/coms.v(130[12] 305[6])
    defparam i13122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_1677_i20_3_lut (.I0(duty[22]), .I1(duty[19]), .I2(n260), 
            .I3(GND_net), .O(n11592));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13787_3_lut (.I0(current_limit[15]), .I1(\data_in_frame[20] [7]), 
            .I2(n22318), .I3(GND_net), .O(n29632));   // verilog/coms.v(130[12] 305[6])
    defparam i13787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14168_2_lut_4_lut (.I0(reset), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2882));   // verilog/coms.v(130[12] 305[6])
    defparam i14168_2_lut_4_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(current[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5708));   // verilog/TinyFPGA_B.v(129[16:24])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13788_3_lut (.I0(current_limit[14]), .I1(\data_in_frame[20] [6]), 
            .I2(n22318), .I3(GND_net), .O(n29633));   // verilog/coms.v(130[12] 305[6])
    defparam i13788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13789_3_lut (.I0(current_limit[13]), .I1(\data_in_frame[20] [5]), 
            .I2(n22318), .I3(GND_net), .O(n29634));   // verilog/coms.v(130[12] 305[6])
    defparam i13789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13790_3_lut (.I0(current_limit[12]), .I1(\data_in_frame[20] [4]), 
            .I2(n22318), .I3(GND_net), .O(n29635));   // verilog/coms.v(130[12] 305[6])
    defparam i13790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13791_3_lut (.I0(current_limit[11]), .I1(\data_in_frame[20] [3]), 
            .I2(n22318), .I3(GND_net), .O(n29636));   // verilog/coms.v(130[12] 305[6])
    defparam i13791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13792_3_lut (.I0(current_limit[10]), .I1(\data_in_frame[20] [2]), 
            .I2(n22318), .I3(GND_net), .O(n29637));   // verilog/coms.v(130[12] 305[6])
    defparam i13792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13793_3_lut (.I0(current_limit[9]), .I1(\data_in_frame[20] [1]), 
            .I2(n22318), .I3(GND_net), .O(n29638));   // verilog/coms.v(130[12] 305[6])
    defparam i13793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13795_3_lut (.I0(current_limit[7]), .I1(\data_in_frame[21] [7]), 
            .I2(n22318), .I3(GND_net), .O(n29640));   // verilog/coms.v(130[12] 305[6])
    defparam i13795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13797_3_lut (.I0(current_limit[5]), .I1(\data_in_frame[21] [5]), 
            .I2(n22318), .I3(GND_net), .O(n29642));   // verilog/coms.v(130[12] 305[6])
    defparam i13797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13798_3_lut (.I0(current_limit[4]), .I1(\data_in_frame[21] [4]), 
            .I2(n22318), .I3(GND_net), .O(n29643));   // verilog/coms.v(130[12] 305[6])
    defparam i13798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13799_3_lut (.I0(current_limit[3]), .I1(\data_in_frame[21] [3]), 
            .I2(n22318), .I3(GND_net), .O(n29644));   // verilog/coms.v(130[12] 305[6])
    defparam i13799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13800_3_lut (.I0(current_limit[2]), .I1(\data_in_frame[21] [2]), 
            .I2(n22318), .I3(GND_net), .O(n29645));   // verilog/coms.v(130[12] 305[6])
    defparam i13800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13801_3_lut (.I0(current_limit[1]), .I1(\data_in_frame[21] [1]), 
            .I2(n22318), .I3(GND_net), .O(n29646));   // verilog/coms.v(130[12] 305[6])
    defparam i13801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18753_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n22318), .I3(GND_net), .O(n29647));
    defparam i18753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13803_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n22318), .I3(GND_net), .O(n29648));   // verilog/coms.v(130[12] 305[6])
    defparam i13803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13804_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n22318), .I3(GND_net), .O(n29649));   // verilog/coms.v(130[12] 305[6])
    defparam i13804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13805_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n22318), .I3(GND_net), .O(n29650));   // verilog/coms.v(130[12] 305[6])
    defparam i13805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [0]), 
            .O(n55454));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h5100;
    SB_LUT4 i13809_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n22369), .I3(GND_net), .O(n29654));   // verilog/coms.v(130[12] 305[6])
    defparam i13809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1776 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [1]), 
            .O(n55453));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1776.LUT_INIT = 16'h5100;
    SB_LUT4 i13810_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n22369), .I3(GND_net), .O(n29655));   // verilog/coms.v(130[12] 305[6])
    defparam i13810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13811_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n22369), .I3(GND_net), .O(n29656));   // verilog/coms.v(130[12] 305[6])
    defparam i13811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13812_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n22369), .I3(GND_net), .O(n29657));   // verilog/coms.v(130[12] 305[6])
    defparam i13812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1777 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [2]), 
            .O(n55452));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1777.LUT_INIT = 16'h5100;
    SB_LUT4 i13815_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n22369), .I3(GND_net), .O(n29660));   // verilog/coms.v(130[12] 305[6])
    defparam i13815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18721_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n22369), .I3(GND_net), .O(n29661));
    defparam i18721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13817_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n22369), .I3(GND_net), .O(n29662));   // verilog/coms.v(130[12] 305[6])
    defparam i13817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13819_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n22369), .I3(GND_net), .O(n29664));   // verilog/coms.v(130[12] 305[6])
    defparam i13819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13820_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n22369), .I3(GND_net), .O(n29665));   // verilog/coms.v(130[12] 305[6])
    defparam i13820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13821_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n22369), .I3(GND_net), .O(n29666));   // verilog/coms.v(130[12] 305[6])
    defparam i13821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13822_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n22369), .I3(GND_net), .O(n29667));   // verilog/coms.v(130[12] 305[6])
    defparam i13822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13823_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n22369), .I3(GND_net), .O(n29668));   // verilog/coms.v(130[12] 305[6])
    defparam i13823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13824_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n22369), .I3(GND_net), .O(n29669));   // verilog/coms.v(130[12] 305[6])
    defparam i13824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13825_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n22369), .I3(GND_net), .O(n29670));   // verilog/coms.v(130[12] 305[6])
    defparam i13825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13826_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n22369), .I3(GND_net), .O(n29671));   // verilog/coms.v(130[12] 305[6])
    defparam i13826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13828_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n22369), .I3(GND_net), .O(n29673));   // verilog/coms.v(130[12] 305[6])
    defparam i13828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13829_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n22369), .I3(GND_net), .O(n29674));   // verilog/coms.v(130[12] 305[6])
    defparam i13829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13116_3_lut (.I0(\data_in_frame[4] [2]), .I1(rx_data[2]), .I2(n27900), 
            .I3(GND_net), .O(n28961));   // verilog/coms.v(130[12] 305[6])
    defparam i13116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13831_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n22369), .I3(GND_net), .O(n29676));   // verilog/coms.v(130[12] 305[6])
    defparam i13831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13832_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n22369), .I3(GND_net), .O(n29677));   // verilog/coms.v(130[12] 305[6])
    defparam i13832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1778 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [3]), 
            .O(n55451));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1778.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1779 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [4]), 
            .O(n55450));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1779.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1780 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [5]), 
            .O(n55445));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1780.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1781 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [6]), 
            .O(n28680));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1781.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1782 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[26] [7]), 
            .O(n55455));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1782.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1783 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [0]), 
            .O(n55446));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1783.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1784 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [1]), 
            .O(n55447));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1784.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1785 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [2]), 
            .O(n55448));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1785.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1786 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [3]), 
            .O(n55449));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1786.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1787 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [4]), 
            .O(n55443));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1787.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1788 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [5]), 
            .O(n55444));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1788.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1789 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [6]), 
            .O(n28672));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1789.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1790 (.I0(reset), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[27] [7]), 
            .O(n55456));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1790.LUT_INIT = 16'h5100;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[16] [4]), 
            .I2(n10_adj_5745), .I3(n25494), .O(n55766));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13529_3_lut_4_lut_4_lut (.I0(reset), .I1(n67), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n29374));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i13529_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13536_3_lut_4_lut_4_lut (.I0(reset), .I1(n67), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n29381));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i13536_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13539_3_lut_4_lut_4_lut (.I0(reset), .I1(n67), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n29384));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i13539_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13523_3_lut_4_lut_4_lut (.I0(reset), .I1(n67), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n29368));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i13523_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13533_3_lut_4_lut_4_lut (.I0(reset), .I1(n67), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n29378));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i13533_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13526_3_lut_4_lut_4_lut (.I0(reset), .I1(n67), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n29371));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i13526_3_lut_4_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(duty[2]), .I1(duty[3]), .I2(current[3]), 
            .I3(GND_net), .O(n6_adj_5739));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_11_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(current[6]), 
            .I3(GND_net), .O(n10_adj_5735));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam LessThan_11_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_11_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(current[8]), 
            .I3(GND_net), .O(n8_adj_5737));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam LessThan_11_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(reset), .I1(n3484), .I2(n37097), 
            .I3(n8_adj_5789), .O(n27929));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i46326_2_lut_4_lut (.I0(duty[8]), .I1(n302), .I2(duty[4]), 
            .I3(n306), .O(n63388));
    defparam i46326_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i46335_2_lut_4_lut (.I0(duty[6]), .I1(n304), .I2(duty[5]), 
            .I3(n305), .O(n63397));
    defparam i46335_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_14_i6_3_lut_3_lut (.I0(current_limit[2]), .I1(current_limit[3]), 
            .I2(current[3]), .I3(GND_net), .O(n6_adj_5724));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam LessThan_14_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46924_2_lut_4_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(current[4]), .I3(current_limit[4]), .O(n63986));
    defparam i46924_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_14_i8_3_lut_3_lut (.I0(current_limit[4]), .I1(current_limit[8]), 
            .I2(current[8]), .I3(GND_net), .O(n8_adj_5722));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam LessThan_14_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1791 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [1]), 
            .O(n55292));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1791.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1792 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [2]), 
            .O(n55291));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1792.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1793 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [3]), 
            .O(n55290));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1793.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1794 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [4]), 
            .O(n55289));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1794.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1795 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [5]), 
            .O(n55288));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1795.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1796 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [6]), 
            .O(n55242));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1796.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1797 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [7]), 
            .O(n55287));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1797.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1798 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [0]), 
            .O(n55286));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1798.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1799 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [1]), 
            .O(n55285));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1799.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1800 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [2]), 
            .O(n55284));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1800.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1801 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [3]), 
            .O(n55283));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1801.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1802 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [4]), 
            .O(n55282));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1802.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1803 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [1]), 
            .O(n55409));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1803.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1804 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [5]), 
            .O(n55281));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1804.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1805 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [6]), 
            .O(n55280));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1805.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1806 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[19] [7]), 
            .O(n55279));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1806.LUT_INIT = 16'h2300;
    SB_LUT4 mux_1677_i21_3_lut (.I0(duty[23]), .I1(duty[20]), .I2(n260), 
            .I3(GND_net), .O(n11590));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1807 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [0]), 
            .O(n55278));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1807.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1808 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [3]), 
            .O(n55408));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1808.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1809 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [4]), 
            .O(n55407));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1809.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1810 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [1]), 
            .O(n55277));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1810.LUT_INIT = 16'h2300;
    SB_LUT4 i13218_3_lut_4_lut (.I0(n1749), .I1(b_prev), .I2(a_new[1]), 
            .I3(position_31__N_3836), .O(n29063));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13218_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1811 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [6]), 
            .O(n55406));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1811.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1812 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[3] [7]), 
            .O(n55405));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1812.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1813 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [2]), 
            .O(n55276));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1813.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1814 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [3]), 
            .O(n55275));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1814.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1815 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [4]), 
            .O(n55274));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1815.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1816 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [5]), 
            .O(n28729));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1816.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1817 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [6]), 
            .O(n55273));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1817.LUT_INIT = 16'h2300;
    SB_LUT4 i13909_3_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(n336), 
            .I2(n27260), .I3(GND_net), .O(n29754));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13113_3_lut (.I0(\data_in_frame[4] [1]), .I1(rx_data[1]), .I2(n27900), 
            .I3(GND_net), .O(n28958));   // verilog/coms.v(130[12] 305[6])
    defparam i13113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1818 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[20] [7]), 
            .O(n55272));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1818.LUT_INIT = 16'h2300;
    SB_LUT4 i49197_3_lut (.I0(rx_data[0]), .I1(\data_in_frame[4] [0]), .I2(n27900), 
            .I3(GND_net), .O(n54733));   // verilog/coms.v(94[13:20])
    defparam i49197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13912_3_lut (.I0(\PID_CONTROLLER.integral [22]), .I1(n337), 
            .I2(n27260), .I3(GND_net), .O(n29757));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13913_3_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n338), 
            .I2(n27260), .I3(GND_net), .O(n29758));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13914_3_lut (.I0(\PID_CONTROLLER.integral [20]), .I1(n339), 
            .I2(n27260), .I3(GND_net), .O(n29759));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13915_3_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n340), 
            .I2(n27260), .I3(GND_net), .O(n29760));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13916_3_lut (.I0(\PID_CONTROLLER.integral [18]), .I1(n341), 
            .I2(n27260), .I3(GND_net), .O(n29761));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13917_3_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n342), 
            .I2(n27260), .I3(GND_net), .O(n29762));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13918_3_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n343), 
            .I2(n27260), .I3(GND_net), .O(n29763));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13919_3_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n344), 
            .I2(n27260), .I3(GND_net), .O(n29764));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13920_3_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n345), 
            .I2(n27260), .I3(GND_net), .O(n29765));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13921_3_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n346), 
            .I2(n27260), .I3(GND_net), .O(n29766));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13922_3_lut (.I0(\PID_CONTROLLER.integral [12]), .I1(n347), 
            .I2(n27260), .I3(GND_net), .O(n29767));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13923_3_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n348), 
            .I2(n27260), .I3(GND_net), .O(n29768));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13924_3_lut (.I0(\PID_CONTROLLER.integral [10]), .I1(n349), 
            .I2(n27260), .I3(GND_net), .O(n29769));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13925_3_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n350), 
            .I2(n27260), .I3(GND_net), .O(n29770));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13926_3_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(n351), 
            .I2(n27260), .I3(GND_net), .O(n29771));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1819 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [0]), 
            .O(n55271));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1819.LUT_INIT = 16'h2300;
    SB_LUT4 i13927_3_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n352), 
            .I2(n27260), .I3(GND_net), .O(n29772));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13928_3_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(n353), 
            .I2(n27260), .I3(GND_net), .O(n29773));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13929_3_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(n354), 
            .I2(n27260), .I3(GND_net), .O(n29774));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13930_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(n355), 
            .I2(n27260), .I3(GND_net), .O(n29775));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13931_3_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(n356), 
            .I2(n27260), .I3(GND_net), .O(n29776));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13932_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(n357), 
            .I2(n27260), .I3(GND_net), .O(n29777));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13933_3_lut (.I0(\PID_CONTROLLER.integral [1]), .I1(n358), 
            .I2(n27260), .I3(GND_net), .O(n29778));   // verilog/motorControl.v(42[14] 73[8])
    defparam i13933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1820 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [1]), 
            .O(n55270));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1820.LUT_INIT = 16'h2300;
    SB_LUT4 i13107_3_lut (.I0(\data_in_frame[3] [7]), .I1(rx_data[7]), .I2(n27898), 
            .I3(GND_net), .O(n28952));   // verilog/coms.v(130[12] 305[6])
    defparam i13107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13104_3_lut (.I0(\data_in_frame[3] [6]), .I1(rx_data[6]), .I2(n27898), 
            .I3(GND_net), .O(n28949));   // verilog/coms.v(130[12] 305[6])
    defparam i13104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13101_3_lut (.I0(\data_in_frame[3] [5]), .I1(rx_data[5]), .I2(n27898), 
            .I3(GND_net), .O(n28946));   // verilog/coms.v(130[12] 305[6])
    defparam i13101_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13095_3_lut (.I0(\data_in_frame[3] [3]), .I1(rx_data[3]), .I2(n27898), 
            .I3(GND_net), .O(n28940));   // verilog/coms.v(130[12] 305[6])
    defparam i13095_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6228_2_lut (.I0(hall3), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(n21262));   // verilog/TinyFPGA_B.v(168[4] 170[7])
    defparam i6228_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i46864_4_lut (.I0(data_ready), .I1(n6911), .I2(n24_adj_5828), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n63121));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i46864_4_lut.LUT_INIT = 16'hdccc;
    SB_LUT4 i46907_2_lut (.I0(n24_adj_5828), .I1(n6911), .I2(GND_net), 
            .I3(GND_net), .O(n63124));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i46907_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i49_4_lut (.I0(n63124), .I1(n63121), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(n6_adj_5815), .O(n53719));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i49_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1821 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [2]), 
            .O(n55269));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1821.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1822 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [3]), 
            .O(n55268));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1822.LUT_INIT = 16'h2300;
    SB_LUT4 i6232_2_lut (.I0(hall3), .I1(hall1), .I2(GND_net), .I3(GND_net), 
            .O(commutation_state_7__N_27[2]));   // verilog/TinyFPGA_B.v(174[4] 176[7])
    defparam i6232_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1823 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [4]), 
            .O(n55267));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1823.LUT_INIT = 16'h2300;
    SB_LUT4 i39300_3_lut (.I0(n4_adj_5835), .I1(commutation_state_7__N_27[2]), 
            .I2(commutation_state[2]), .I3(GND_net), .O(n56301));   // verilog/TinyFPGA_B.v(151[9] 230[5])
    defparam i39300_3_lut.LUT_INIT = 16'hdcdc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1824 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [5]), 
            .O(n28721));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1824.LUT_INIT = 16'h2300;
    SB_LUT4 i13747_4_lut (.I0(n58594), .I1(r_Bit_Index[0]), .I2(n56281), 
            .I3(n27312), .O(n29592));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i13747_4_lut.LUT_INIT = 16'h32c8;
    SB_LUT4 i13744_4_lut (.I0(n58374), .I1(r_Bit_Index_adj_5924[0]), .I2(n57036), 
            .I3(n27315), .O(n29589));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i13744_4_lut.LUT_INIT = 16'h31c4;
    SB_LUT4 i13729_4_lut (.I0(commutation_state_7__N_27[2]), .I1(commutation_state[1]), 
            .I2(n21262), .I3(n4_adj_5835), .O(n29574));   // verilog/TinyFPGA_B.v(151[9] 230[5])
    defparam i13729_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i11_4_lut (.I0(\data_in_frame[23] [6]), .I1(n38695), .I2(n27939), 
            .I3(rx_data[6]), .O(n54695));   // verilog/coms.v(130[12] 305[6])
    defparam i11_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1825 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [6]), 
            .O(n55241));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1825.LUT_INIT = 16'h2300;
    SB_LUT4 i3_4_lut_adj_1826 (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), 
            .I2(delay_counter[31]), .I3(\ID_READOUT_FSM.state [0]), .O(n58312));
    defparam i3_4_lut_adj_1826.LUT_INIT = 16'h0004;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1827 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[21] [7]), 
            .O(n55266));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1827.LUT_INIT = 16'h2300;
    SB_LUT4 i11_4_lut_adj_1828 (.I0(\data_in_frame[23] [5]), .I1(n38695), 
            .I2(n27939), .I3(rx_data[5]), .O(n54697));   // verilog/coms.v(130[12] 305[6])
    defparam i11_4_lut_adj_1828.LUT_INIT = 16'hca0a;
    SB_LUT4 i13713_3_lut (.I0(\data_in_frame[23] [4]), .I1(rx_data[4]), 
            .I2(n27939), .I3(GND_net), .O(n29558));   // verilog/coms.v(130[12] 305[6])
    defparam i13713_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13710_3_lut (.I0(\data_in_frame[23] [3]), .I1(rx_data[3]), 
            .I2(n27939), .I3(GND_net), .O(n29555));   // verilog/coms.v(130[12] 305[6])
    defparam i13710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13707_3_lut (.I0(\data_in_frame[23] [2]), .I1(rx_data[2]), 
            .I2(n27939), .I3(GND_net), .O(n29552));   // verilog/coms.v(130[12] 305[6])
    defparam i13707_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13704_3_lut (.I0(\data_in_frame[23] [1]), .I1(rx_data[1]), 
            .I2(n27939), .I3(GND_net), .O(n29549));   // verilog/coms.v(130[12] 305[6])
    defparam i13704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1829 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [0]), 
            .O(n55265));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1829.LUT_INIT = 16'h2300;
    SB_LUT4 i13701_3_lut (.I0(\data_in_frame[23] [0]), .I1(rx_data[0]), 
            .I2(n27939), .I3(GND_net), .O(n29546));   // verilog/coms.v(130[12] 305[6])
    defparam i13701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1830 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [1]), 
            .O(n55264));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1830.LUT_INIT = 16'h2300;
    SB_LUT4 i13216_3_lut_3_lut (.I0(\FRAME_MATCHER.rx_data_ready_prev ), .I1(rx_data_ready), 
            .I2(reset), .I3(GND_net), .O(n29061));   // verilog/coms.v(130[12] 305[6])
    defparam i13216_3_lut_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1831 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [2]), 
            .O(n55263));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1831.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1832 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [3]), 
            .O(n55262));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1832.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1833 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [4]), 
            .O(n55261));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1833.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1834 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [5]), 
            .O(n28713));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1834.LUT_INIT = 16'h2300;
    SB_LUT4 i13961_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5899[6]), 
            .I2(n38386), .I3(n25100), .O(n29806));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13961_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1835 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [0]), 
            .O(n55404));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1835.LUT_INIT = 16'h2300;
    SB_LUT4 i13963_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5899[1]), 
            .I2(n10_adj_5812), .I3(n25095), .O(n29808));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13963_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13964_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5899[2]), 
            .I2(n4_adj_5742), .I3(n25100), .O(n29809));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13964_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13965_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5899[3]), 
            .I2(n4_adj_5742), .I3(n25095), .O(n29810));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13965_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13966_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5899[4]), 
            .I2(n4_adj_5743), .I3(n25100), .O(n29811));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13966_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13967_4_lut (.I0(state_7__N_4126[3]), .I1(data_adj_5899[5]), 
            .I2(n4_adj_5743), .I3(n25095), .O(n29812));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13967_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1836 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [1]), 
            .O(n55403));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1836.LUT_INIT = 16'h2300;
    SB_LUT4 i13969_4_lut (.I0(CS_MISO_c), .I1(data_adj_5906[1]), .I2(n5_adj_5746), 
            .I3(n25110), .O(n29814));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13969_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13970_4_lut (.I0(CS_MISO_c), .I1(data_adj_5906[2]), .I2(n5_adj_5771), 
            .I3(n25110), .O(n29815));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13970_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1837 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [6]), 
            .O(n55260));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1837.LUT_INIT = 16'h2300;
    SB_LUT4 i13971_4_lut (.I0(CS_MISO_c), .I1(data_adj_5906[3]), .I2(n38316), 
            .I3(n25110), .O(n29816));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13971_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i13972_4_lut (.I0(CS_MISO_c), .I1(data_adj_5906[4]), .I2(n5_adj_5761), 
            .I3(n25141), .O(n29817));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13972_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13973_4_lut (.I0(CS_MISO_c), .I1(data_adj_5906[5]), .I2(n5_adj_5746), 
            .I3(n25141), .O(n29818));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13973_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1838 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[22] [7]), 
            .O(n28711));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1838.LUT_INIT = 16'h2300;
    SB_LUT4 i13974_4_lut (.I0(CS_MISO_c), .I1(data_adj_5906[6]), .I2(n5_adj_5771), 
            .I3(n25141), .O(n29819));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13974_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1839 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [0]), 
            .O(n55259));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1839.LUT_INIT = 16'h2300;
    SB_LUT4 i13975_4_lut (.I0(CS_MISO_c), .I1(data_adj_5906[7]), .I2(n38316), 
            .I3(n25141), .O(n29820));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13975_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1840 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [2]), 
            .O(n55419));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1840.LUT_INIT = 16'h2300;
    SB_LUT4 i13976_4_lut (.I0(CS_MISO_c), .I1(data_adj_5906[8]), .I2(n5_adj_5761), 
            .I3(n25133), .O(n29821));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13976_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13977_4_lut (.I0(CS_MISO_c), .I1(data_adj_5906[9]), .I2(n5_adj_5746), 
            .I3(n25133), .O(n29822));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13977_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13978_4_lut (.I0(CS_MISO_c), .I1(data_adj_5906[10]), .I2(n5_adj_5771), 
            .I3(n25133), .O(n29823));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13978_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1841 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [3]), 
            .O(n55402));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1841.LUT_INIT = 16'h2300;
    SB_LUT4 i13979_4_lut (.I0(CS_MISO_c), .I1(data_adj_5906[11]), .I2(n38316), 
            .I3(n25133), .O(n29824));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13979_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i13980_4_lut (.I0(CS_MISO_c), .I1(data_adj_5906[12]), .I2(n5_adj_5761), 
            .I3(n25130), .O(n29825));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13980_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1842 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [4]), 
            .O(n55401));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1842.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1843 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [5]), 
            .O(n55400));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1843.LUT_INIT = 16'h2300;
    SB_LUT4 i13981_4_lut (.I0(CS_MISO_c), .I1(data_adj_5906[15]), .I2(n38316), 
            .I3(n25130), .O(n29826));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13981_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1844 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [6]), 
            .O(n55399));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1844.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1845 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[4] [7]), 
            .O(n55398));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1845.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1846 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [0]), 
            .O(n55397));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1846.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1847 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [1]), 
            .O(n55396));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1847.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1848 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [2]), 
            .O(n55395));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1848.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1849 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [3]), 
            .O(n55300));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1849.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1850 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [4]), 
            .O(n55394));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1850.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1851 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [5]), 
            .O(n55393));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1851.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1852 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [1]), 
            .O(n55258));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1852.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1853 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [2]), 
            .O(n55257));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1853.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1854 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [3]), 
            .O(n55256));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1854.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1855 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [4]), 
            .O(n28706));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1855.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1856 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [6]), 
            .O(n55392));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1856.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1857 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [5]), 
            .O(n55255));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1857.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1858 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[5] [7]), 
            .O(n55391));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1858.LUT_INIT = 16'h2300;
    SB_LUT4 i13215_3_lut (.I0(b_prev), .I1(b_new[1]), .I2(debounce_cnt_N_3833), 
            .I3(GND_net), .O(n29060));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13215_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13217_3_lut (.I0(a_prev), .I1(a_new[1]), .I2(debounce_cnt_N_3833), 
            .I3(GND_net), .O(n29062));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13217_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_4_lut (.I0(rx_data_ready), .I1(r_SM_Main[1]), .I2(r_SM_Main[2]), 
            .I3(n27308), .O(n51425));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h0caa;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1859 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [6]), 
            .O(n55254));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1859.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_adj_1860 (.I0(\data_out_frame[18] [6]), .I1(n55884), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5834));
    defparam i1_2_lut_adj_1860.LUT_INIT = 16'h6666;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .clk16MHz(clk16MHz), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(42[10] 46[2])
    SB_LUT4 i4_4_lut_adj_1861 (.I0(n51161), .I1(n25494), .I2(n55766), 
            .I3(n6_adj_5834), .O(n50591));
    defparam i4_4_lut_adj_1861.LUT_INIT = 16'h6996;
    \quadrature_decoder(0)_U0  quad_counter0 (.ENCODER0_B_N_keep(ENCODER0_B_N), 
            .n1795(clk16MHz), .ENCODER0_A_N_keep(ENCODER0_A_N), .n1751(n1751), 
            .GND_net(GND_net), .n1753(n1753), .n1755(n1755), .n1757(n1757), 
            .n1759(n1759), .n1761(n1761), .n1763(n1763), .n1765(n1765), 
            .n1767(n1767), .n1769(n1769), .\encoder0_position[21] (encoder0_position[21]), 
            .\encoder0_position[20] (encoder0_position[20]), .\encoder0_position[19] (encoder0_position[19]), 
            .\encoder0_position[18] (encoder0_position[18]), .\encoder0_position[17] (encoder0_position[17]), 
            .\encoder0_position[16] (encoder0_position[16]), .\encoder0_position[15] (encoder0_position[15]), 
            .\encoder0_position[14] (encoder0_position[14]), .\encoder0_position[13] (encoder0_position[13]), 
            .\encoder0_position[12] (encoder0_position[12]), .\encoder0_position[11] (encoder0_position[11]), 
            .\encoder0_position[10] (encoder0_position[10]), .\encoder0_position[9] (encoder0_position[9]), 
            .\encoder0_position[8] (encoder0_position[8]), .\encoder0_position[7] (encoder0_position[7]), 
            .\encoder0_position[6] (encoder0_position[6]), .\encoder0_position[5] (encoder0_position[5]), 
            .\encoder0_position[4] (encoder0_position[4]), .\encoder0_position[3] (encoder0_position[3]), 
            .\encoder0_position[2] (encoder0_position[2]), .\encoder0_position[1] (encoder0_position[1]), 
            .\encoder0_position[0] (encoder0_position[0]), .VCC_net(VCC_net), 
            .\a_new[1] (a_new[1]), .\b_new[1] (b_new[1]), .b_prev(b_prev), 
            .n29063(n29063), .n1749(n1749), .n29062(n29062), .a_prev(a_prev), 
            .n29060(n29060), .position_31__N_3836(position_31__N_3836), 
            .debounce_cnt_N_3833(debounce_cnt_N_3833)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(313[27] 319[6])
    SB_LUT4 i13219_3_lut (.I0(a_prev_adj_5751), .I1(a_new_adj_5885[1]), 
            .I2(debounce_cnt_N_3833_adj_5753), .I3(GND_net), .O(n29064));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13219_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_4_lut_adj_1862 (.I0(n62), .I1(delay_counter[31]), .I2(data_ready), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n6_adj_5815));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i2_3_lut_4_lut_adj_1862.LUT_INIT = 16'h2022;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1863 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[23] [7]), 
            .O(n28703));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1863.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_adj_1864 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1325), .I3(n38194), .O(n24_adj_5828));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_adj_1864.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1865 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [0]), 
            .O(n55390));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1865.LUT_INIT = 16'h2300;
    SB_LUT4 n66669_bdd_4_lut (.I0(n66669), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(byte_transmit_counter[2]), 
            .O(n66672));
    defparam n66669_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5115_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_372));   // verilog/TinyFPGA_B.v(187[7] 206[15])
    defparam i5115_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1866 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [0]), 
            .O(n55301));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1866.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1867 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [1]), 
            .O(n55389));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1867.LUT_INIT = 16'h2300;
    SB_LUT4 i5113_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_355));   // verilog/TinyFPGA_B.v(187[7] 206[15])
    defparam i5113_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1868 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [2]), 
            .O(n55388));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1868.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(current[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5727));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1869 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [3]), 
            .O(n55387));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1869.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_11_i7_2_lut (.I0(current[3]), .I1(duty[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5738));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam LessThan_11_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(current[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5736));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(current[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5730));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(current[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5729));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1870 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [4]), 
            .O(n55386));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1870.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(current[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5728));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(current[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5734));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(current[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5733));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(current[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5732));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1871 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [1]), 
            .O(n55253));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1871.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_14_i13_2_lut (.I0(current[6]), .I1(current_limit[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5719));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam LessThan_14_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i15_2_lut (.I0(current[7]), .I1(current_limit[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5718));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam LessThan_14_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1872 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [2]), 
            .O(n55252));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1872.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_14_i19_2_lut (.I0(current[9]), .I1(current_limit[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5715));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam LessThan_14_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i17_2_lut (.I0(current[8]), .I1(current_limit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5716));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam LessThan_14_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i7_2_lut (.I0(current[3]), .I1(current_limit[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5723));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam LessThan_14_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i9_2_lut (.I0(current[4]), .I1(current_limit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5721));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam LessThan_14_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1873 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [3]), 
            .O(n55251));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1873.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_14_i11_2_lut (.I0(current[5]), .I1(current_limit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5720));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam LessThan_14_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_14_i5_2_lut (.I0(current[2]), .I1(current_limit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5725));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam LessThan_14_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1874 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [4]), 
            .O(n55250));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1874.LUT_INIT = 16'h2300;
    SB_LUT4 i46946_4_lut (.I0(n11_adj_5720), .I1(n9_adj_5721), .I2(n7_adj_5723), 
            .I3(n5_adj_5725), .O(n64008));
    defparam i46946_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1875 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [5]), 
            .O(n55249));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1875.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1876 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [6]), 
            .O(n28696));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1876.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_adj_1877 (.I0(n50591), .I1(\data_out_frame[16] [5]), 
            .I2(\data_out_frame[18] [6]), .I3(\data_out_frame[18] [5]), 
            .O(n51296));
    defparam i1_2_lut_4_lut_adj_1877.LUT_INIT = 16'h6996;
    SB_LUT4 LessThan_14_i16_3_lut (.I0(n8_adj_5722), .I1(current_limit[9]), 
            .I2(n19_adj_5715), .I3(GND_net), .O(n16_adj_5717));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam LessThan_14_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_14_i4_4_lut (.I0(current_limit[0]), .I1(current_limit[1]), 
            .I2(current[1]), .I3(current[0]), .O(n4_adj_5726));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam LessThan_14_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i48609_3_lut (.I0(n4_adj_5726), .I1(current_limit[5]), .I2(n11_adj_5720), 
            .I3(GND_net), .O(n65671));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam i48609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48610_3_lut (.I0(n65671), .I1(current_limit[6]), .I2(n13_adj_5719), 
            .I3(GND_net), .O(n65672));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam i48610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46926_4_lut (.I0(n17_adj_5716), .I1(n15_adj_5718), .I2(n13_adj_5719), 
            .I3(n64008), .O(n63988));
    defparam i46926_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1878 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[24] [7]), 
            .O(n55299));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1878.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1879 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [0]), 
            .O(n55248));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1879.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1880 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [1]), 
            .O(n55247));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1880.LUT_INIT = 16'h2300;
    SB_LUT4 i48855_4_lut (.I0(n16_adj_5717), .I1(n6_adj_5724), .I2(n19_adj_5715), 
            .I3(n63986), .O(n65917));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam i48855_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47236_3_lut (.I0(n65672), .I1(current_limit[7]), .I2(n15_adj_5718), 
            .I3(GND_net), .O(n64298));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam i47236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49138_4_lut (.I0(n64298), .I1(n65917), .I2(n19_adj_5715), 
            .I3(n63988), .O(n66200));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam i49138_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49139_3_lut (.I0(n66200), .I1(current_limit[10]), .I2(current[10]), 
            .I3(GND_net), .O(n66201));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam i49139_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1881 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [2]), 
            .O(n55246));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1881.LUT_INIT = 16'h2300;
    SB_LUT4 i49052_3_lut (.I0(n66201), .I1(current_limit[11]), .I2(current[11]), 
            .I3(GND_net), .O(n24_adj_5714));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam i49052_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1882 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [3]), 
            .O(n55245));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1882.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1883 (.I0(current_limit[13]), .I1(n24_adj_5714), 
            .I2(current_limit[14]), .I3(current_limit[12]), .O(n58026));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam i1_4_lut_adj_1883.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1884 (.I0(current_limit[13]), .I1(n24_adj_5714), 
            .I2(current_limit[14]), .I3(current_limit[12]), .O(n58029));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam i1_4_lut_adj_1884.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_1885 (.I0(current[15]), .I1(current_limit[15]), 
            .I2(n58029), .I3(n58026), .O(n260));   // verilog/TinyFPGA_B.v(126[9:30])
    defparam i1_4_lut_adj_1885.LUT_INIT = 16'hb3a2;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1886 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [4]), 
            .O(n55244));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1886.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i25_2_lut (.I0(duty[12]), .I1(n298), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam LessThan_17_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i23_2_lut (.I0(duty[11]), .I1(n299), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam LessThan_17_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i21_2_lut (.I0(duty[10]), .I1(n300), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam LessThan_17_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(duty[9]), .I1(n301), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5693));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i7_2_lut (.I0(duty[3]), .I1(n307), .I2(GND_net), 
            .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam LessThan_17_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1887 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [5]), 
            .O(n28689));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1887.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i9_2_lut (.I0(duty[4]), .I1(n306), .I2(GND_net), 
            .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(duty[5]), .I1(n305), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_Bit_Index[0]), .I1(r_SM_Main[1]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main[2]), .O(n58932));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(duty[6]), .I1(n304), .I2(GND_net), 
            .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(duty[7]), .I1(n303), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1888 (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[1]), .I3(r_Bit_Index[0]), .O(n58896));
    defparam i1_3_lut_4_lut_adj_1888.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1889 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [5]), 
            .O(n55385));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1889.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1890 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [6]), 
            .O(n28688));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1890.LUT_INIT = 16'h2300;
    SB_LUT4 i13092_3_lut_4_lut (.I0(n1800), .I1(b_prev_adj_5752), .I2(a_new_adj_5885[1]), 
            .I3(position_31__N_3836_adj_5754), .O(n28937));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    defparam i13092_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(duty[8]), .I1(n302), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i5_2_lut (.I0(duty[2]), .I1(n308), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam LessThan_17_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46337_4_lut (.I0(n11), .I1(n9), .I2(n7), .I3(n5), .O(n63399));
    defparam i46337_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46330_4_lut (.I0(n17), .I1(n15), .I2(n13), .I3(n63399), 
            .O(n63392));
    defparam i46330_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1891 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[25] [7]), 
            .O(n55243));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1891.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_17_i10_3_lut (.I0(n305), .I1(n304), .I2(n13), .I3(GND_net), 
            .O(n10));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam LessThan_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i4_3_lut (.I0(n62960), .I1(n309), .I2(duty[1]), 
            .I3(GND_net), .O(n4));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam LessThan_17_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_17_i12_3_lut (.I0(n10), .I1(n303), .I2(n15), .I3(GND_net), 
            .O(n12));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam LessThan_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1892 (.I0(duty[15]), .I1(duty[20]), .I2(n294), 
            .I3(GND_net), .O(n12_adj_5820));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam i2_3_lut_adj_1892.LUT_INIT = 16'h7e7e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1893 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [6]), 
            .O(n55384));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1893.LUT_INIT = 16'h2300;
    SB_LUT4 mux_1677_i22_3_lut (.I0(duty[23]), .I1(duty[21]), .I2(n260), 
            .I3(GND_net), .O(n11588));   // verilog/TinyFPGA_B.v(125[13] 136[7])
    defparam mux_1677_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i6_4_lut_adj_1894 (.I0(duty[13]), .I1(n12_adj_5820), .I2(duty[21]), 
            .I3(n294), .O(n16_adj_5818));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam i6_4_lut_adj_1894.LUT_INIT = 16'hdffe;
    SB_LUT4 i4_3_lut (.I0(duty[19]), .I1(duty[16]), .I2(n294), .I3(GND_net), 
            .O(n14_adj_5819));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam i4_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 LessThan_17_i8_3_lut (.I0(n306), .I1(n302), .I2(n17), .I3(GND_net), 
            .O(n8_adj_5713));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam LessThan_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i6_3_lut (.I0(n308), .I1(n307), .I2(n7), .I3(GND_net), 
            .O(n6));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam LessThan_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n8_adj_5713), .I1(n301), .I2(n19_adj_5693), 
            .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48947_4_lut (.I0(n16), .I1(n6), .I2(n19_adj_5693), .I3(n63388), 
            .O(n66009));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam i48947_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1895 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[6] [7]), 
            .O(n55383));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1895.LUT_INIT = 16'h2300;
    SB_LUT4 i48948_3_lut (.I0(n66009), .I1(n300), .I2(n21), .I3(GND_net), 
            .O(n66010));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam i48948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48694_3_lut (.I0(n66010), .I1(n299), .I2(n23), .I3(GND_net), 
            .O(n65756));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam i48694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48422_4_lut (.I0(n23), .I1(n21), .I2(n19_adj_5693), .I3(n63392), 
            .O(n65484));
    defparam i48422_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48387_4_lut (.I0(n12), .I1(n4), .I2(n15), .I3(n63397), 
            .O(n65449));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam i48387_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48036_3_lut (.I0(n65756), .I1(n298), .I2(n25), .I3(GND_net), 
            .O(n65098));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam i48036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1896 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [0]), 
            .O(n55382));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1896.LUT_INIT = 16'h2300;
    SB_LUT4 i8_4_lut_adj_1897 (.I0(duty[14]), .I1(n16_adj_5818), .I2(duty[18]), 
            .I3(n294), .O(n18_adj_5816));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam i8_4_lut_adj_1897.LUT_INIT = 16'hdffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1898 (.I0(n2882), .I1(n56366), .I2(n38266), 
            .I3(\FRAME_MATCHER.i [0]), .O(n27939));
    defparam i1_2_lut_3_lut_4_lut_adj_1898.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1899 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [1]), 
            .O(n55381));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1899.LUT_INIT = 16'h2300;
    SB_LUT4 i7_4_lut_adj_1900 (.I0(duty[22]), .I1(n14_adj_5819), .I2(duty[17]), 
            .I3(n294), .O(n17_adj_5817));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam i7_4_lut_adj_1900.LUT_INIT = 16'hdffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1901 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [2]), 
            .O(n55380));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1901.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1902 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [3]), 
            .O(n55379));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1902.LUT_INIT = 16'h2300;
    SB_LUT4 i48460_4_lut (.I0(n65098), .I1(n65449), .I2(n25), .I3(n65484), 
            .O(n65522));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam i48460_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48461_4_lut (.I0(n65522), .I1(n294), .I2(n17_adj_5817), .I3(n18_adj_5816), 
            .O(n65523));   // verilog/TinyFPGA_B.v(129[11:24])
    defparam i48461_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i39506_4_lut (.I0(n260), .I1(duty[23]), .I2(n294), .I3(n65523), 
            .O(n9939));
    defparam i39506_4_lut.LUT_INIT = 16'h1151;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1903 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [4]), 
            .O(n55378));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1903.LUT_INIT = 16'h2300;
    SB_LUT4 i47498_3_lut (.I0(n15_adj_5732), .I1(n13_adj_5733), .I2(n11_adj_5734), 
            .I3(GND_net), .O(n64560));
    defparam i47498_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1904 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [5]), 
            .O(n55377));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1904.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1905 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [6]), 
            .O(n55302));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1905.LUT_INIT = 16'h2300;
    SB_LUT4 i47377_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n64560), .O(n64439));
    defparam i47377_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i46476_4_lut (.I0(n21_adj_5728), .I1(n19_adj_5729), .I2(n17_adj_5730), 
            .I3(n9_adj_5736), .O(n63538));
    defparam i46476_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47520_4_lut (.I0(n9_adj_5736), .I1(n7_adj_5738), .I2(current[2]), 
            .I3(duty[2]), .O(n64582));
    defparam i47520_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1906 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [2]), 
            .O(n55418));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1906.LUT_INIT = 16'h2300;
    SB_LUT4 i48105_4_lut (.I0(n15_adj_5732), .I1(n13_adj_5733), .I2(n11_adj_5734), 
            .I3(n64582), .O(n65167));
    defparam i48105_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48097_4_lut (.I0(n21_adj_5728), .I1(n19_adj_5729), .I2(n17_adj_5730), 
            .I3(n65167), .O(n65159));
    defparam i48097_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1907 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [3]), 
            .O(n55417));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1907.LUT_INIT = 16'h2300;
    SB_LUT4 i48789_4_lut (.I0(current[15]), .I1(n23_adj_5727), .I2(duty[12]), 
            .I3(n65159), .O(n65851));
    defparam i48789_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i47446_4_lut (.I0(current[15]), .I1(duty[13]), .I2(duty[14]), 
            .I3(n65851), .O(n64508));
    defparam i47446_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(current[0]), .I1(duty[1]), .I2(current[1]), 
            .I3(duty[0]), .O(n4_adj_5740));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i48163_3_lut (.I0(n4_adj_5740), .I1(duty[13]), .I2(current[15]), 
            .I3(GND_net), .O(n65225));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam i48163_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47363_4_lut (.I0(current[15]), .I1(duty[16]), .I2(duty[17]), 
            .I3(n15_adj_5732), .O(n64425));
    defparam i47363_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1908 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[0] [4]), 
            .O(n55416));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1908.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1909 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [0]), 
            .O(n55415));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1909.LUT_INIT = 16'h2300;
    SB_LUT4 LessThan_11_i30_4_lut (.I0(duty[7]), .I1(duty[17]), .I2(current[15]), 
            .I3(duty[16]), .O(n30));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam LessThan_11_i30_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i46428_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n64439), .O(n63490));
    defparam i46428_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 i13251_3_lut (.I0(current[11]), .I1(data_adj_5906[11]), .I2(n27290), 
            .I3(GND_net), .O(n29096));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i35_rep_309_2_lut (.I0(current[15]), .I1(duty[17]), 
            .I2(GND_net), .I3(GND_net), .O(n67455));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam LessThan_11_i35_rep_309_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49035_3_lut (.I0(n30), .I1(n10_adj_5735), .I2(n64425), .I3(GND_net), 
            .O(n66097));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam i49035_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1910 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [1]), 
            .O(n55414));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1910.LUT_INIT = 16'h2300;
    SB_LUT4 i47246_4_lut (.I0(n65225), .I1(duty[15]), .I2(current[15]), 
            .I3(duty[14]), .O(n64308));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam i47246_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i48159_3_lut (.I0(n6_adj_5739), .I1(duty[10]), .I2(n21_adj_5728), 
            .I3(GND_net), .O(n65221));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam i48159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48160_3_lut (.I0(n65221), .I1(duty[11]), .I2(n23_adj_5727), 
            .I3(GND_net), .O(n65222));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam i48160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13252_3_lut (.I0(current[10]), .I1(data_adj_5906[10]), .I2(n27290), 
            .I3(GND_net), .O(n29097));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48089_4_lut (.I0(current[15]), .I1(n23_adj_5727), .I2(duty[12]), 
            .I3(n63538), .O(n65151));
    defparam i48089_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n8_adj_5737), .I1(duty[9]), .I2(n19_adj_5729), 
            .I3(GND_net), .O(n16_adj_5731));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1911 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [3]), 
            .O(n55413));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1911.LUT_INIT = 16'h2300;
    SB_LUT4 i47248_3_lut (.I0(n65222), .I1(duty[12]), .I2(current[15]), 
            .I3(GND_net), .O(n64310));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam i47248_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48464_4_lut (.I0(current[15]), .I1(duty[15]), .I2(duty[16]), 
            .I3(n64508), .O(n65526));
    defparam i48464_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i49169_4_lut (.I0(n64308), .I1(n66097), .I2(n67455), .I3(n63490), 
            .O(n66231));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam i49169_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1912 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [5]), 
            .O(n55412));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1912.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1913 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [6]), 
            .O(n55411));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1913.LUT_INIT = 16'h2300;
    SB_LUT4 i48395_3_lut (.I0(n64310), .I1(n16_adj_5731), .I2(n65151), 
            .I3(GND_net), .O(n65457));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam i48395_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i49191_4_lut (.I0(n65457), .I1(n66231), .I2(n67455), .I3(n65526), 
            .O(n66253));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam i49191_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1914 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[1] [7]), 
            .O(n55410));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1914.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1915 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[7] [7]), 
            .O(n55376));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1915.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1916 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [2]), 
            .O(n55303));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1916.LUT_INIT = 16'h2300;
    SB_LUT4 i13253_3_lut (.I0(current[9]), .I1(data_adj_5906[9]), .I2(n27290), 
            .I3(GND_net), .O(n29098));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49182_4_lut (.I0(n66253), .I1(duty[19]), .I2(current[15]), 
            .I3(duty[18]), .O(n66244));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam i49182_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i2_2_lut_adj_1917 (.I0(current[15]), .I1(duty[22]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5809));
    defparam i2_2_lut_adj_1917.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1918 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [3]), 
            .O(n55375));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1918.LUT_INIT = 16'h2300;
    SB_LUT4 i48716_4_lut (.I0(n66244), .I1(duty[21]), .I2(current[15]), 
            .I3(duty[20]), .O(n65778));   // verilog/TinyFPGA_B.v(118[10:22])
    defparam i48716_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i7_4_lut_adj_1919 (.I0(n65778), .I1(duty[23]), .I2(n6_adj_5809), 
            .I3(n260), .O(n9941));
    defparam i7_4_lut_adj_1919.LUT_INIT = 16'h3332;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1920 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [4]), 
            .O(n55374));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1920.LUT_INIT = 16'h2300;
    SB_LUT4 i13254_3_lut (.I0(current[8]), .I1(data_adj_5906[8]), .I2(n27290), 
            .I3(GND_net), .O(n29099));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1921 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [5]), 
            .O(n55373));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1921.LUT_INIT = 16'h2300;
    SB_LUT4 i13255_3_lut (.I0(current[7]), .I1(data_adj_5906[7]), .I2(n27290), 
            .I3(GND_net), .O(n29100));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1922 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [6]), 
            .O(n55372));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1922.LUT_INIT = 16'h2300;
    SB_LUT4 i13256_3_lut (.I0(current[6]), .I1(data_adj_5906[6]), .I2(n27290), 
            .I3(GND_net), .O(n29101));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1923 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[8] [7]), 
            .O(n55371));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1923.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1924 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [0]), 
            .O(n55370));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1924.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1925 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [1]), 
            .O(n55369));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1925.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1926 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [2]), 
            .O(n55368));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1926.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1927 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [3]), 
            .O(n55367));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1927.LUT_INIT = 16'h2300;
    SB_LUT4 i5117_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_377));
    defparam i5117_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 i5119_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_386));
    defparam i5119_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1928 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [4]), 
            .O(n55366));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1928.LUT_INIT = 16'h2300;
    SB_LUT4 i13257_3_lut (.I0(current[5]), .I1(data_adj_5906[5]), .I2(n27290), 
            .I3(GND_net), .O(n29102));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1929 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [5]), 
            .O(n55365));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1929.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1930 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [6]), 
            .O(n55364));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1930.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1931 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[9] [7]), 
            .O(n55363));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1931.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1932 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [0]), 
            .O(n55362));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1932.LUT_INIT = 16'h2300;
    SB_LUT4 i13258_3_lut (.I0(current[4]), .I1(data_adj_5906[4]), .I2(n27290), 
            .I3(GND_net), .O(n29103));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1933 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [1]), 
            .O(n55361));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1933.LUT_INIT = 16'h2300;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49582 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [7]), .I2(\data_out_frame[23] [7]), 
            .I3(byte_transmit_counter[2]), .O(n66651));
    defparam byte_transmit_counter_0__bdd_4_lut_49582.LUT_INIT = 16'he4aa;
    SB_LUT4 i13259_3_lut (.I0(current[3]), .I1(data_adj_5906[3]), .I2(n27290), 
            .I3(GND_net), .O(n29104));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_245_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15_adj_5712), .I3(n15_adj_5770), .O(motor_state_23__N_91[9]));   // verilog/TinyFPGA_B.v(294[5] 296[10])
    defparam mux_245_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_243_i10_3_lut (.I0(encoder0_position_scaled[9]), .I1(motor_state_23__N_91[9]), 
            .I2(n15_adj_5748), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(293[5] 296[10])
    defparam mux_243_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1934 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [2]), 
            .O(n55360));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1934.LUT_INIT = 16'h2300;
    SB_LUT4 i13260_3_lut (.I0(current[2]), .I1(data_adj_5906[2]), .I2(n27290), 
            .I3(GND_net), .O(n29105));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1935 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [3]), 
            .O(n55359));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1935.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1936 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [4]), 
            .O(n55358));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1936.LUT_INIT = 16'h2300;
    SB_LUT4 i13261_3_lut (.I0(current[1]), .I1(data_adj_5906[1]), .I2(n27290), 
            .I3(GND_net), .O(n29106));   // verilog/tli4970.v(35[10] 68[6])
    defparam i13261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1937 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [5]), 
            .O(n55357));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1937.LUT_INIT = 16'h2300;
    SB_LUT4 i13262_3_lut (.I0(baudrate[31]), .I1(data_adj_5899[7]), .I2(n57999), 
            .I3(GND_net), .O(n29107));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13262_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1938 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [6]), 
            .O(n55356));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1938.LUT_INIT = 16'h2300;
    SB_LUT4 n66651_bdd_4_lut (.I0(n66651), .I1(\data_out_frame[19] [7]), 
            .I2(\data_out_frame[18] [7]), .I3(byte_transmit_counter[2]), 
            .O(n66654));
    defparam n66651_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1939 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[10] [7]), 
            .O(n55355));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1939.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1940 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [0]), 
            .O(n55354));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1940.LUT_INIT = 16'h2300;
    SB_LUT4 i13263_3_lut (.I0(baudrate[30]), .I1(data_adj_5899[6]), .I2(n57999), 
            .I3(GND_net), .O(n29108));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13263_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1941 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [1]), 
            .O(n55353));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1941.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1942 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [2]), 
            .O(n55352));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1942.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1943 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [3]), 
            .O(n55351));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1943.LUT_INIT = 16'h2300;
    SB_LUT4 i13264_3_lut (.I0(baudrate[29]), .I1(data_adj_5899[5]), .I2(n57999), 
            .I3(GND_net), .O(n29109));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13264_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1944 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [4]), 
            .O(n55350));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1944.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1945 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [5]), 
            .O(n55349));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1945.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1946 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [6]), 
            .O(n55348));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1946.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1947 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[11] [7]), 
            .O(n55347));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1947.LUT_INIT = 16'h2300;
    SB_LUT4 i13265_3_lut (.I0(baudrate[28]), .I1(data_adj_5899[4]), .I2(n57999), 
            .I3(GND_net), .O(n29110));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13265_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1948 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [0]), 
            .O(n55346));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1948.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1949 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [1]), 
            .O(n55345));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1949.LUT_INIT = 16'h2300;
    SB_LUT4 i13266_3_lut (.I0(baudrate[27]), .I1(data_adj_5899[3]), .I2(n57999), 
            .I3(GND_net), .O(n29111));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13266_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1950 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [2]), 
            .O(n55344));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1950.LUT_INIT = 16'h2300;
    SB_LUT4 i13267_3_lut (.I0(baudrate[26]), .I1(data_adj_5899[2]), .I2(n57999), 
            .I3(GND_net), .O(n29112));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13267_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1951 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [3]), 
            .O(n55343));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1951.LUT_INIT = 16'h2300;
    SB_LUT4 i49479_4_lut_4_lut_4_lut (.I0(hall3), .I1(hall1), .I2(commutation_state_7__N_27[2]), 
            .I3(hall2), .O(n7_adj_5846));
    defparam i49479_4_lut_4_lut_4_lut.LUT_INIT = 16'h77fc;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1952 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [4]), 
            .O(n55342));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1952.LUT_INIT = 16'h2300;
    SB_LUT4 i13268_3_lut (.I0(baudrate[25]), .I1(data_adj_5899[1]), .I2(n57999), 
            .I3(GND_net), .O(n29113));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13268_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1953 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [5]), 
            .O(n55341));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1953.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1954 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [6]), 
            .O(n55340));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1954.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1955 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[12] [7]), 
            .O(n55339));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1955.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1956 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [0]), 
            .O(n55338));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1956.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1957 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [1]), 
            .O(n55337));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1957.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1958 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [2]), 
            .O(n55336));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1958.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1959 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [3]), 
            .O(n55335));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1959.LUT_INIT = 16'h2300;
    SB_LUT4 i13269_3_lut (.I0(baudrate[24]), .I1(data_adj_5899[0]), .I2(n57999), 
            .I3(GND_net), .O(n29114));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13269_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1960 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [4]), 
            .O(n55334));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1960.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1961 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [5]), 
            .O(n55333));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1961.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1962 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [6]), 
            .O(n55332));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1962.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1963 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[13] [7]), 
            .O(n55331));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1963.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1964 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [0]), 
            .O(n55330));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1964.LUT_INIT = 16'h2300;
    SB_LUT4 i13586_3_lut (.I0(\data_in_frame[18] [4]), .I1(rx_data[4]), 
            .I2(n27929), .I3(GND_net), .O(n29431));   // verilog/coms.v(130[12] 305[6])
    defparam i13586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1965 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [1]), 
            .O(n55329));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1965.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1966 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [2]), 
            .O(n55328));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1966.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1967 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [3]), 
            .O(n55327));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1967.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1968 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [4]), 
            .O(n55326));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1968.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1969 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [5]), 
            .O(n55325));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1969.LUT_INIT = 16'h2300;
    SB_LUT4 i21362_4_lut (.I0(n78), .I1(n67), .I2(rx_data[6]), .I3(\data_in_frame[16] [6]), 
            .O(n37128));   // verilog/coms.v(94[13:20])
    defparam i21362_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i2_2_lut_adj_1970 (.I0(dti_counter[1]), .I1(dti_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5832));   // verilog/TinyFPGA_B.v(179[9:23])
    defparam i2_2_lut_adj_1970.LUT_INIT = 16'heeee;
    SB_LUT4 i21363_3_lut (.I0(n37128), .I1(\data_in_frame[16] [6]), .I2(reset), 
            .I3(GND_net), .O(n29389));   // verilog/TinyFPGA_B.v(55[5:10])
    defparam i21363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1971 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [6]), 
            .O(n55305));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1971.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1972 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[14] [7]), 
            .O(n55324));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1972.LUT_INIT = 16'h2300;
    SB_LUT4 i49240_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n38194), .I3(GND_net), .O(n27321));
    defparam i49240_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 i46358_2_lut_3_lut (.I0(n62), .I1(delay_counter[31]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n63020));
    defparam i46358_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_adj_1973 (.I0(\FRAME_MATCHER.i [5]), .I1(n8_adj_5711), 
            .I2(GND_net), .I3(GND_net), .O(n76));
    defparam i1_2_lut_adj_1973.LUT_INIT = 16'heeee;
    SB_LUT4 i22539_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n38194), .I3(GND_net), .O(n38279));
    defparam i22539_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i6_4_lut_adj_1974 (.I0(dti_counter[7]), .I1(dti_counter[4]), 
            .I2(dti_counter[5]), .I3(dti_counter[6]), .O(n14_adj_5831));   // verilog/TinyFPGA_B.v(179[9:23])
    defparam i6_4_lut_adj_1974.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1975 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [0]), 
            .O(n55323));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1975.LUT_INIT = 16'h2300;
    SB_LUT4 i3_4_lut_adj_1976 (.I0(n76), .I1(\FRAME_MATCHER.i [3]), .I2(\FRAME_MATCHER.i [4]), 
            .I3(n56368), .O(n78));
    defparam i3_4_lut_adj_1976.LUT_INIT = 16'hefff;
    SB_LUT4 i21347_4_lut (.I0(n78), .I1(n67), .I2(rx_data[7]), .I3(\data_in_frame[16] [7]), 
            .O(n37113));   // verilog/coms.v(94[13:20])
    defparam i21347_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i21348_3_lut (.I0(n37113), .I1(\data_in_frame[16] [7]), .I2(reset), 
            .I3(GND_net), .O(n29392));   // verilog/TinyFPGA_B.v(55[5:10])
    defparam i21348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1977 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [1]), 
            .O(n55322));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1977.LUT_INIT = 16'h2300;
    SB_LUT4 i13164_3_lut (.I0(\data_in_frame[6] [2]), .I1(rx_data[2]), .I2(n27904), 
            .I3(GND_net), .O(n29009));   // verilog/coms.v(130[12] 305[6])
    defparam i13164_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1978 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [2]), 
            .O(n55321));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1978.LUT_INIT = 16'h2300;
    SB_LUT4 i7_4_lut_adj_1979 (.I0(dti_counter[0]), .I1(n14_adj_5831), .I2(n10_adj_5832), 
            .I3(dti_counter[3]), .O(n22471));   // verilog/TinyFPGA_B.v(179[9:23])
    defparam i7_4_lut_adj_1979.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1980 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [3]), 
            .O(n55320));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1980.LUT_INIT = 16'h2300;
    SB_LUT4 i1_4_lut_adj_1981 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5833));   // verilog/TinyFPGA_B.v(154[7:48])
    defparam i1_4_lut_adj_1981.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1982 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [4]), 
            .O(n55319));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1982.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1983 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [5]), 
            .O(n55318));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1983.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1984 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [6]), 
            .O(n55317));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1984.LUT_INIT = 16'h2300;
    SB_LUT4 i2_3_lut_adj_1985 (.I0(commutation_state[0]), .I1(n4_adj_5833), 
            .I2(commutation_state_prev[0]), .I3(GND_net), .O(n15_adj_5741));   // verilog/TinyFPGA_B.v(154[7:48])
    defparam i2_3_lut_adj_1985.LUT_INIT = 16'hdede;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1986 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[15] [7]), 
            .O(n55304));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1986.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1987 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [0]), 
            .O(n55316));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1987.LUT_INIT = 16'h2300;
    SB_LUT4 i13549_3_lut (.I0(\data_in_frame[17] [0]), .I1(rx_data[0]), 
            .I2(n27926), .I3(GND_net), .O(n29394));   // verilog/coms.v(130[12] 305[6])
    defparam i13549_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1988 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [1]), 
            .O(n55315));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1988.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1989 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [2]), 
            .O(n55314));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1989.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1990 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [3]), 
            .O(n55313));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1990.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1991 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [4]), 
            .O(n55312));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1991.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1992 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [5]), 
            .O(n55311));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1992.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1993 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [6]), 
            .O(n55310));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1993.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1994 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[16] [7]), 
            .O(n55309));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1994.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1995 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [0]), 
            .O(n55308));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1995.LUT_INIT = 16'h2300;
    SB_LUT4 i13552_3_lut (.I0(\data_in_frame[17] [1]), .I1(rx_data[1]), 
            .I2(n27926), .I3(GND_net), .O(n29397));   // verilog/coms.v(130[12] 305[6])
    defparam i13552_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1996 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [1]), 
            .O(n55307));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1996.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1997 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [2]), 
            .O(n55306));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1997.LUT_INIT = 16'h2300;
    SB_LUT4 i13555_3_lut (.I0(\data_in_frame[17] [2]), .I1(rx_data[2]), 
            .I2(n27926), .I3(GND_net), .O(n29400));   // verilog/coms.v(130[12] 305[6])
    defparam i13555_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(read_N_409), .I3(n2829), .O(n25_adj_5827));   // verilog/TinyFPGA_B.v(385[7:11])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h5450;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1998 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [3]), 
            .O(n55298));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1998.LUT_INIT = 16'h2300;
    SB_LUT4 i13558_3_lut (.I0(\data_in_frame[17] [3]), .I1(rx_data[3]), 
            .I2(n27926), .I3(GND_net), .O(n29403));   // verilog/coms.v(130[12] 305[6])
    defparam i13558_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_1999 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [4]), 
            .O(n55297));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_1999.LUT_INIT = 16'h2300;
    SB_LUT4 i13561_3_lut (.I0(\data_in_frame[17] [4]), .I1(rx_data[4]), 
            .I2(n27926), .I3(GND_net), .O(n29406));   // verilog/coms.v(130[12] 305[6])
    defparam i13561_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13564_3_lut (.I0(\data_in_frame[17] [5]), .I1(rx_data[5]), 
            .I2(n27926), .I3(GND_net), .O(n29409));   // verilog/coms.v(130[12] 305[6])
    defparam i13564_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2000 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [5]), 
            .O(n55296));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2000.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_3_lut_adj_2001 (.I0(hall1), .I1(hall2), .I2(n21262), 
            .I3(GND_net), .O(n4_adj_5835));   // verilog/TinyFPGA_B.v(159[7:22])
    defparam i1_2_lut_3_lut_adj_2001.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2002 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [6]), 
            .O(n55295));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2002.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2003 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[17] [7]), 
            .O(n55294));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2003.LUT_INIT = 16'h2300;
    SB_LUT4 i1_2_lut_4_lut_4_lut_adj_2004 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(reset), .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(\data_out_frame[18] [0]), 
            .O(n55293));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_2_lut_4_lut_4_lut_adj_2004.LUT_INIT = 16'h2300;
    SB_LUT4 i13570_3_lut (.I0(\data_in_frame[17] [7]), .I1(rx_data[7]), 
            .I2(n27926), .I3(GND_net), .O(n29415));   // verilog/coms.v(130[12] 305[6])
    defparam i13570_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[18] [6]), 
            .I2(n10_adj_5837), .I3(\data_out_frame[18] [4]), .O(n24633));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_2005 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[18] [6]), 
            .I2(\data_out_frame[18] [5]), .I3(GND_net), .O(n56109));
    defparam i1_2_lut_3_lut_adj_2005.LUT_INIT = 16'h9696;
    SB_LUT4 i13573_3_lut (.I0(\data_in_frame[18] [0]), .I1(rx_data[0]), 
            .I2(n27929), .I3(GND_net), .O(n29418));   // verilog/coms.v(130[12] 305[6])
    defparam i13573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13278_3_lut (.I0(baudrate[15]), .I1(data_adj_5899[7]), .I2(n55526), 
            .I3(GND_net), .O(n29123));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13278_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i49410_2_lut (.I0(n22471), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_404));
    defparam i49410_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i13279_3_lut (.I0(baudrate[14]), .I1(data_adj_5899[6]), .I2(n55526), 
            .I3(GND_net), .O(n29124));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13279_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13280_3_lut (.I0(baudrate[13]), .I1(data_adj_5899[5]), .I2(n55526), 
            .I3(GND_net), .O(n29125));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13280_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13281_3_lut (.I0(baudrate[12]), .I1(data_adj_5899[4]), .I2(n55526), 
            .I3(GND_net), .O(n29126));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13281_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49543 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [6]), .I2(\data_out_frame[23] [6]), 
            .I3(byte_transmit_counter[1]), .O(n66615));
    defparam byte_transmit_counter_0__bdd_4_lut_49543.LUT_INIT = 16'he4aa;
    SB_LUT4 i13576_3_lut (.I0(\data_in_frame[18] [1]), .I1(rx_data[1]), 
            .I2(n27929), .I3(GND_net), .O(n29421));   // verilog/coms.v(130[12] 305[6])
    defparam i13576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n66615_bdd_4_lut (.I0(n66615), .I1(\data_out_frame[21] [6]), 
            .I2(\data_out_frame[20] [6]), .I3(byte_transmit_counter[1]), 
            .O(n66618));
    defparam n66615_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13579_3_lut (.I0(\data_in_frame[18] [2]), .I1(rx_data[2]), 
            .I2(n27929), .I3(GND_net), .O(n29424));   // verilog/coms.v(130[12] 305[6])
    defparam i13579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13589_3_lut (.I0(\data_in_frame[18] [5]), .I1(rx_data[5]), 
            .I2(n27929), .I3(GND_net), .O(n29434));   // verilog/coms.v(130[12] 305[6])
    defparam i13589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13282_3_lut (.I0(baudrate[11]), .I1(data_adj_5899[3]), .I2(n55526), 
            .I3(GND_net), .O(n29127));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13282_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut_adj_2006 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [7]), 
            .I2(n55587), .I3(n6_adj_5825), .O(Kp_23__N_748));   // verilog/coms.v(99[12:25])
    defparam i4_4_lut_adj_2006.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_4_lut_adj_2007 (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(reset), .I3(n38194), .O(n53805));   // verilog/TinyFPGA_B.v(367[10] 397[6])
    defparam i1_4_lut_4_lut_adj_2007.LUT_INIT = 16'hb1f1;
    SB_LUT4 LessThan_1178_i6_3_lut_3_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(GND_net), .O(n6_adj_5806));   // verilog/uart_rx.v(119[17:57])
    defparam LessThan_1178_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i46364_3_lut_4_lut (.I0(r_Clock_Count[3]), .I1(o_Rx_DV_N_3488[3]), 
            .I2(o_Rx_DV_N_3488[2]), .I3(r_Clock_Count[2]), .O(n63426));   // verilog/uart_rx.v(119[17:57])
    defparam i46364_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i13283_3_lut (.I0(baudrate[10]), .I1(data_adj_5899[2]), .I2(n55526), 
            .I3(GND_net), .O(n29128));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13283_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13284_3_lut (.I0(baudrate[9]), .I1(data_adj_5899[1]), .I2(n55526), 
            .I3(GND_net), .O(n29129));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13284_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13331_4_lut_4_lut (.I0(n27441), .I1(state[1]), .I2(bit_ctr[1]), 
            .I3(bit_ctr[0]), .O(n29176));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13331_4_lut_4_lut.LUT_INIT = 16'h5270;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5691));   // verilog/TinyFPGA_B.v(332[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12797_2_lut_3_lut (.I0(n22471), .I1(dti), .I2(n15_adj_5741), 
            .I3(GND_net), .O(n28642));
    defparam i12797_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i13161_3_lut (.I0(\data_in_frame[6] [1]), .I1(rx_data[1]), .I2(n27904), 
            .I3(GND_net), .O(n29006));   // verilog/coms.v(130[12] 305[6])
    defparam i13161_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut_adj_2008 (.I0(n22471), .I1(dti), .I2(n15_adj_5741), 
            .I3(GND_net), .O(n27460));
    defparam i1_2_lut_3_lut_adj_2008.LUT_INIT = 16'hf8f8;
    SB_LUT4 i13285_3_lut (.I0(baudrate[8]), .I1(data_adj_5899[0]), .I2(n55526), 
            .I3(GND_net), .O(n29130));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13285_3_lut.LUT_INIT = 16'hacac;
    TLI4970 tli (.state_7__N_4319(state_7__N_4319), .GND_net(GND_net), .clk16MHz(clk16MHz), 
            .CS_c(CS_c), .CS_CLK_c(CS_CLK_c), .VCC_net(VCC_net), .n27290(n27290), 
            .\current[15] (current[15]), .n29106(n29106), .\current[1] (current[1]), 
            .n29105(n29105), .\current[2] (current[2]), .n29104(n29104), 
            .\current[3] (current[3]), .n29103(n29103), .\current[4] (current[4]), 
            .n29102(n29102), .\current[5] (current[5]), .n29101(n29101), 
            .\current[6] (current[6]), .n29100(n29100), .\current[7] (current[7]), 
            .n29099(n29099), .\current[8] (current[8]), .n29098(n29098), 
            .\current[9] (current[9]), .n29097(n29097), .\current[10] (current[10]), 
            .n29096(n29096), .\current[11] (current[11]), .n29826(n29826), 
            .\data[15] (data_adj_5906[15]), .n29825(n29825), .\data[12] (data_adj_5906[12]), 
            .n29824(n29824), .\data[11] (data_adj_5906[11]), .n29823(n29823), 
            .\data[10] (data_adj_5906[10]), .n29822(n29822), .\data[9] (data_adj_5906[9]), 
            .n29821(n29821), .\data[8] (data_adj_5906[8]), .n29820(n29820), 
            .\data[7] (data_adj_5906[7]), .n29819(n29819), .\data[6] (data_adj_5906[6]), 
            .n29818(n29818), .\data[5] (data_adj_5906[5]), .n29817(n29817), 
            .\data[4] (data_adj_5906[4]), .n29816(n29816), .\data[3] (data_adj_5906[3]), 
            .n29815(n29815), .\data[2] (data_adj_5906[2]), .n29814(n29814), 
            .\data[1] (data_adj_5906[1]), .n29600(n29600), .\data[0] (data_adj_5906[0]), 
            .n28927(n28927), .\current[0] (current[0]), .n5(n5_adj_5761), 
            .n11(n11_adj_5747), .n25130(n25130), .n25133(n25133), .n5_adj_21(n5_adj_5746), 
            .n5_adj_22(n5_adj_5771), .n38316(n38316), .n25141(n25141), 
            .n25110(n25110)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(413[11] 419[4])
    SB_LUT4 i13583_3_lut (.I0(\data_in_frame[18] [3]), .I1(rx_data[3]), 
            .I2(n27929), .I3(GND_net), .O(n29428));   // verilog/coms.v(130[12] 305[6])
    defparam i13583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13286_3_lut (.I0(baudrate[7]), .I1(data_adj_5899[7]), .I2(n55533), 
            .I3(GND_net), .O(n29131));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13286_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1956_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n1325), .I3(n38194), .O(n6911));   // verilog/TinyFPGA_B.v(370[5] 396[12])
    defparam i1956_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 i9_2_lut (.I0(PWMLimit[12]), .I1(setpoint[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5791));   // verilog/TinyFPGA_B.v(250[22:30])
    defparam i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13287_3_lut (.I0(baudrate[6]), .I1(data_adj_5899[6]), .I2(n55533), 
            .I3(GND_net), .O(n29132));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13287_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i9_2_lut_adj_2009 (.I0(PWMLimit[10]), .I1(setpoint[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5790));   // verilog/TinyFPGA_B.v(250[22:30])
    defparam i9_2_lut_adj_2009.LUT_INIT = 16'h6666;
    SB_LUT4 i13288_3_lut (.I0(baudrate[5]), .I1(data_adj_5899[5]), .I2(n55533), 
            .I3(GND_net), .O(n29133));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13288_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13289_3_lut (.I0(baudrate[4]), .I1(data_adj_5899[4]), .I2(n55533), 
            .I3(GND_net), .O(n29134));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13289_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i18014_3_lut (.I0(n36), .I1(PWMLimit[18]), .I2(setpoint[18]), 
            .I3(GND_net), .O(n33833));   // verilog/TinyFPGA_B.v(250[22:30])
    defparam i18014_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i13290_3_lut (.I0(baudrate[3]), .I1(data_adj_5899[3]), .I2(n55533), 
            .I3(GND_net), .O(n29135));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13290_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17971_3_lut (.I0(n40), .I1(PWMLimit[20]), .I2(setpoint[20]), 
            .I3(GND_net), .O(n33791));   // verilog/TinyFPGA_B.v(250[22:30])
    defparam i17971_3_lut.LUT_INIT = 16'hb2b2;
    SB_LUT4 i13291_3_lut (.I0(baudrate[2]), .I1(data_adj_5899[2]), .I2(n55533), 
            .I3(GND_net), .O(n29136));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13291_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13292_3_lut (.I0(baudrate[1]), .I1(data_adj_5899[1]), .I2(n55533), 
            .I3(GND_net), .O(n29137));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13292_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13293_3_lut (.I0(baudrate[0]), .I1(data_adj_5899[0]), .I2(n55533), 
            .I3(GND_net), .O(n29138));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13293_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13294_3_lut (.I0(ID[7]), .I1(data_adj_5899[7]), .I2(n55524), 
            .I3(GND_net), .O(n29139));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13294_3_lut.LUT_INIT = 16'hacac;
    \quadrature_decoder(0)  quad_counter1 (.ENCODER1_B_N_keep(ENCODER1_B_N), 
            .n1795(clk16MHz), .ENCODER1_A_N_keep(ENCODER1_A_N), .b_prev(b_prev_adj_5752), 
            .\a_new[1] (a_new_adj_5885[1]), .GND_net(GND_net), .encoder1_position({encoder1_position}), 
            .VCC_net(VCC_net), .\b_new[1] (b_new_adj_5886[1]), .n29064(n29064), 
            .a_prev(a_prev_adj_5751), .position_31__N_3836(position_31__N_3836_adj_5754), 
            .n28938(n28938), .n28937(n28937), .n1800(n1800), .debounce_cnt_N_3833(debounce_cnt_N_3833_adj_5753)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(321[27] 327[6])
    SB_LUT4 i13295_3_lut (.I0(ID[6]), .I1(data_adj_5899[6]), .I2(n55524), 
            .I3(GND_net), .O(n29140));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13295_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13296_3_lut (.I0(ID[5]), .I1(data_adj_5899[5]), .I2(n55524), 
            .I3(GND_net), .O(n29141));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13296_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13297_3_lut (.I0(ID[4]), .I1(data_adj_5899[4]), .I2(n55524), 
            .I3(GND_net), .O(n29142));   // verilog/eeprom.v(35[8] 81[4])
    defparam i13297_3_lut.LUT_INIT = 16'hacac;
    coms neopxl_color_23__I_0 (.n2882(n2882), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .clk16MHz(clk16MHz), .n55292(n55292), .n29434(n29434), .VCC_net(VCC_net), 
         .\data_in_frame[18] ({\data_in_frame[18] }), .n55291(n55291), .n55290(n55290), 
         .n29431(n29431), .n55289(n55289), .n55288(n55288), .n55242(n55242), 
         .n55287(n55287), .\data_out_frame[9] ({\data_out_frame[9] }), .\FRAME_MATCHER.i_31__N_2509 (\FRAME_MATCHER.i_31__N_2509 ), 
         .encoder1_position_scaled({encoder1_position_scaled}), .n8(n8_adj_5789), 
         .rx_data({rx_data}), .\data_in_frame[2] ({Open_3, Open_4, Open_5, 
         Open_6, Open_7, Open_8, Open_9, \data_in_frame[2] [0]}), 
         .\data_in_frame[12] ({\data_in_frame[12] }), .IntegralLimit({IntegralLimit}), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .n55286(n55286), 
         .n55285(n55285), .n55284(n55284), .n55283(n55283), .n55282(n55282), 
         .\data_out_frame[3][1] (\data_out_frame[3] [1]), .n55409(n55409), 
         .\data_out_frame[8][7] (\data_out_frame[8] [7]), .\encoder0_position_scaled[7] (encoder0_position_scaled[7]), 
         .n55281(n55281), .n55280(n55280), .n55279(n55279), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .n55278(n55278), .\data_out_frame[8][6] (\data_out_frame[8] [6]), 
         .\encoder0_position_scaled[6] (encoder0_position_scaled[6]), .\data_out_frame[3][3] (\data_out_frame[3] [3]), 
         .n55408(n55408), .n29428(n29428), .\data_out_frame[3][4] (\data_out_frame[3] [4]), 
         .n55407(n55407), .\data_out_frame[8][5] (\data_out_frame[8] [5]), 
         .\encoder0_position_scaled[5] (encoder0_position_scaled[5]), .n55277(n55277), 
         .\data_out_frame[3][6] (\data_out_frame[3] [6]), .n55406(n55406), 
         .n29006(n29006), .\data_in_frame[6] ({Open_10, Open_11, Open_12, 
         \data_in_frame[6] [4:1], Open_13}), .\data_out_frame[3][7] (\data_out_frame[3] [7]), 
         .n55405(n55405), .n55276(n55276), .\data_out_frame[8][4] (\data_out_frame[8] [4]), 
         .\encoder0_position_scaled[4] (encoder0_position_scaled[4]), .\data_out_frame[8][3] (\data_out_frame[8] [3]), 
         .\encoder0_position_scaled[3] (encoder0_position_scaled[3]), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .\data_out_frame[8][2] (\data_out_frame[8] [2]), .\encoder0_position_scaled[2] (encoder0_position_scaled[2]), 
         .n55275(n55275), .n55274(n55274), .\data_out_frame[7] ({\data_out_frame[7] }), 
         .\encoder0_position_scaled[15] (encoder0_position_scaled[15]), .n28729(n28729), 
         .n55273(n55273), .n55272(n55272), .\data_out_frame[21] ({\data_out_frame[21] }), 
         .n55271(n55271), .n55270(n55270), .n55269(n55269), .n55268(n55268), 
         .\data_out_frame[1][7] (\data_out_frame[1] [7]), .GND_net(GND_net), 
         .n55267(n55267), .n28721(n28721), .n55241(n55241), .n55266(n55266), 
         .\data_out_frame[1][6] (\data_out_frame[1] [6]), .\data_out_frame[22] ({\data_out_frame[22] }), 
         .n55265(n55265), .n55264(n55264), .n55263(n55263), .n55262(n55262), 
         .n55261(n55261), .n28713(n28713), .n29424(n29424), .\data_out_frame[4] ({\data_out_frame[4] }), 
         .n55404(n55404), .n55403(n55403), .\data_out_frame[1][5] (\data_out_frame[1] [5]), 
         .\data_out_frame[1][3] (\data_out_frame[1] [3]), .\data_out_frame[1][1] (\data_out_frame[1] [1]), 
         .n29421(n29421), .n55260(n55260), .n28711(n28711), .\data_out_frame[1][0] (\data_out_frame[1] [0]), 
         .\data_out_frame[0][4] (\data_out_frame[0] [4]), .\data_out_frame[0][3] (\data_out_frame[0] [3]), 
         .\data_out_frame[0][2] (\data_out_frame[0] [2]), .\data_out_frame[23] ({\data_out_frame[23] }), 
         .n55259(n55259), .\data_in_frame[21] ({\data_in_frame[21] [7], 
         Open_14, Open_15, Open_16, Open_17, Open_18, Open_19, Open_20}), 
         .n27934(n27934), .n55419(n55419), .n55402(n55402), .displacement({displacement}), 
         .n55401(n55401), .n29418(n29418), .n55400(n55400), .n55399(n55399), 
         .n55398(n55398), .n29415(n29415), .\data_in_frame[17] ({\data_in_frame[17] [7], 
         Open_21, Open_22, Open_23, Open_24, Open_25, Open_26, Open_27}), 
         .\data_out_frame[5] ({\data_out_frame[5] }), .n55397(n55397), .n55396(n55396), 
         .n29409(n29409), .\data_in_frame[17][5] (\data_in_frame[17] [5]), 
         .n29406(n29406), .\data_in_frame[17][4] (\data_in_frame[17] [4]), 
         .n55395(n55395), .n29403(n29403), .\data_in_frame[17][3] (\data_in_frame[17] [3]), 
         .n55300(n55300), .n29400(n29400), .\data_in_frame[17][2] (\data_in_frame[17] [2]), 
         .n55394(n55394), .n29397(n29397), .\data_in_frame[17][1] (\data_in_frame[17] [1]), 
         .n55393(n55393), .n55258(n55258), .n55257(n55257), .n55256(n55256), 
         .n28706(n28706), .n55392(n55392), .n55255(n55255), .n55391(n55391), 
         .n55254(n55254), .n29394(n29394), .\data_in_frame[17][0] (\data_in_frame[17] [0]), 
         .n28703(n28703), .\data_out_frame[6] ({\data_out_frame[6] }), .n55390(n55390), 
         .\data_out_frame[24] ({\data_out_frame[24] }), .n55301(n55301), 
         .n29009(n29009), .n55389(n55389), .n29392(n29392), .\data_in_frame[16] ({\data_in_frame[16] }), 
         .n55388(n55388), .n29389(n29389), .n55387(n55387), .n29384(n29384), 
         .n55386(n55386), .deadband({deadband}), .n55253(n55253), .\data_in_frame[14][6] (\data_in_frame[14] [6]), 
         .n55252(n55252), .n55251(n55251), .n29381(n29381), .n55250(n55250), 
         .n55249(n55249), .n28696(n28696), .n55299(n55299), .\data_out_frame[25] ({\data_out_frame[25] }), 
         .n55248(n55248), .n55247(n55247), .\data_in_frame[20] ({\data_in_frame[20] }), 
         .n27932(n27932), .n29378(n29378), .n55246(n55246), .n55245(n55245), 
         .n55244(n55244), .n28689(n28689), .n55385(n55385), .\encoder0_position_scaled[11] (encoder0_position_scaled[11]), 
         .\data_in_frame[15] ({\data_in_frame[15] }), .n28688(n28688), .\encoder0_position_scaled[10] (encoder0_position_scaled[10]), 
         .n55243(n55243), .\data_out_frame[26] ({\data_out_frame[26] }), 
         .n55454(n55454), .n55453(n55453), .n55384(n55384), .n55452(n55452), 
         .n55451(n55451), .n55450(n55450), .n55445(n55445), .byte_transmit_counter({Open_28, 
         Open_29, Open_30, Open_31, Open_32, byte_transmit_counter[2:0]}), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .n28680(n28680), .n55455(n55455), .\data_out_frame[27] ({\data_out_frame[27] }), 
         .n55446(n55446), .n55447(n55447), .n55448(n55448), .n55449(n55449), 
         .n55443(n55443), .reset(reset), .n55444(n55444), .n29012(n29012), 
         .n27898(n27898), .setpoint({setpoint}), .n28672(n28672), .n29374(n29374), 
         .\r_SM_Main_2__N_3545[0] (r_SM_Main_2__N_3545[0]), .tx_active(tx_active), 
         .n53(n53), .n55456(n55456), .\encoder0_position_scaled[9] (encoder0_position_scaled[9]), 
         .\FRAME_MATCHER.i[3] (\FRAME_MATCHER.i [3]), .\FRAME_MATCHER.i[4] (\FRAME_MATCHER.i [4]), 
         .\encoder0_position_scaled[8] (encoder0_position_scaled[8]), .\FRAME_MATCHER.i[5] (\FRAME_MATCHER.i [5]), 
         .\byte_transmit_counter[5] (byte_transmit_counter[5]), .\byte_transmit_counter[6] (byte_transmit_counter[6]), 
         .\byte_transmit_counter[7] (byte_transmit_counter[7]), .n29371(n29371), 
         .n55383(n55383), .n29368(n29368), .\encoder0_position_scaled[14] (encoder0_position_scaled[14]), 
         .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), .n8_adj_4(n8_adj_5711), 
         .n56368(n56368), .n29365(n29365), .\data_in_frame[19] ({Open_33, 
         Open_34, Open_35, Open_36, Open_37, \data_in_frame[19] [2:1], 
         Open_38}), .n55382(n55382), .n58202(n58202), .n29362(n29362), 
         .n55381(n55381), .\FRAME_MATCHER.i[0] (\FRAME_MATCHER.i [0]), .\data_in_frame[3][3] (\data_in_frame[3] [3]), 
         .n29359(n29359), .n29356(n29356), .n29353(n29353), .n29015(n29015), 
         .n29349(n29349), .n55380(n55380), .n3484(n3484), .n29346(n29346), 
         .n55379(n55379), .n29343(n29343), .\data_in_frame[3][5] (\data_in_frame[3] [5]), 
         .\data_in_frame[3][6] (\data_in_frame[3] [6]), .\data_in_frame[1] ({\data_in_frame[1] [7:4], 
         Open_39, Open_40, Open_41, \data_in_frame[1] [0]}), .\encoder0_position_scaled[23] (encoder0_position_scaled[23]), 
         .\data_in_frame[3][0] (\data_in_frame[3] [0]), .\data_in_frame[19][0] (\data_in_frame[19] [0]), 
         .n29316(n29316), .n29313(n29313), .n29309(n29309), .n29306(n29306), 
         .n29303(n29303), .n29300(n29300), .n29297(n29297), .n55378(n55378), 
         .n29294(n29294), .n29291(n29291), .n29288(n29288), .n29285(n29285), 
         .n29282(n29282), .\data_in_frame[6][6] (\data_in_frame[6] [6]), 
         .n29278(n29278), .n29275(n29275), .n29272(n29272), .n29269(n29269), 
         .n29266(n29266), .\data_in_frame[11] ({\data_in_frame[11] }), .n29263(n29263), 
         .n29024(n29024), .\data_in_frame[6][7] (\data_in_frame[6] [7]), 
         .n29258(n29258), .n29255(n29255), .n29252(n29252), .n55377(n55377), 
         .n29249(n29249), .n29246(n29246), .n29243(n29243), .n29030(n29030), 
         .\data_in_frame[7][1] (\data_in_frame[7] [1]), .n29033(n29033), 
         .\data_in_frame[7][2] (\data_in_frame[7] [2]), .n29042(n29042), 
         .\data_in_frame[7][4] (\data_in_frame[7] [4]), .\data_in_frame[3][7] (\data_in_frame[3] [7]), 
         .n29045(n29045), .\data_in_frame[7][5] (\data_in_frame[7] [5]), 
         .n29048(n29048), .\data_in_frame[7][6] (\data_in_frame[7] [6]), 
         .n29051(n29051), .\data_in_frame[7][7] (\data_in_frame[7] [7]), 
         .n66714(n66714), .n55302(n55302), .n66702(n66702), .n56366(n56366), 
         .n56162(n56162), .n56050(n56050), .n27906(n27906), .\data_in_frame[21][1] (\data_in_frame[21] [1]), 
         .n25895(n25895), .n55418(n55418), .n55417(n55417), .n55416(n55416), 
         .n55415(n55415), .n55414(n55414), .n55413(n55413), .n55412(n55412), 
         .n55411(n55411), .n55410(n55410), .n55376(n55376), .n55303(n55303), 
         .n55375(n55375), .n55374(n55374), .n55373(n55373), .n55372(n55372), 
         .n55371(n55371), .n55370(n55370), .n55369(n55369), .n55368(n55368), 
         .n55367(n55367), .n55366(n55366), .n55365(n55365), .n55364(n55364), 
         .n55363(n55363), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .n55362(n55362), .n55361(n55361), .n55360(n55360), .n55359(n55359), 
         .n55358(n55358), .n55357(n55357), .n55356(n55356), .n55355(n55355), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .n55354(n55354), 
         .n55353(n55353), .n55352(n55352), .n55351(n55351), .n55350(n55350), 
         .n55349(n55349), .n55348(n55348), .n55347(n55347), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .n55346(n55346), .n55345(n55345), .n55344(n55344), .n55343(n55343), 
         .n55342(n55342), .n55341(n55341), .n55340(n55340), .n55339(n55339), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .n55338(n55338), 
         .n55337(n55337), .n55336(n55336), .n55335(n55335), .n55334(n55334), 
         .n55333(n55333), .n55332(n55332), .n55331(n55331), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .n55330(n55330), .n55329(n55329), .n55328(n55328), .n55327(n55327), 
         .n55326(n55326), .n55325(n55325), .n55305(n55305), .n55324(n55324), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .n55323(n55323), 
         .n55322(n55322), .n55321(n55321), .n55320(n55320), .n55319(n55319), 
         .n55318(n55318), .n55317(n55317), .n55304(n55304), .n55316(n55316), 
         .n55315(n55315), .n55314(n55314), .n55313(n55313), .n55312(n55312), 
         .n29061(n29061), .\FRAME_MATCHER.rx_data_ready_prev (\FRAME_MATCHER.rx_data_ready_prev ), 
         .n55311(n55311), .n55310(n55310), .n55309(n55309), .n55308(n55308), 
         .n55307(n55307), .n55306(n55306), .n55298(n55298), .n55297(n55297), 
         .n55296(n55296), .n55295(n55295), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .LED_c(LED_c), .n56120(n56120), .n55985(n55985), .DE_c(DE_c), 
         .n55294(n55294), .\data_in_frame[0] ({\data_in_frame[0] [7], Open_42, 
         Open_43, Open_44, Open_45, Open_46, Open_47, Open_48}), 
         .n50260(n50260), .n24804(n24804), .n25941(n25941), .n55648(n55648), 
         .\data_in_frame[6][0] (\data_in_frame[6] [0]), .Kp_23__N_875(Kp_23__N_875), 
         .n50264(n50264), .n55624(n55624), .n55775(n55775), .\data_in_frame[21][2] (\data_in_frame[21] [2]), 
         .n25705(n25705), .n32987(n32987), .\data_in_frame[21][3] (\data_in_frame[21] [3]), 
         .n25490(n25490), .n55681(n55681), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .n56062(n56062), .n27900(n27900), .n29437(n29437), .\encoder0_position_scaled[13] (encoder0_position_scaled[13]), 
         .n29440(n29440), .n28912(n28912), .n29468(n29468), .n29477(n29477), 
         .n29481(n29481), .n29484(n29484), .n29487(n29487), .n29493(n29493), 
         .\data_in_frame[21][0] (\data_in_frame[21] [0]), .n29496(n29496), 
         .n29499(n29499), .n29506(n29506), .n29509(n29509), .\data_in_frame[21][4] (\data_in_frame[21] [4]), 
         .n29512(n29512), .\data_in_frame[21][5] (\data_in_frame[21] [5]), 
         .\data_in_frame[0][4] (\data_in_frame[0] [4]), .n29546(n29546), 
         .\data_in_frame[23] ({Open_49, \data_in_frame[23] [6:0]}), .n29549(n29549), 
         .n29552(n29552), .n29555(n29555), .n29558(n29558), .n54697(n54697), 
         .n54695(n54695), .n28940(n28940), .n28946(n28946), .n28949(n28949), 
         .n28952(n28952), .n54733(n54733), .n28958(n28958), .\Kp[1] (Kp[1]), 
         .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), 
         .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), 
         .\Kp[10] (Kp[10]), .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .\Kp[13] (Kp[13]), 
         .\Kp[14] (Kp[14]), .\Kp[15] (Kp[15]), .\Ki[1] (Ki[1]), .\Ki[2] (Ki[2]), 
         .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), 
         .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), 
         .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), 
         .\Ki[15] (Ki[15]), .n29677(n29677), .neopxl_color({neopxl_color}), 
         .n29676(n29676), .n28961(n28961), .n29674(n29674), .n29673(n29673), 
         .n29671(n29671), .n29670(n29670), .n29669(n29669), .n29668(n29668), 
         .n29667(n29667), .n29666(n29666), .n29665(n29665), .n29664(n29664), 
         .n29662(n29662), .n29661(n29661), .n29660(n29660), .n29659(n29659), 
         .n29658(n29658), .n29657(n29657), .n29656(n29656), .n29655(n29655), 
         .n29654(n29654), .control_mode({control_mode}), .n29650(n29650), 
         .n29649(n29649), .n29648(n29648), .n29647(n29647), .n29646(n29646), 
         .current_limit({current_limit}), .n29645(n29645), .n29644(n29644), 
         .n29643(n29643), .n29642(n29642), .n29640(n29640), .n29638(n29638), 
         .n29637(n29637), .n29636(n29636), .n29635(n29635), .n29634(n29634), 
         .n29633(n29633), .n29632(n29632), .PWMLimit({PWMLimit}), .n28964(n28964), 
         .n28967(n28967), .n28976(n28976), .n55293(n55293), .n28982(n28982), 
         .ID({ID}), .n28988(n28988), .n28991(n28991), .n28994(n28994), 
         .n28997(n28997), .n28923(n28923), .n28922(n28922), .n28921(n28921), 
         .\Ki[0] (Ki[0]), .\Kp[0] (Kp[0]), .n29000(n29000), .n29003(n29003), 
         .n56059(n56059), .n63134(n63134), .n27904(n27904), .n25933(n25933), 
         .n55668(n55668), .pwm_setpoint({pwm_setpoint}), .\encoder0_position_scaled[12] (encoder0_position_scaled[12]), 
         .n57376(n57376), .n27513(n27513), .n66672(n66672), .n66654(n66654), 
         .n50946(n50946), .n56231(n56231), .n56201(n56201), .n24633(n24633), 
         .n56165(n56165), .n22318(n22318), .n50377(n50377), .n66864(n66864), 
         .n66618(n66618), .n56183(n56183), .Kp_23__N_748(Kp_23__N_748), 
         .\encoder0_position_scaled[22] (encoder0_position_scaled[22]), .n73(n73), 
         .rx_data_ready(rx_data_ready), .n51197(n51197), .n51161(n51161), 
         .n51296(n51296), .n37097(n37097), .n27926(n27926), .n27902(n27902), 
         .n55952(n55952), .n55152(n55152), .n56109(n56109), .n22369(n22369), 
         .n50927(n50927), .n50183(n50183), .n25803(n25803), .n26439(n26439), 
         .n51232(n51232), .n55884(n55884), .n27939(n27939), .n55989(n55989), 
         .n63131(n63131), .n25494(n25494), .n4(n4_adj_5836), .n55181(n55181), 
         .n105(n105), .control_update(control_update), .n7064(n7064), 
         .n38328(n38328), .n24981(n24981), .n38638(n38638), .n6(n6_adj_5825), 
         .n55149(n55149), .n10(n10_adj_5745), .n15(n15_adj_5770), .n27260(n27260), 
         .n15_adj_5(n15_adj_5748), .n15_adj_6(n15_adj_5712), .n55766(n55766), 
         .n56024(n56024), .n38266(n38266), .n38695(n38695), .\encoder0_position_scaled[21] (encoder0_position_scaled[21]), 
         .\encoder0_position_scaled[20] (encoder0_position_scaled[20]), .\encoder0_position_scaled[19] (encoder0_position_scaled[19]), 
         .\encoder0_position_scaled[18] (encoder0_position_scaled[18]), .\encoder0_position_scaled[17] (encoder0_position_scaled[17]), 
         .n50591(n50591), .\encoder0_position_scaled[16] (encoder0_position_scaled[16]), 
         .n55151(n55151), .n57943(n57943), .\current[7] (current[7]), 
         .\current[6] (current[6]), .n55587(n55587), .\current[5] (current[5]), 
         .\current[4] (current[4]), .\current[3] (current[3]), .\current[2] (current[2]), 
         .\current[1] (current[1]), .\current[0] (current[0]), .\current[15] (current[15]), 
         .n55153(n55153), .n60056(n60056), .n60054(n60054), .\current[11] (current[11]), 
         .\current[10] (current[10]), .\current[9] (current[9]), .\current[8] (current[8]), 
         .\r_SM_Main[1] (r_SM_Main_adj_5922[1]), .r_Clock_Count({r_Clock_Count_adj_5923}), 
         .n39972(n39972), .tx_o(tx_o), .n20722(n20722), .\r_SM_Main[0] (r_SM_Main_adj_5922[0]), 
         .n27315(n27315), .n23(n23_adj_5830), .\o_Rx_DV_N_3488[12] (o_Rx_DV_N_3488[12]), 
         .n5228(n5228), .\o_Rx_DV_N_3488[24] (o_Rx_DV_N_3488[24]), .n27(n27), 
         .n29(n29), .n39919(n39919), .n29589(n29589), .\r_Bit_Index[0] (r_Bit_Index_adj_5924[0]), 
         .n51433(n51433), .n39937(n39937), .n57036(n57036), .n31(n31), 
         .n58374(n58374), .n58502(n58502), .o_Tx_Serial_N_3598(o_Tx_Serial_N_3598), 
         .tx_enable(tx_enable), .baudrate({baudrate}), .r_SM_Main({r_SM_Main}), 
         .r_Rx_Data(r_Rx_Data), .RX_N_2(RX_N_2), .r_Clock_Count_adj_20({r_Clock_Count}), 
         .n25108(n25108), .n5225(n5225), .\o_Rx_DV_N_3488[8] (o_Rx_DV_N_3488[8]), 
         .\o_Rx_DV_N_3488[7] (o_Rx_DV_N_3488[7]), .\o_Rx_DV_N_3488[6] (o_Rx_DV_N_3488[6]), 
         .\o_Rx_DV_N_3488[5] (o_Rx_DV_N_3488[5]), .\o_Rx_DV_N_3488[4] (o_Rx_DV_N_3488[4]), 
         .\o_Rx_DV_N_3488[3] (o_Rx_DV_N_3488[3]), .\o_Rx_DV_N_3488[2] (o_Rx_DV_N_3488[2]), 
         .\o_Rx_DV_N_3488[1] (o_Rx_DV_N_3488[1]), .\o_Rx_DV_N_3488[0] (o_Rx_DV_N_3488[0]), 
         .n27312(n27312), .n29592(n29592), .\r_Bit_Index[0]_adj_17 (r_Bit_Index[0]), 
         .n51425(n51425), .n29596(n29596), .n29582(n29582), .n29581(n29581), 
         .n29580(n29580), .n29578(n29578), .n29577(n29577), .n29576(n29576), 
         .n29575(n29575), .\r_SM_Main_2__N_3446[1] (r_SM_Main_2__N_3446[1]), 
         .n56281(n56281), .n6_adj_18(n6_adj_5838), .n55184(n55184), .n58618(n58618), 
         .n4_adj_19(n4_adj_5744), .n27308(n27308), .n58594(n58594), .n58896(n58896), 
         .n58898(n58898), .n58932(n58932), .n58844(n58844), .n58970(n58970), 
         .n58934(n58934), .n58880(n58880), .n58952(n58952)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(263[22] 288[4])
    SB_LUT4 unary_minus_15_inv_0_i24_1_lut (.I0(duty[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_setpoint_23__N_207));   // verilog/TinyFPGA_B.v(127[24:29])
    defparam unary_minus_15_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    EEPROM eeprom (.GND_net(GND_net), .enable_slow_N_4213(enable_slow_N_4213), 
           .clk16MHz(clk16MHz), .\state_7__N_4110[0] (state_7__N_4110[0]), 
           .n29153(n29153), .ID({ID}), .n29152(n29152), .n29143(n29143), 
           .n29142(n29142), .n29141(n29141), .n29140(n29140), .n29139(n29139), 
           .n29138(n29138), .baudrate({baudrate}), .n29137(n29137), .n29136(n29136), 
           .n29135(n29135), .n29134(n29134), .n29133(n29133), .n29132(n29132), 
           .n29131(n29131), .n29130(n29130), .n29129(n29129), .n29128(n29128), 
           .n29127(n29127), .n29126(n29126), .n29125(n29125), .n29124(n29124), 
           .n29123(n29123), .n29114(n29114), .n29113(n29113), .n29112(n29112), 
           .n29111(n29111), .n29110(n29110), .n29109(n29109), .n29108(n29108), 
           .n29107(n29107), .data_ready(data_ready), .n28925(n28925), 
           .n55526(n55526), .n55533(n55533), .\state_7__N_3918[0] (state_7__N_3918[0]), 
           .data({data_adj_5899}), .n55524(n55524), .n57999(n57999), .n25095(n25095), 
           .VCC_net(VCC_net), .n38386(n38386), .scl_enable(scl_enable), 
           .\state[0] (state_adj_5935[0]), .n29156(n29156), .scl(scl), 
           .sda_enable(sda_enable), .sda_out(sda_out), .n29812(n29812), 
           .n29811(n29811), .n29810(n29810), .n29809(n29809), .n29808(n29808), 
           .n29806(n29806), .n29586(n29586), .n6(n6_adj_5842), .n6715(n6715), 
           .n10(n10_adj_5812), .\state_7__N_4126[3] (state_7__N_4126[3]), 
           .n38223(n38223), .n38221(n38221), .n4(n4_adj_5742), .n25100(n25100), 
           .n4_adj_3(n4_adj_5743)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(399[10] 411[6])
    pwm PWM (.n2882(n2882), .pwm_out(pwm_out), .clk32MHz(clk32MHz), .GND_net(GND_net), 
        .VCC_net(VCC_net), .pwm_setpoint({pwm_setpoint}), .reset(reset)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(105[6] 110[3])
    motorControl control (.GND_net(GND_net), .\Ki[2] (Ki[2]), .n335({n336, 
            n337, n338, n339, n340, n341, n342, n343, n344, 
            n345, n346, n347, n348, n349, n350, n351, n352, 
            n353, n354, n355, n356, n357, n358, n359}), .setpoint({setpoint}), 
            .deadband({deadband}), .\Ki[3] (Ki[3]), .\Kp[7] (Kp[7]), .IntegralLimit({IntegralLimit}), 
            .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), 
            .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), 
            .\Kp[6] (Kp[6]), .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), 
            .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .\Kp[13] (Kp[13]), .\Kp[14] (Kp[14]), 
            .\Ki[6] (Ki[6]), .\Kp[15] (Kp[15]), .\encoder1_position_scaled[0] (encoder1_position_scaled[0]), 
            .n15(n15_adj_5748), .n62934(n62934), .n15_adj_1(n15_adj_5712), 
            .\encoder1_position_scaled[1] (encoder1_position_scaled[1]), .n62948(n62948), 
            .\motor_state[9] (motor_state[9]), .control_update(control_update), 
            .duty({duty}), .clk16MHz(clk16MHz), .reset(reset), .\motor_state[8] (motor_state[8]), 
            .\Ki[1] (Ki[1]), .\Ki[0] (Ki[0]), .PWMLimit({PWMLimit}), .\Ki[7] (Ki[7]), 
            .\Ki[8] (Ki[8]), .\Ki[9] (Ki[9]), .\motor_state[7] (motor_state[7]), 
            .VCC_net(VCC_net), .\motor_state[6] (motor_state[6]), .\Ki[10] (Ki[10]), 
            .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), .\Ki[13] (Ki[13]), .\motor_state[5] (motor_state[5]), 
            .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), .\motor_state[4] (motor_state[4]), 
            .\motor_state[10] (motor_state[10]), .\motor_state[3] (motor_state[3]), 
            .n3(n3_adj_5811), .control_mode({control_mode}), .n55181(n55181), 
            .n105(n105), .n7064(n7064), .n38638(n38638), .n29778(n29778), 
            .\PID_CONTROLLER.integral ({\PID_CONTROLLER.integral }), .n29777(n29777), 
            .n29776(n29776), .n29775(n29775), .n29774(n29774), .n29773(n29773), 
            .n29772(n29772), .n29771(n29771), .n29770(n29770), .n29769(n29769), 
            .n29768(n29768), .n29767(n29767), .n29766(n29766), .n29765(n29765), 
            .n29764(n29764), .n29763(n29763), .n29762(n29762), .n29761(n29761), 
            .n29760(n29760), .n29759(n29759), .n29758(n29758), .n29757(n29757), 
            .n29754(n29754), .n28910(n28910), .\motor_state[23] (motor_state[23]), 
            .\motor_state[22] (motor_state[22]), .\motor_state[21] (motor_state[21]), 
            .\motor_state[20] (motor_state[20]), .\motor_state[19] (motor_state[19]), 
            .\motor_state[18] (motor_state[18]), .\motor_state[17] (motor_state[17]), 
            .\motor_state[16] (motor_state[16]), .\motor_state[15] (motor_state[15]), 
            .n9(n9_adj_5792), .\motor_state[13] (motor_state[13]), .\motor_state[12] (motor_state[12]), 
            .\motor_state[11] (motor_state[11]), .n38659(n38659), .n24981(n24981), 
            .n38328(n38328), .n21(n21_adj_5790), .n25(n25_adj_5791), .n36(n36), 
            .n33833(n33833), .n40(n40), .n33791(n33791)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(298[16] 311[4])
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (clk16MHz, bit_ctr, GND_net, 
            state, n3173, neopxl_color, t0, n23, n38711, timer, 
            n35156, n27441, VCC_net, n29176, n5, n29155, n29154, 
            n29151, n29150, n29149, n29148, n29147, n29146, n29145, 
            n29144, NEOPXL_c, n28939, \data_in_frame[4][2] , \data_in_frame[4][3] , 
            n56059, \data_in_frame[1][6] , \data_in_frame[1][7] , n55668, 
            n56216, n25933, Kp_23__N_875, \data_out_frame[23][2] , \data_out_frame[23][3] , 
            n55952, \data_out_frame[24][7] , n50377, n56165, \rx_data[3] , 
            n27900, n28964, n22369, n29658, n29659, LED_c, n24633, 
            \data_out_frame[21][0] , n56162, \data_in_frame[2][0] ) /* synthesis syn_module_defined=1 */ ;
    input clk16MHz;
    output [4:0]bit_ctr;
    input GND_net;
    output [1:0]state;
    output n3173;
    input [23:0]neopxl_color;
    output [10:0]t0;
    output n23;
    output n38711;
    output [10:0]timer;
    output n35156;
    output n27441;
    input VCC_net;
    input n29176;
    input n5;
    input n29155;
    input n29154;
    input n29151;
    input n29150;
    input n29149;
    input n29148;
    input n29147;
    input n29146;
    input n29145;
    input n29144;
    output NEOPXL_c;
    input n28939;
    input \data_in_frame[4][2] ;
    input \data_in_frame[4][3] ;
    output n56059;
    input \data_in_frame[1][6] ;
    input \data_in_frame[1][7] ;
    output n55668;
    output n56216;
    input n25933;
    output Kp_23__N_875;
    input \data_out_frame[23][2] ;
    input \data_out_frame[23][3] ;
    output n55952;
    input \data_out_frame[24][7] ;
    input n50377;
    output n56165;
    input \rx_data[3] ;
    input n27900;
    output n28964;
    input n22369;
    output n29658;
    output n29659;
    input LED_c;
    input n24633;
    input \data_out_frame[21][0] ;
    output n56162;
    input \data_in_frame[2][0] ;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(41[6:14])
    wire [10:0]t1_10__N_432;
    wire [10:0]t1;   // verilog/neopixel.v(11[12:14])
    
    wire \neo_pixel_transmitter.done_N_516 , n57853, \neo_pixel_transmitter.done , 
        start_N_507, n7, start, n7201, n38255, n61, n67026, n63144, 
        n14, n66759;
    wire [5:0]color_bit_N_502;
    
    wire n66762;
    wire [10:0]n13;
    wire [4:0]bit_ctr_c;   // verilog/neopixel.v(20[11:18])
    
    wire n41, n50325, n56287;
    wire [10:0]n49;
    
    wire n49118, n49117, n59, n49116, n49115, n49114, n27435, 
        n28875, n49113, n49112, n49111, n49110, n49109, n63, n57899, 
        n63156, n56384, n56484, n57623, n57_adj_5683, n43, n32, 
        one_wire_N_499;
    wire [31:0]n149;
    
    wire n20625, n28352;
    wire [1:0]state_1__N_451;
    
    wire n6_adj_5684, n28351, n48543, n48542, n48541, n48540, n48539, 
        n48538, n48537, n48536, n48535, n48534, n66879, n66882, 
        n38340, n50292, n66, n66696, n65381, n66612, n65597, n66822, 
        n63137, n60006, n60007, n60010, n60009, n44, n1, n66693, 
        n66819, n50_adj_5685, n4_adj_5686, n59884, n6_adj_5687, n66609, 
        n56_adj_5688, n25124, n63013, n38251, n63012, n12_adj_5689;
    
    SB_DFF t1_i0 (.Q(t1[0]), .C(clk16MHz), .D(t1_10__N_432[0]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFFE \neo_pixel_transmitter.done_96  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk16MHz), .E(n57853), .D(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFE start_95 (.Q(start), .C(clk16MHz), .E(n7), .D(start_N_507));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 i2203_2_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(n7201));   // verilog/neopixel.v(65[23:32])
    defparam i2203_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22515_2_lut (.I0(state[1]), .I1(t1[0]), .I2(GND_net), .I3(GND_net), 
            .O(n38255));
    defparam i22515_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i47125_4_lut (.I0(n38255), .I1(n61), .I2(t1[10]), .I3(n67026), 
            .O(n63144));   // verilog/neopixel.v(19[11:16])
    defparam i47125_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i44_4_lut (.I0(n63144), .I1(state[1]), .I2(start), .I3(n14), 
            .O(n3173));   // verilog/neopixel.v(19[11:16])
    defparam i44_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 n66759_bdd_4_lut (.I0(n66759), .I1(neopxl_color[21]), .I2(neopxl_color[20]), 
            .I3(color_bit_N_502[1]), .O(n66762));
    defparam n66759_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2201_2_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(color_bit_N_502[1]));   // verilog/neopixel.v(65[23:32])
    defparam i2201_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 timer_10__I_0_inv_0_i1_1_lut (.I0(t0[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[0]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i2_1_lut (.I0(t0[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[1]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i52_3_lut (.I0(bit_ctr_c[2]), .I1(bit_ctr_c[3]), .I2(bit_ctr[1]), 
            .I3(GND_net), .O(n41));
    defparam i52_3_lut.LUT_INIT = 16'h2424;
    SB_LUT4 timer_10__I_0_inv_0_i3_1_lut (.I0(t0[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[2]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut (.I0(n50325), .I1(n41), .I2(bit_ctr[1]), .I3(bit_ctr[0]), 
            .O(n23));
    defparam i3_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i39287_2_lut (.I0(n23), .I1(n38711), .I2(GND_net), .I3(GND_net), 
            .O(n56287));
    defparam i39287_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 timer_2039_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n49118), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2039_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n49117), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_11 (.CI(n49117), .I0(GND_net), .I1(timer[9]), 
            .CO(n49118));
    SB_LUT4 i1_2_lut (.I0(start), .I1(n59), .I2(GND_net), .I3(GND_net), 
            .O(n35156));   // verilog/neopixel.v(19[11:16])
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 timer_2039_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n49116), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_10 (.CI(n49116), .I0(GND_net), .I1(timer[8]), 
            .CO(n49117));
    SB_LUT4 timer_2039_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n49115), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_9 (.CI(n49115), .I0(GND_net), .I1(timer[7]), 
            .CO(n49116));
    SB_LUT4 timer_2039_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n49114), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_8 (.CI(n49114), .I0(GND_net), .I1(timer[6]), 
            .CO(n49115));
    SB_LUT4 timer_10__I_0_inv_0_i4_1_lut (.I0(t0[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[3]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i5_1_lut (.I0(t0[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[4]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut (.I0(n27435), .I1(n35156), .I2(state[1]), .I3(GND_net), 
            .O(n27441));
    defparam i1_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i13030_2_lut (.I0(n27441), .I1(state[1]), .I2(GND_net), .I3(GND_net), 
            .O(n28875));   // verilog/neopixel.v(34[12] 113[6])
    defparam i13030_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 timer_2039_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n49113), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_7 (.CI(n49113), .I0(GND_net), .I1(timer[5]), 
            .CO(n49114));
    SB_LUT4 timer_2039_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n49112), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_6 (.CI(n49112), .I0(GND_net), .I1(timer[4]), 
            .CO(n49113));
    SB_LUT4 timer_2039_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n49111), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_5 (.CI(n49111), .I0(GND_net), .I1(timer[3]), 
            .CO(n49112));
    SB_LUT4 timer_2039_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n49110), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_4 (.CI(n49110), .I0(GND_net), .I1(timer[2]), 
            .CO(n49111));
    SB_LUT4 timer_2039_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n49109), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_3 (.CI(n49109), .I0(GND_net), .I1(timer[1]), 
            .CO(n49110));
    SB_LUT4 timer_2039_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2039_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2039_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n49109));
    SB_LUT4 timer_10__I_0_inv_0_i6_1_lut (.I0(t0[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[5]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i7_1_lut (.I0(t0[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[6]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i8_1_lut (.I0(t0[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[7]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i9_1_lut (.I0(t0[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[8]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i10_1_lut (.I0(t0[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[9]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_10__I_0_inv_0_i11_1_lut (.I0(t0[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n13[10]));   // verilog/neopixel.v(15[9:21])
    defparam timer_10__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_4_lut (.I0(state[1]), .I1(state[0]), .I2(n63), .I3(\neo_pixel_transmitter.done ), 
            .O(n57899));   // verilog/neopixel.v(34[12] 113[6])
    defparam i2_4_lut.LUT_INIT = 16'h0020;
    SB_DFFE bit_ctr_i1 (.Q(bit_ctr[1]), .C(clk16MHz), .E(VCC_net), .D(n29176));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(VCC_net), .D(n5));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 i47043_3_lut (.I0(n63), .I1(state[0]), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n63156));
    defparam i47043_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i2_4_lut_adj_1712 (.I0(n56384), .I1(n56484), .I2(state[0]), 
            .I3(\neo_pixel_transmitter.done ), .O(n57623));
    defparam i2_4_lut_adj_1712.LUT_INIT = 16'hfffe;
    SB_LUT4 i61_4_lut (.I0(n57623), .I1(n63156), .I2(state[1]), .I3(start), 
            .O(n57_adj_5683));
    defparam i61_4_lut.LUT_INIT = 16'hcfc5;
    SB_LUT4 i49477_3_lut (.I0(n43), .I1(n57_adj_5683), .I2(n56484), .I3(GND_net), 
            .O(n32));
    defparam i49477_3_lut.LUT_INIT = 16'h3131;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(one_wire_N_499));   // verilog/neopixel.v(34[12] 113[6])
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_DFF t0_i0_i1 (.Q(t0[1]), .C(clk16MHz), .D(n29155));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF timer_2039__i0 (.Q(timer[0]), .C(clk16MHz), .D(n49[0]));   // verilog/neopixel.v(14[12:21])
    SB_DFF t0_i0_i2 (.Q(t0[2]), .C(clk16MHz), .D(n29154));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i3 (.Q(t0[3]), .C(clk16MHz), .D(n29151));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR bit_ctr_i2 (.Q(bit_ctr_c[2]), .C(clk16MHz), .E(n27441), 
            .D(n149[2]), .R(n28875));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR bit_ctr_i3 (.Q(bit_ctr_c[3]), .C(clk16MHz), .E(n27441), 
            .D(n149[3]), .R(n28875));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR bit_ctr_i4 (.Q(bit_ctr_c[4]), .C(clk16MHz), .E(n27441), 
            .D(n149[4]), .R(n28875));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i4 (.Q(t0[4]), .C(clk16MHz), .D(n29150));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i5 (.Q(t0[5]), .C(clk16MHz), .D(n29149));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i6 (.Q(t0[6]), .C(clk16MHz), .D(n29148));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i7 (.Q(t0[7]), .C(clk16MHz), .D(n29147));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i8 (.Q(t0[8]), .C(clk16MHz), .D(n29146));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i9 (.Q(t0[9]), .C(clk16MHz), .D(n29145));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFF t0_i0_i10 (.Q(t0[10]), .C(clk16MHz), .D(n29144));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR bit_ctr_i0 (.Q(bit_ctr[0]), .C(clk16MHz), .E(n27435), .D(n20625), 
            .R(n28352));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESS state_i0 (.Q(state[0]), .C(clk16MHz), .E(n6_adj_5684), .D(state_1__N_451[0]), 
            .S(n28351));   // verilog/neopixel.v(34[12] 113[6])
    SB_DFFESR one_wire_99 (.Q(NEOPXL_c), .C(clk16MHz), .E(n32), .D(one_wire_N_499), 
            .R(n57899));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 timer_10__I_0_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n13[10]), 
            .I3(n48543), .O(t1_10__N_432[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_10__I_0_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n13[9]), 
            .I3(n48542), .O(t1_10__N_432[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_11 (.CI(n48542), .I0(timer[9]), .I1(n13[9]), 
            .CO(n48543));
    SB_LUT4 timer_10__I_0_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n13[8]), 
            .I3(n48541), .O(t1_10__N_432[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_10 (.CI(n48541), .I0(timer[8]), .I1(n13[8]), 
            .CO(n48542));
    SB_LUT4 timer_10__I_0_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n13[7]), 
            .I3(n48540), .O(t1_10__N_432[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_9 (.CI(n48540), .I0(timer[7]), .I1(n13[7]), 
            .CO(n48541));
    SB_LUT4 timer_10__I_0_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n13[6]), 
            .I3(n48539), .O(t1_10__N_432[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_8 (.CI(n48539), .I0(timer[6]), .I1(n13[6]), 
            .CO(n48540));
    SB_LUT4 timer_10__I_0_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n13[5]), 
            .I3(n48538), .O(t1_10__N_432[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_7 (.CI(n48538), .I0(timer[5]), .I1(n13[5]), 
            .CO(n48539));
    SB_LUT4 timer_10__I_0_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n13[4]), 
            .I3(n48537), .O(t1_10__N_432[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_6 (.CI(n48537), .I0(timer[4]), .I1(n13[4]), 
            .CO(n48538));
    SB_LUT4 timer_10__I_0_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n13[3]), 
            .I3(n48536), .O(t1_10__N_432[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_5 (.CI(n48536), .I0(timer[3]), .I1(n13[3]), 
            .CO(n48537));
    SB_LUT4 timer_10__I_0_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n13[2]), 
            .I3(n48535), .O(t1_10__N_432[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_4 (.CI(n48535), .I0(timer[2]), .I1(n13[2]), 
            .CO(n48536));
    SB_LUT4 timer_10__I_0_add_2_3_lut (.I0(GND_net), .I1(timer[1]), .I2(n13[1]), 
            .I3(n48534), .O(t1_10__N_432[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_3 (.CI(n48534), .I0(timer[1]), .I1(n13[1]), 
            .CO(n48535));
    SB_LUT4 timer_10__I_0_add_2_2_lut (.I0(GND_net), .I1(timer[0]), .I2(n13[0]), 
            .I3(VCC_net), .O(t1_10__N_432[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_10__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_10__I_0_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n13[0]), 
            .CO(n48534));
    SB_DFF t1_i10 (.Q(t1[10]), .C(clk16MHz), .D(t1_10__N_432[10]));   // verilog/neopixel.v(13[8] 16[4])
    SB_LUT4 n66879_bdd_4_lut (.I0(n66879), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(color_bit_N_502[1]), .O(n66882));
    defparam n66879_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF t1_i9 (.Q(t1[9]), .C(clk16MHz), .D(t1_10__N_432[9]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i8 (.Q(t1[8]), .C(clk16MHz), .D(t1_10__N_432[8]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i7 (.Q(t1[7]), .C(clk16MHz), .D(t1_10__N_432[7]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i6 (.Q(t1[6]), .C(clk16MHz), .D(t1_10__N_432[6]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i5 (.Q(t1[5]), .C(clk16MHz), .D(t1_10__N_432[5]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i4 (.Q(t1[4]), .C(clk16MHz), .D(t1_10__N_432[4]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i3 (.Q(t1[3]), .C(clk16MHz), .D(t1_10__N_432[3]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i2 (.Q(t1[2]), .C(clk16MHz), .D(t1_10__N_432[2]));   // verilog/neopixel.v(13[8] 16[4])
    SB_DFF t1_i1 (.Q(t1[1]), .C(clk16MHz), .D(t1_10__N_432[1]));   // verilog/neopixel.v(13[8] 16[4])
    SB_LUT4 i1_2_lut_adj_1713 (.I0(bit_ctr_c[3]), .I1(n38340), .I2(GND_net), 
            .I3(GND_net), .O(n50292));
    defparam i1_2_lut_adj_1713.LUT_INIT = 16'h6666;
    SB_DFF t0_i0_i0 (.Q(t0[0]), .C(clk16MHz), .D(n28939));   // verilog/neopixel.v(34[12] 113[6])
    SB_LUT4 i14_4_lut (.I0(n35156), .I1(n66), .I2(state[1]), .I3(state[0]), 
            .O(n6_adj_5684));
    defparam i14_4_lut.LUT_INIT = 16'hfa3a;
    SB_DFF timer_2039__i1 (.Q(timer[1]), .C(clk16MHz), .D(n49[1]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i2 (.Q(timer[2]), .C(clk16MHz), .D(n49[2]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i3 (.Q(timer[3]), .C(clk16MHz), .D(n49[3]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i4 (.Q(timer[4]), .C(clk16MHz), .D(n49[4]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i5 (.Q(timer[5]), .C(clk16MHz), .D(n49[5]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i6 (.Q(timer[6]), .C(clk16MHz), .D(n49[6]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i7 (.Q(timer[7]), .C(clk16MHz), .D(n49[7]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i8 (.Q(timer[8]), .C(clk16MHz), .D(n49[8]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i9 (.Q(timer[9]), .C(clk16MHz), .D(n49[9]));   // verilog/neopixel.v(14[12:21])
    SB_DFF timer_2039__i10 (.Q(timer[10]), .C(clk16MHz), .D(n49[10]));   // verilog/neopixel.v(14[12:21])
    SB_LUT4 i48319_3_lut (.I0(n66696), .I1(n66882), .I2(color_bit_N_502[2]), 
            .I3(GND_net), .O(n65381));
    defparam i48319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i48535_3_lut (.I0(n65381), .I1(n66612), .I2(n50292), .I3(GND_net), 
            .O(n65597));   // verilog/neopixel.v(24[26:38])
    defparam i48535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46475_4_lut (.I0(n66822), .I1(n50292), .I2(n66762), .I3(color_bit_N_502[2]), 
            .O(n63137));
    defparam i46475_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i22456_4_lut (.I0(n63137), .I1(n56287), .I2(n65597), .I3(n50325), 
            .O(state_1__N_451[0]));   // verilog/neopixel.v(39[18] 44[12])
    defparam i22456_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1_2_lut_adj_1714 (.I0(\data_in_frame[4][2] ), .I1(\data_in_frame[4][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n56059));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1714.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1715 (.I0(\data_in_frame[1][6] ), .I1(\data_in_frame[1][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n55668));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1715.LUT_INIT = 16'h6666;
    SB_LUT4 i42944_3_lut (.I0(neopxl_color[0]), .I1(neopxl_color[1]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n60006));
    defparam i42944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42945_3_lut (.I0(neopxl_color[2]), .I1(neopxl_color[3]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n60007));
    defparam i42945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42948_3_lut (.I0(neopxl_color[6]), .I1(neopxl_color[7]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n60010));
    defparam i42948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42947_3_lut (.I0(neopxl_color[4]), .I1(neopxl_color[5]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n60009));
    defparam i42947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i63_4_lut_4_lut (.I0(t1[3]), .I1(t1[1]), .I2(\neo_pixel_transmitter.done ), 
            .I3(state[0]), .O(n44));
    defparam i63_4_lut_4_lut.LUT_INIT = 16'h1881;
    SB_LUT4 i85_2_lut_3_lut (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(n63), .I3(GND_net), .O(n1));
    defparam i85_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2215_2_lut_3_lut_4_lut (.I0(bit_ctr_c[2]), .I1(bit_ctr[1]), 
            .I2(bit_ctr[0]), .I3(bit_ctr_c[3]), .O(n149[3]));   // verilog/neopixel.v(65[23:32])
    defparam i2215_2_lut_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i60_4_lut_4_lut_4_lut (.I0(t1[3]), .I1(t1[1]), .I2(state[0]), 
            .I3(\neo_pixel_transmitter.done ), .O(n43));
    defparam i60_4_lut_4_lut_4_lut.LUT_INIT = 16'h1880;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[4][2] ), .I1(\data_in_frame[4][3] ), 
            .I2(n56216), .I3(n25933), .O(Kp_23__N_875));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1716 (.I0(\data_out_frame[23][2] ), .I1(\data_out_frame[23][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n55952));
    defparam i1_2_lut_adj_1716.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1717 (.I0(\data_out_frame[24][7] ), .I1(n50377), 
            .I2(GND_net), .I3(GND_net), .O(n56165));
    defparam i1_2_lut_adj_1717.LUT_INIT = 16'h6666;
    SB_LUT4 bit_ctr_0__bdd_4_lut_49656_4_lut_4_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), 
            .I2(neopxl_color[13]), .I3(neopxl_color[12]), .O(n66693));   // verilog/neopixel.v(65[23:32])
    defparam bit_ctr_0__bdd_4_lut_49656_4_lut_4_lut.LUT_INIT = 16'hd5c4;
    SB_LUT4 i13119_3_lut (.I0(\data_in_frame[4][3] ), .I1(\rx_data[3] ), 
            .I2(n27900), .I3(GND_net), .O(n28964));   // verilog/coms.v(130[12] 305[6])
    defparam i13119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i18672_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4][3] ), 
            .I2(n22369), .I3(GND_net), .O(n29658));
    defparam i18672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18678_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4][2] ), 
            .I2(n22369), .I3(GND_net), .O(n29659));
    defparam i18678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 color_bit_N_502_1__bdd_4_lut_4_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), 
            .I2(neopxl_color[17]), .I3(neopxl_color[19]), .O(n66819));
    defparam color_bit_N_502_1__bdd_4_lut_4_lut.LUT_INIT = 16'he6a2;
    SB_LUT4 i2_3_lut_4_lut_adj_1718 (.I0(t1[4]), .I1(t1[0]), .I2(t1[2]), 
            .I3(n50_adj_5685), .O(n56484));
    defparam i2_3_lut_4_lut_adj_1718.LUT_INIT = 16'hffef;
    SB_LUT4 i42831_3_lut_4_lut (.I0(t1[4]), .I1(t1[0]), .I2(t1[10]), .I3(n4_adj_5686), 
            .O(n59884));
    defparam i42831_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut (.I0(n61), .I1(n4_adj_5686), .I2(t1[2]), .I3(GND_net), 
            .O(n6_adj_5687));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_1719 (.I0(n61), .I1(n4_adj_5686), .I2(t1[8]), 
            .I3(t1[10]), .O(n50_adj_5685));
    defparam i2_3_lut_4_lut_adj_1719.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut (.I0(state[0]), .I1(n56287), .I2(LED_c), .I3(state[1]), 
            .O(n27435));   // verilog/neopixel.v(35[4] 112[11])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h80ff;
    SB_LUT4 i12507_2_lut_4_lut (.I0(state[0]), .I1(n56287), .I2(LED_c), 
            .I3(state[1]), .O(n28352));   // verilog/neopixel.v(35[4] 112[11])
    defparam i12507_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i22964_2_lut_3_lut (.I0(bit_ctr_c[3]), .I1(n38340), .I2(bit_ctr_c[4]), 
            .I3(GND_net), .O(n38711));
    defparam i22964_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1720 (.I0(bit_ctr_c[3]), .I1(n38340), .I2(bit_ctr_c[4]), 
            .I3(GND_net), .O(n50325));
    defparam i1_2_lut_3_lut_adj_1720.LUT_INIT = 16'h7878;
    SB_LUT4 i1_2_lut_3_lut_adj_1721 (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr_c[2]), 
            .I3(GND_net), .O(color_bit_N_502[2]));
    defparam i1_2_lut_3_lut_adj_1721.LUT_INIT = 16'h1e1e;
    SB_LUT4 n66819_bdd_4_lut (.I0(n66819), .I1(neopxl_color[18]), .I2(neopxl_color[16]), 
            .I3(bit_ctr[0]), .O(n66822));
    defparam n66819_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i22599_2_lut_3_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr_c[2]), 
            .I3(GND_net), .O(n38340));
    defparam i22599_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 n67023_bdd_4_lut_4_lut_4_lut_4_lut (.I0(t1[3]), .I1(t1[1]), 
            .I2(state[0]), .I3(\neo_pixel_transmitter.done ), .O(n67026));
    defparam n67023_bdd_4_lut_4_lut_4_lut_4_lut.LUT_INIT = 16'h1881;
    SB_LUT4 i2_3_lut_4_lut_adj_1722 (.I0(n24633), .I1(\data_out_frame[23][2] ), 
            .I2(\data_out_frame[23][3] ), .I3(\data_out_frame[21][0] ), 
            .O(n56162));
    defparam i2_3_lut_4_lut_adj_1722.LUT_INIT = 16'h6996;
    SB_LUT4 n66693_bdd_4_lut_4_lut (.I0(color_bit_N_502[1]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(n66693), .O(n66696));   // verilog/neopixel.v(65[23:32])
    defparam n66693_bdd_4_lut_4_lut.LUT_INIT = 16'hf588;
    SB_LUT4 i1_2_lut_3_lut_adj_1723 (.I0(\data_in_frame[2][0] ), .I1(\data_in_frame[1][6] ), 
            .I2(\data_in_frame[1][7] ), .I3(GND_net), .O(n56216));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_adj_1723.LUT_INIT = 16'h9696;
    SB_LUT4 i12_3_lut_4_lut (.I0(start), .I1(n59), .I2(n1), .I3(state[1]), 
            .O(n28351));   // verilog/neopixel.v(34[12] 113[6])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h0f44;
    SB_LUT4 i16_2_lut_3_lut (.I0(start), .I1(n59), .I2(bit_ctr[0]), .I3(GND_net), 
            .O(n20625));   // verilog/neopixel.v(20[11:18])
    defparam i16_2_lut_3_lut.LUT_INIT = 16'hb4b4;
    SB_LUT4 bit_ctr_0__bdd_4_lut_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n66879));
    defparam bit_ctr_0__bdd_4_lut_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 color_bit_N_502_1__bdd_4_lut_49706 (.I0(color_bit_N_502[1]), .I1(n60009), 
            .I2(n60010), .I3(color_bit_N_502[2]), .O(n66609));
    defparam color_bit_N_502_1__bdd_4_lut_49706.LUT_INIT = 16'he4aa;
    SB_LUT4 n66609_bdd_4_lut (.I0(n66609), .I1(n60007), .I2(n60006), .I3(color_bit_N_502[2]), 
            .O(n66612));
    defparam n66609_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_49756_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[22]), 
            .I2(neopxl_color[23]), .I3(bit_ctr[1]), .O(n66759));
    defparam bit_ctr_0__bdd_4_lut_49756_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 i6_3_lut_4_lut (.I0(t1[8]), .I1(t1[5]), .I2(t1[6]), .I3(n56_adj_5688), 
            .O(n14));
    defparam i6_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i2222_3_lut_4_lut (.I0(bit_ctr_c[2]), .I1(n7201), .I2(bit_ctr_c[3]), 
            .I3(bit_ctr_c[4]), .O(n149[4]));   // verilog/neopixel.v(65[23:32])
    defparam i2222_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 i3_4_lut_adj_1724 (.I0(t1[3]), .I1(t1[1]), .I2(t1[4]), .I3(t1[0]), 
            .O(n25124));   // verilog/neopixel.v(60[15:45])
    defparam i3_4_lut_adj_1724.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut (.I0(n25124), .I1(t1[10]), .I2(t1[8]), .I3(n6_adj_5687), 
            .O(n63));
    defparam i4_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_adj_1725 (.I0(t1[2]), .I1(t1[4]), .I2(GND_net), .I3(GND_net), 
            .O(n56_adj_5688));   // verilog/neopixel.v(13[8] 16[4])
    defparam i1_2_lut_adj_1725.LUT_INIT = 16'h2222;
    SB_LUT4 i83_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(n63), .I2(GND_net), 
            .I3(GND_net), .O(n66));
    defparam i83_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i46885_3_lut (.I0(n25124), .I1(n50_adj_5685), .I2(t1[2]), 
            .I3(GND_net), .O(n63013));   // verilog/neopixel.v(19[11:16])
    defparam i46885_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i47730_4_lut (.I0(n56_adj_5688), .I1(n50_adj_5685), .I2(n38251), 
            .I3(t1[0]), .O(n63012));   // verilog/neopixel.v(19[11:16])
    defparam i47730_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i1_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(n63012), .I2(n63013), 
            .I3(state[0]), .O(n59));   // verilog/neopixel.v(19[11:16])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i15_4_lut (.I0(n59), .I1(n1), .I2(state[1]), .I3(start), 
            .O(n7));
    defparam i15_4_lut.LUT_INIT = 16'h3f3a;
    SB_LUT4 i2208_2_lut_3_lut (.I0(bit_ctr_c[2]), .I1(bit_ctr[1]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n149[2]));   // verilog/neopixel.v(65[23:32])
    defparam i2208_2_lut_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i49407_2_lut (.I0(state[1]), .I1(start), .I2(GND_net), .I3(GND_net), 
            .O(start_N_507));   // verilog/neopixel.v(35[4] 112[11])
    defparam i49407_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_1726 (.I0(t1[5]), .I1(t1[6]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_5686));   // verilog/neopixel.v(60[15:45])
    defparam i1_2_lut_adj_1726.LUT_INIT = 16'heeee;
    SB_LUT4 i22511_2_lut (.I0(t1[1]), .I1(t1[3]), .I2(GND_net), .I3(GND_net), 
            .O(n38251));
    defparam i22511_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i39377_2_lut (.I0(t1[3]), .I1(t1[1]), .I2(GND_net), .I3(GND_net), 
            .O(n56384));
    defparam i39377_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1727 (.I0(t1[9]), .I1(t1[7]), .I2(GND_net), .I3(GND_net), 
            .O(n61));
    defparam i1_2_lut_adj_1727.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(t1[2]), .I1(t1[8]), .I2(n44), .I3(n61), .O(n12_adj_5689));
    defparam i5_4_lut.LUT_INIT = 16'h0020;
    SB_LUT4 i2_4_lut_adj_1728 (.I0(state[1]), .I1(n59884), .I2(start), 
            .I3(n12_adj_5689), .O(n57853));
    defparam i2_4_lut_adj_1728.LUT_INIT = 16'hfbfa;
    SB_LUT4 i19392_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[1]), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_516 ));   // verilog/neopixel.v(19[11:16])
    defparam i19392_3_lut.LUT_INIT = 16'hc1c1;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, clk16MHz, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk16MHz;
    input VCC_net;
    output clk32MHz;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(41[6:14])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(41[16:24])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(clk16MHz), .PLLOUTCORE(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=42, LSE_RLINE=46 */ ;   // verilog/TinyFPGA_B.v(42[10] 46[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(0)_U0 
//

module \quadrature_decoder(0)_U0  (ENCODER0_B_N_keep, n1795, ENCODER0_A_N_keep, 
            n1751, GND_net, n1753, n1755, n1757, n1759, n1761, 
            n1763, n1765, n1767, n1769, \encoder0_position[21] , \encoder0_position[20] , 
            \encoder0_position[19] , \encoder0_position[18] , \encoder0_position[17] , 
            \encoder0_position[16] , \encoder0_position[15] , \encoder0_position[14] , 
            \encoder0_position[13] , \encoder0_position[12] , \encoder0_position[11] , 
            \encoder0_position[10] , \encoder0_position[9] , \encoder0_position[8] , 
            \encoder0_position[7] , \encoder0_position[6] , \encoder0_position[5] , 
            \encoder0_position[4] , \encoder0_position[3] , \encoder0_position[2] , 
            \encoder0_position[1] , \encoder0_position[0] , VCC_net, \a_new[1] , 
            \b_new[1] , b_prev, n29063, n1749, n29062, a_prev, n29060, 
            position_31__N_3836, debounce_cnt_N_3833) /* synthesis lattice_noprune=1 */ ;
    input ENCODER0_B_N_keep;
    input n1795;
    input ENCODER0_A_N_keep;
    output n1751;
    input GND_net;
    output n1753;
    output n1755;
    output n1757;
    output n1759;
    output n1761;
    output n1763;
    output n1765;
    output n1767;
    output n1769;
    output \encoder0_position[21] ;
    output \encoder0_position[20] ;
    output \encoder0_position[19] ;
    output \encoder0_position[18] ;
    output \encoder0_position[17] ;
    output \encoder0_position[16] ;
    output \encoder0_position[15] ;
    output \encoder0_position[14] ;
    output \encoder0_position[13] ;
    output \encoder0_position[12] ;
    output \encoder0_position[11] ;
    output \encoder0_position[10] ;
    output \encoder0_position[9] ;
    output \encoder0_position[8] ;
    output \encoder0_position[7] ;
    output \encoder0_position[6] ;
    output \encoder0_position[5] ;
    output \encoder0_position[4] ;
    output \encoder0_position[3] ;
    output \encoder0_position[2] ;
    output \encoder0_position[1] ;
    output \encoder0_position[0] ;
    input VCC_net;
    output \a_new[1] ;
    output \b_new[1] ;
    output b_prev;
    input n29063;
    output n1749;
    input n29062;
    output a_prev;
    input n29060;
    output position_31__N_3836;
    output debounce_cnt_N_3833;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    wire [31:0]n133;
    
    wire direction_N_3840, n49274, n49273, n49272, n49271, n49270, 
        n49269, n49268, n49267, n49266, n49265, n49264, n49263, 
        n49262, n49261, n49260, n49259, n49258, n49257, n49256, 
        n49255, n49254, n49253, n49252, n49251, n49250, n49249, 
        n49248, n49247, n49246, n49245, n49244;
    
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1795), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1795), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 position_2054_add_4_33_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1751), .I3(n49274), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2054_add_4_32_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1753), .I3(n49273), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_32 (.CI(n49273), .I0(direction_N_3840), 
            .I1(n1753), .CO(n49274));
    SB_LUT4 position_2054_add_4_31_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1755), .I3(n49272), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_31 (.CI(n49272), .I0(direction_N_3840), 
            .I1(n1755), .CO(n49273));
    SB_LUT4 position_2054_add_4_30_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1757), .I3(n49271), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_30 (.CI(n49271), .I0(direction_N_3840), 
            .I1(n1757), .CO(n49272));
    SB_LUT4 position_2054_add_4_29_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1759), .I3(n49270), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_29 (.CI(n49270), .I0(direction_N_3840), 
            .I1(n1759), .CO(n49271));
    SB_LUT4 position_2054_add_4_28_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1761), .I3(n49269), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_28 (.CI(n49269), .I0(direction_N_3840), 
            .I1(n1761), .CO(n49270));
    SB_LUT4 position_2054_add_4_27_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1763), .I3(n49268), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_27 (.CI(n49268), .I0(direction_N_3840), 
            .I1(n1763), .CO(n49269));
    SB_LUT4 position_2054_add_4_26_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1765), .I3(n49267), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_26 (.CI(n49267), .I0(direction_N_3840), 
            .I1(n1765), .CO(n49268));
    SB_LUT4 position_2054_add_4_25_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1767), .I3(n49266), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_25 (.CI(n49266), .I0(direction_N_3840), 
            .I1(n1767), .CO(n49267));
    SB_LUT4 position_2054_add_4_24_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(n1769), .I3(n49265), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_24 (.CI(n49265), .I0(direction_N_3840), 
            .I1(n1769), .CO(n49266));
    SB_LUT4 position_2054_add_4_23_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[21] ), .I3(n49264), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_23 (.CI(n49264), .I0(direction_N_3840), 
            .I1(\encoder0_position[21] ), .CO(n49265));
    SB_LUT4 position_2054_add_4_22_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[20] ), .I3(n49263), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_22 (.CI(n49263), .I0(direction_N_3840), 
            .I1(\encoder0_position[20] ), .CO(n49264));
    SB_LUT4 position_2054_add_4_21_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[19] ), .I3(n49262), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_21 (.CI(n49262), .I0(direction_N_3840), 
            .I1(\encoder0_position[19] ), .CO(n49263));
    SB_LUT4 position_2054_add_4_20_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[18] ), .I3(n49261), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_20 (.CI(n49261), .I0(direction_N_3840), 
            .I1(\encoder0_position[18] ), .CO(n49262));
    SB_LUT4 position_2054_add_4_19_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[17] ), .I3(n49260), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_19 (.CI(n49260), .I0(direction_N_3840), 
            .I1(\encoder0_position[17] ), .CO(n49261));
    SB_LUT4 position_2054_add_4_18_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[16] ), .I3(n49259), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_18 (.CI(n49259), .I0(direction_N_3840), 
            .I1(\encoder0_position[16] ), .CO(n49260));
    SB_LUT4 position_2054_add_4_17_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[15] ), .I3(n49258), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_17 (.CI(n49258), .I0(direction_N_3840), 
            .I1(\encoder0_position[15] ), .CO(n49259));
    SB_LUT4 position_2054_add_4_16_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[14] ), .I3(n49257), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_16 (.CI(n49257), .I0(direction_N_3840), 
            .I1(\encoder0_position[14] ), .CO(n49258));
    SB_LUT4 position_2054_add_4_15_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[13] ), .I3(n49256), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_15 (.CI(n49256), .I0(direction_N_3840), 
            .I1(\encoder0_position[13] ), .CO(n49257));
    SB_LUT4 position_2054_add_4_14_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[12] ), .I3(n49255), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_14 (.CI(n49255), .I0(direction_N_3840), 
            .I1(\encoder0_position[12] ), .CO(n49256));
    SB_LUT4 position_2054_add_4_13_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[11] ), .I3(n49254), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_13 (.CI(n49254), .I0(direction_N_3840), 
            .I1(\encoder0_position[11] ), .CO(n49255));
    SB_LUT4 position_2054_add_4_12_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[10] ), .I3(n49253), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_12 (.CI(n49253), .I0(direction_N_3840), 
            .I1(\encoder0_position[10] ), .CO(n49254));
    SB_LUT4 position_2054_add_4_11_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[9] ), .I3(n49252), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_11 (.CI(n49252), .I0(direction_N_3840), 
            .I1(\encoder0_position[9] ), .CO(n49253));
    SB_LUT4 position_2054_add_4_10_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[8] ), .I3(n49251), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_10 (.CI(n49251), .I0(direction_N_3840), 
            .I1(\encoder0_position[8] ), .CO(n49252));
    SB_LUT4 position_2054_add_4_9_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[7] ), .I3(n49250), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_9 (.CI(n49250), .I0(direction_N_3840), 
            .I1(\encoder0_position[7] ), .CO(n49251));
    SB_LUT4 position_2054_add_4_8_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[6] ), .I3(n49249), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_8 (.CI(n49249), .I0(direction_N_3840), 
            .I1(\encoder0_position[6] ), .CO(n49250));
    SB_LUT4 position_2054_add_4_7_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[5] ), .I3(n49248), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_7 (.CI(n49248), .I0(direction_N_3840), 
            .I1(\encoder0_position[5] ), .CO(n49249));
    SB_LUT4 position_2054_add_4_6_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[4] ), .I3(n49247), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_6 (.CI(n49247), .I0(direction_N_3840), 
            .I1(\encoder0_position[4] ), .CO(n49248));
    SB_LUT4 position_2054_add_4_5_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[3] ), .I3(n49246), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_5 (.CI(n49246), .I0(direction_N_3840), 
            .I1(\encoder0_position[3] ), .CO(n49247));
    SB_LUT4 position_2054_add_4_4_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[2] ), .I3(n49245), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_4 (.CI(n49245), .I0(direction_N_3840), 
            .I1(\encoder0_position[2] ), .CO(n49246));
    SB_LUT4 position_2054_add_4_3_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(\encoder0_position[1] ), .I3(n49244), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_3 (.CI(n49244), .I0(direction_N_3840), 
            .I1(\encoder0_position[1] ), .CO(n49245));
    SB_LUT4 position_2054_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\encoder0_position[0] ), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2054_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2054_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\encoder0_position[0] ), 
            .CO(n49244));
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1795), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(\b_new[1] ), .C(n1795), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 b_prev_I_0_48_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3840));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_48_2_lut.LUT_INIT = 16'h9999;
    SB_DFF direction_42 (.Q(n1749), .C(n1795), .D(n29063));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_prev_40 (.Q(a_prev), .C(n1795), .D(n29062));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_prev_41 (.Q(b_prev), .C(n1795), .D(n29060));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_2054__i0 (.Q(\encoder0_position[0] ), .C(n1795), .E(position_31__N_3836), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i1 (.Q(\encoder0_position[1] ), .C(n1795), .E(position_31__N_3836), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i2 (.Q(\encoder0_position[2] ), .C(n1795), .E(position_31__N_3836), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i3 (.Q(\encoder0_position[3] ), .C(n1795), .E(position_31__N_3836), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i4 (.Q(\encoder0_position[4] ), .C(n1795), .E(position_31__N_3836), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i5 (.Q(\encoder0_position[5] ), .C(n1795), .E(position_31__N_3836), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i6 (.Q(\encoder0_position[6] ), .C(n1795), .E(position_31__N_3836), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i7 (.Q(\encoder0_position[7] ), .C(n1795), .E(position_31__N_3836), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i8 (.Q(\encoder0_position[8] ), .C(n1795), .E(position_31__N_3836), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i9 (.Q(\encoder0_position[9] ), .C(n1795), .E(position_31__N_3836), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i10 (.Q(\encoder0_position[10] ), .C(n1795), 
            .E(position_31__N_3836), .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i11 (.Q(\encoder0_position[11] ), .C(n1795), 
            .E(position_31__N_3836), .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i12 (.Q(\encoder0_position[12] ), .C(n1795), 
            .E(position_31__N_3836), .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i13 (.Q(\encoder0_position[13] ), .C(n1795), 
            .E(position_31__N_3836), .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i14 (.Q(\encoder0_position[14] ), .C(n1795), 
            .E(position_31__N_3836), .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i15 (.Q(\encoder0_position[15] ), .C(n1795), 
            .E(position_31__N_3836), .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i16 (.Q(\encoder0_position[16] ), .C(n1795), 
            .E(position_31__N_3836), .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i17 (.Q(\encoder0_position[17] ), .C(n1795), 
            .E(position_31__N_3836), .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i18 (.Q(\encoder0_position[18] ), .C(n1795), 
            .E(position_31__N_3836), .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i19 (.Q(\encoder0_position[19] ), .C(n1795), 
            .E(position_31__N_3836), .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i20 (.Q(\encoder0_position[20] ), .C(n1795), 
            .E(position_31__N_3836), .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i21 (.Q(\encoder0_position[21] ), .C(n1795), 
            .E(position_31__N_3836), .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i22 (.Q(n1769), .C(n1795), .E(position_31__N_3836), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i23 (.Q(n1767), .C(n1795), .E(position_31__N_3836), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i24 (.Q(n1765), .C(n1795), .E(position_31__N_3836), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i25 (.Q(n1763), .C(n1795), .E(position_31__N_3836), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i26 (.Q(n1761), .C(n1795), .E(position_31__N_3836), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i27 (.Q(n1759), .C(n1795), .E(position_31__N_3836), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i28 (.Q(n1757), .C(n1795), .E(position_31__N_3836), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i29 (.Q(n1755), .C(n1795), .E(position_31__N_3836), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i30 (.Q(n1753), .C(n1795), .E(position_31__N_3836), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2054__i31 (.Q(n1751), .C(n1795), .E(position_31__N_3836), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 debounce_cnt_I_936_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(debounce_cnt_N_3833));   // vhdl/quadrature_decoder.vhd(53[8:58])
    defparam debounce_cnt_I_936_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 position_31__I_937_4_lut (.I0(a_prev), .I1(b_prev), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(position_31__N_3836));   // vhdl/quadrature_decoder.vhd(63[11:57])
    defparam position_31__I_937_4_lut.LUT_INIT = 16'h7bde;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (state_7__N_4319, GND_net, clk16MHz, CS_c, CS_CLK_c, 
            VCC_net, n27290, \current[15] , n29106, \current[1] , 
            n29105, \current[2] , n29104, \current[3] , n29103, \current[4] , 
            n29102, \current[5] , n29101, \current[6] , n29100, \current[7] , 
            n29099, \current[8] , n29098, \current[9] , n29097, \current[10] , 
            n29096, \current[11] , n29826, \data[15] , n29825, \data[12] , 
            n29824, \data[11] , n29823, \data[10] , n29822, \data[9] , 
            n29821, \data[8] , n29820, \data[7] , n29819, \data[6] , 
            n29818, \data[5] , n29817, \data[4] , n29816, \data[3] , 
            n29815, \data[2] , n29814, \data[1] , n29600, \data[0] , 
            n28927, \current[0] , n5, n11, n25130, n25133, n5_adj_21, 
            n5_adj_22, n38316, n25141, n25110) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output state_7__N_4319;
    input GND_net;
    input clk16MHz;
    output CS_c;
    output CS_CLK_c;
    input VCC_net;
    output n27290;
    output \current[15] ;
    input n29106;
    output \current[1] ;
    input n29105;
    output \current[2] ;
    input n29104;
    output \current[3] ;
    input n29103;
    output \current[4] ;
    input n29102;
    output \current[5] ;
    input n29101;
    output \current[6] ;
    input n29100;
    output \current[7] ;
    input n29099;
    output \current[8] ;
    input n29098;
    output \current[9] ;
    input n29097;
    output \current[10] ;
    input n29096;
    output \current[11] ;
    input n29826;
    output \data[15] ;
    input n29825;
    output \data[12] ;
    input n29824;
    output \data[11] ;
    input n29823;
    output \data[10] ;
    input n29822;
    output \data[9] ;
    input n29821;
    output \data[8] ;
    input n29820;
    output \data[7] ;
    input n29819;
    output \data[6] ;
    input n29818;
    output \data[5] ;
    input n29817;
    output \data[4] ;
    input n29816;
    output \data[3] ;
    input n29815;
    output \data[2] ;
    input n29814;
    output \data[1] ;
    input n29600;
    output \data[0] ;
    input n28927;
    output \current[0] ;
    output n5;
    output n11;
    output n25130;
    output n25133;
    output n5_adj_21;
    output n5_adj_22;
    output n38316;
    output n25141;
    output n25110;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(41[6:14])
    wire [7:0]state;   // verilog/tli4970.v(29[13:18])
    
    wire n27421, clk_slow_N_4232, clk_out;
    wire [2:0]n17;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire n49236, n49235;
    wire [11:0]n53;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire n49234, n49233, n49232, n49231, n49230, n49229, n49228, 
        n49227, n49226, n49225, n49224;
    wire [7:0]n37;
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    
    wire n49210, n49209, n49208, n49207, n63059, n49206, n2, n63063, 
        n49205, n63064, n49204, n63044;
    wire [13:0]n241;
    
    wire n28888, n22219, delay_counter_15__N_4314, clk_slow_N_4233, 
        n38650, n27371, n28359, n9, n11039, n22223, n28929, n22225, 
        n22227, n6, n15, n8, n12, n10;
    
    SB_LUT4 state_7__I_0_77_i9_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(state_7__N_4319));   // verilog/tli4970.v(53[7:17])
    defparam state_7__I_0_77_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i11655_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n27421));
    defparam i11655_2_lut.LUT_INIT = 16'h6666;
    SB_DFF clk_slow_63 (.Q(clk_slow), .C(clk16MHz), .D(clk_slow_N_4232));   // verilog/tli4970.v(13[10] 19[6])
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 counter_2050_2051_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n49236), .O(n17[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2050_2051_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2050_2051_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n49235), .O(n17[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2050_2051_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2050_2051_add_4_3 (.CI(n49235), .I0(GND_net), .I1(counter[1]), 
            .CO(n49236));
    SB_LUT4 counter_2050_2051_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n17[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2050_2051_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2050_2051_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n49235));
    SB_LUT4 delay_counter_2048_2049_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n49234), .O(n53[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_2048_2049_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n49233), .O(n53[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_12 (.CI(n49233), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n49234));
    SB_LUT4 delay_counter_2048_2049_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n49232), .O(n53[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_11 (.CI(n49232), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n49233));
    SB_LUT4 delay_counter_2048_2049_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n49231), .O(n53[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_10 (.CI(n49231), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n49232));
    SB_LUT4 delay_counter_2048_2049_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n49230), .O(n53[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_9 (.CI(n49230), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n49231));
    SB_LUT4 delay_counter_2048_2049_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n49229), .O(n53[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_8 (.CI(n49229), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n49230));
    SB_LUT4 delay_counter_2048_2049_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n49228), .O(n53[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_7 (.CI(n49228), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n49229));
    SB_LUT4 delay_counter_2048_2049_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n49227), .O(n53[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_6 (.CI(n49227), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n49228));
    SB_LUT4 delay_counter_2048_2049_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n49226), .O(n53[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_5 (.CI(n49226), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n49227));
    SB_LUT4 delay_counter_2048_2049_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n49225), .O(n53[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_4 (.CI(n49225), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n49226));
    SB_LUT4 delay_counter_2048_2049_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n49224), .O(n53[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_3 (.CI(n49224), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n49225));
    SB_LUT4 delay_counter_2048_2049_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n53[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2048_2049_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2048_2049_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n49224));
    SB_LUT4 bit_counter_2044_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n49210), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_2044_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n49209), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2044_add_4_8 (.CI(n49209), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n49210));
    SB_LUT4 bit_counter_2044_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n49208), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2044_add_4_7 (.CI(n49208), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n49209));
    SB_LUT4 bit_counter_2044_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n49207), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2044_add_4_6 (.CI(n49207), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n49208));
    SB_LUT4 bit_counter_2044_add_4_5_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n49206), .O(n63059)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_5 (.CI(n49206), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n49207));
    SB_LUT4 bit_counter_2044_add_4_4_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n49205), .O(n63063)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_4 (.CI(n49205), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n49206));
    SB_LUT4 bit_counter_2044_add_4_3_lut (.I0(n2), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n49204), .O(n63064)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_3 (.CI(n49204), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n49205));
    SB_LUT4 bit_counter_2044_add_4_2_lut (.I0(n2), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n63044)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2044_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2044_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n49204));
    SB_LUT4 i2521_1_lut (.I0(state[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2));
    defparam i2521_1_lut.LUT_INIT = 16'h5555;
    SB_DFFNE current__i13 (.Q(\current[15] ), .C(clk_slow), .E(n27290), 
            .D(n241[13]));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNESR bit_counter_2044__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n27421), 
            .D(n37[7]), .R(n28888));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2044__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n27421), 
            .D(n37[6]), .R(n28888));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2044__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n27421), 
            .D(n37[5]), .R(n28888));   // verilog/tli4970.v(55[24:39])
    SB_DFFNESR bit_counter_2044__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n27421), 
            .D(n37[4]), .R(n28888));   // verilog/tli4970.v(55[24:39])
    SB_DFFN current__i2 (.Q(\current[1] ), .C(clk_slow), .D(n29106));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i3 (.Q(\current[2] ), .C(clk_slow), .D(n29105));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i4 (.Q(\current[3] ), .C(clk_slow), .D(n29104));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i5 (.Q(\current[4] ), .C(clk_slow), .D(n29103));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i6 (.Q(\current[5] ), .C(clk_slow), .D(n29102));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i7 (.Q(\current[6] ), .C(clk_slow), .D(n29101));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i8 (.Q(\current[7] ), .C(clk_slow), .D(n29100));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i9 (.Q(\current[8] ), .C(clk_slow), .D(n29099));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i10 (.Q(\current[9] ), .C(clk_slow), .D(n29098));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i11 (.Q(\current[10] ), .C(clk_slow), .D(n29097));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i12 (.Q(\current[11] ), .C(clk_slow), .D(n29096));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_2044__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n27421), 
            .D(n22219));   // verilog/tli4970.v(55[24:39])
    SB_DFFNSR delay_counter_2048_2049__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n53[0]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_2050_2051__i1 (.Q(counter[0]), .C(clk16MHz), .D(n17[0]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_DFFNESS state_i0 (.Q(state[0]), .C(clk_slow), .E(n27371), .D(n38650), 
            .S(n28359));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n29826));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n29825));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n29824));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n29823));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n29822));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n29821));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n29820));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n29819));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n29818));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n29817));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n29816));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n29815));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n29814));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n29600));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN clk_out_67 (.Q(clk_out), .C(clk_slow), .D(n9));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNESR state_i1 (.Q(state[1]), .C(clk_slow), .E(n27371), .D(n11039), 
            .R(n28359));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_2044__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n27421), 
            .D(n22223));   // verilog/tli4970.v(55[24:39])
    SB_DFFN slave_select_66 (.Q(CS_c), .C(clk_slow), .D(n28929));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFN current__i1 (.Q(\current[0] ), .C(clk_slow), .D(n28927));   // verilog/tli4970.v(35[10] 68[6])
    SB_DFFNE bit_counter_2044__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n27421), 
            .D(n22225));   // verilog/tli4970.v(55[24:39])
    SB_DFFNE bit_counter_2044__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n27421), 
            .D(n22227));   // verilog/tli4970.v(55[24:39])
    SB_DFFNSR delay_counter_2048_2049__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n53[1]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n53[2]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n53[3]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n53[4]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n53[5]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n53[6]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n53[7]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n53[8]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n53[9]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n53[10]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFNSR delay_counter_2048_2049__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n53[11]), .R(delay_counter_15__N_4314));   // verilog/tli4970.v(40[24:39])
    SB_DFFSR counter_2050_2051__i2 (.Q(counter[1]), .C(clk16MHz), .D(n17[1]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2050_2051__i3 (.Q(counter[2]), .C(clk16MHz), .D(n17[2]), 
            .R(clk_slow_N_4233));   // verilog/tli4970.v(14[16:27])
    SB_LUT4 equal_330_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(54[9:26])
    defparam equal_330_i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut (.I0(bit_counter[5]), .I1(bit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6));   // verilog/tli4970.v(56[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(bit_counter[6]), .I1(bit_counter[7]), .I2(n11), 
            .I3(n6), .O(n15));   // verilog/tli4970.v(56[12:26])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i49256_2_lut (.I0(n15), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n38650));
    defparam i49256_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i2179_3_lut (.I0(counter[0]), .I1(counter[2]), .I2(counter[1]), 
            .I3(GND_net), .O(clk_slow_N_4233));
    defparam i2179_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 clk_slow_I_0_72_2_lut (.I0(clk_slow), .I1(clk_slow_N_4233), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4232));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_72_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49242_3_lut (.I0(\data[15] ), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n27290));
    defparam i49242_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i2243_1_lut (.I0(\data[12] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n241[13]));
    defparam i2243_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6638_3_lut (.I0(state[0]), .I1(n63059), .I2(state[1]), .I3(GND_net), 
            .O(n22227));   // verilog/tli4970.v(55[24:39])
    defparam i6638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6636_3_lut (.I0(state[0]), .I1(n63063), .I2(state[1]), .I3(GND_net), 
            .O(n22225));   // verilog/tli4970.v(55[24:39])
    defparam i6636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6634_3_lut (.I0(state[0]), .I1(n63064), .I2(state[1]), .I3(GND_net), 
            .O(n22223));   // verilog/tli4970.v(55[24:39])
    defparam i6634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2153_i2_3_lut (.I0(n15), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n11039));
    defparam mux_2153_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(bit_counter[3]), 
            .I3(bit_counter[2]), .O(n25130));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1709 (.I0(state[0]), .I1(state[1]), 
            .I2(bit_counter[3]), .I3(bit_counter[2]), .O(n25133));   // verilog/tli4970.v(43[5] 67[12])
    defparam i1_2_lut_3_lut_4_lut_adj_1709.LUT_INIT = 16'hffbf;
    SB_LUT4 i3_3_lut (.I0(delay_counter[1]), .I1(delay_counter[2]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2180_4_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(n8), 
            .I3(delay_counter[0]), .O(n12));
    defparam i2180_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i4_4_lut_adj_1710 (.I0(delay_counter[11]), .I1(delay_counter[7]), 
            .I2(delay_counter[8]), .I3(delay_counter[9]), .O(n10));
    defparam i4_4_lut_adj_1710.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut (.I0(delay_counter[10]), .I1(n10), .I2(n12), .I3(delay_counter[6]), 
            .O(delay_counter_15__N_4314));
    defparam i5_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 i6631_3_lut (.I0(state[0]), .I1(n63044), .I2(state[1]), .I3(GND_net), 
            .O(n22219));   // verilog/tli4970.v(55[24:39])
    defparam i6631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_337_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_21));   // verilog/tli4970.v(54[9:26])
    defparam equal_337_i5_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_328_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_22));   // verilog/tli4970.v(54[9:26])
    defparam equal_328_i5_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i22576_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n38316));
    defparam i22576_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(state[0]), 
            .I3(state[1]), .O(n25141));   // verilog/tli4970.v(43[5] 67[12])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i13084_3_lut_3_lut (.I0(state[0]), .I1(state[1]), .I2(CS_c), 
            .I3(GND_net), .O(n28929));
    defparam i13084_3_lut_3_lut.LUT_INIT = 16'hd1d1;
    SB_LUT4 i49470_4_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(clk_out), 
            .I3(n15), .O(n9));
    defparam i49470_4_lut_4_lut.LUT_INIT = 16'hf2b2;
    SB_LUT4 i1_2_lut_4_lut (.I0(delay_counter_15__N_4314), .I1(state[0]), 
            .I2(state[1]), .I3(n15), .O(n27371));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'heefe;
    SB_LUT4 i12514_2_lut_4_lut (.I0(delay_counter_15__N_4314), .I1(state[0]), 
            .I2(state[1]), .I3(n15), .O(n28359));   // verilog/tli4970.v(35[10] 68[6])
    defparam i12514_2_lut_4_lut.LUT_INIT = 16'h2202;
    SB_LUT4 equal_268_i11_2_lut_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(bit_counter[0]), .I3(bit_counter[1]), .O(n11));   // verilog/tli4970.v(54[9:26])
    defparam equal_268_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1711 (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(state[0]), .I3(state[1]), .O(n25110));   // verilog/tli4970.v(54[9:26])
    defparam i1_2_lut_3_lut_4_lut_adj_1711.LUT_INIT = 16'hfeff;
    SB_LUT4 i13043_2_lut_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n28888));   // verilog/tli4970.v(55[24:39])
    defparam i13043_2_lut_2_lut.LUT_INIT = 16'h4444;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(0) 
//

module \quadrature_decoder(0)  (ENCODER1_B_N_keep, n1795, ENCODER1_A_N_keep, 
            b_prev, \a_new[1] , GND_net, encoder1_position, VCC_net, 
            \b_new[1] , n29064, a_prev, position_31__N_3836, n28938, 
            n28937, n1800, debounce_cnt_N_3833) /* synthesis lattice_noprune=1 */ ;
    input ENCODER1_B_N_keep;
    input n1795;
    input ENCODER1_A_N_keep;
    output b_prev;
    output \a_new[1] ;
    input GND_net;
    output [31:0]encoder1_position;
    input VCC_net;
    output \b_new[1] ;
    input n29064;
    output a_prev;
    output position_31__N_3836;
    input n28938;
    input n28937;
    output n1800;
    output debounce_cnt_N_3833;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(39[9:14])
    
    wire direction_N_3840;
    wire [31:0]n133;
    
    wire n49172, n49171, n49170, n49169, n49168, n49167, n49166, 
        n49165, n49164, n49163, n49162, n49161, n49160, n49159, 
        n49158, n49157, n49156, n49155, n49154, n49153, n49152, 
        n49151, n49150, n49149, n49148, n49147, n49146, n49145, 
        n49144, n49143, n49142;
    
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1795), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1795), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_LUT4 b_prev_I_0_48_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3840));   // vhdl/quadrature_decoder.vhd(64[18:37])
    defparam b_prev_I_0_48_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 position_2041_add_4_33_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[31]), .I3(n49172), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2041_add_4_32_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[30]), .I3(n49171), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_32 (.CI(n49171), .I0(direction_N_3840), 
            .I1(encoder1_position[30]), .CO(n49172));
    SB_LUT4 position_2041_add_4_31_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[29]), .I3(n49170), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_31 (.CI(n49170), .I0(direction_N_3840), 
            .I1(encoder1_position[29]), .CO(n49171));
    SB_LUT4 position_2041_add_4_30_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[28]), .I3(n49169), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_30 (.CI(n49169), .I0(direction_N_3840), 
            .I1(encoder1_position[28]), .CO(n49170));
    SB_LUT4 position_2041_add_4_29_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[27]), .I3(n49168), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_29 (.CI(n49168), .I0(direction_N_3840), 
            .I1(encoder1_position[27]), .CO(n49169));
    SB_LUT4 position_2041_add_4_28_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[26]), .I3(n49167), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_28 (.CI(n49167), .I0(direction_N_3840), 
            .I1(encoder1_position[26]), .CO(n49168));
    SB_LUT4 position_2041_add_4_27_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[25]), .I3(n49166), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_27 (.CI(n49166), .I0(direction_N_3840), 
            .I1(encoder1_position[25]), .CO(n49167));
    SB_LUT4 position_2041_add_4_26_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[24]), .I3(n49165), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_26 (.CI(n49165), .I0(direction_N_3840), 
            .I1(encoder1_position[24]), .CO(n49166));
    SB_LUT4 position_2041_add_4_25_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[23]), .I3(n49164), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_25 (.CI(n49164), .I0(direction_N_3840), 
            .I1(encoder1_position[23]), .CO(n49165));
    SB_LUT4 position_2041_add_4_24_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[22]), .I3(n49163), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_24 (.CI(n49163), .I0(direction_N_3840), 
            .I1(encoder1_position[22]), .CO(n49164));
    SB_LUT4 position_2041_add_4_23_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[21]), .I3(n49162), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_23 (.CI(n49162), .I0(direction_N_3840), 
            .I1(encoder1_position[21]), .CO(n49163));
    SB_LUT4 position_2041_add_4_22_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[20]), .I3(n49161), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_22 (.CI(n49161), .I0(direction_N_3840), 
            .I1(encoder1_position[20]), .CO(n49162));
    SB_LUT4 position_2041_add_4_21_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[19]), .I3(n49160), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_21 (.CI(n49160), .I0(direction_N_3840), 
            .I1(encoder1_position[19]), .CO(n49161));
    SB_LUT4 position_2041_add_4_20_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[18]), .I3(n49159), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_20 (.CI(n49159), .I0(direction_N_3840), 
            .I1(encoder1_position[18]), .CO(n49160));
    SB_LUT4 position_2041_add_4_19_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[17]), .I3(n49158), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_19 (.CI(n49158), .I0(direction_N_3840), 
            .I1(encoder1_position[17]), .CO(n49159));
    SB_LUT4 position_2041_add_4_18_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[16]), .I3(n49157), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_18 (.CI(n49157), .I0(direction_N_3840), 
            .I1(encoder1_position[16]), .CO(n49158));
    SB_LUT4 position_2041_add_4_17_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[15]), .I3(n49156), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_17 (.CI(n49156), .I0(direction_N_3840), 
            .I1(encoder1_position[15]), .CO(n49157));
    SB_LUT4 position_2041_add_4_16_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[14]), .I3(n49155), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_16 (.CI(n49155), .I0(direction_N_3840), 
            .I1(encoder1_position[14]), .CO(n49156));
    SB_LUT4 position_2041_add_4_15_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[13]), .I3(n49154), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_15 (.CI(n49154), .I0(direction_N_3840), 
            .I1(encoder1_position[13]), .CO(n49155));
    SB_LUT4 position_2041_add_4_14_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[12]), .I3(n49153), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_14 (.CI(n49153), .I0(direction_N_3840), 
            .I1(encoder1_position[12]), .CO(n49154));
    SB_LUT4 position_2041_add_4_13_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[11]), .I3(n49152), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_13 (.CI(n49152), .I0(direction_N_3840), 
            .I1(encoder1_position[11]), .CO(n49153));
    SB_LUT4 position_2041_add_4_12_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[10]), .I3(n49151), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_12 (.CI(n49151), .I0(direction_N_3840), 
            .I1(encoder1_position[10]), .CO(n49152));
    SB_LUT4 position_2041_add_4_11_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[9]), .I3(n49150), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_11 (.CI(n49150), .I0(direction_N_3840), 
            .I1(encoder1_position[9]), .CO(n49151));
    SB_LUT4 position_2041_add_4_10_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[8]), .I3(n49149), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_10 (.CI(n49149), .I0(direction_N_3840), 
            .I1(encoder1_position[8]), .CO(n49150));
    SB_LUT4 position_2041_add_4_9_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[7]), .I3(n49148), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_9 (.CI(n49148), .I0(direction_N_3840), 
            .I1(encoder1_position[7]), .CO(n49149));
    SB_LUT4 position_2041_add_4_8_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[6]), .I3(n49147), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_8 (.CI(n49147), .I0(direction_N_3840), 
            .I1(encoder1_position[6]), .CO(n49148));
    SB_LUT4 position_2041_add_4_7_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[5]), .I3(n49146), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_7 (.CI(n49146), .I0(direction_N_3840), 
            .I1(encoder1_position[5]), .CO(n49147));
    SB_LUT4 position_2041_add_4_6_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[4]), .I3(n49145), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_6 (.CI(n49145), .I0(direction_N_3840), 
            .I1(encoder1_position[4]), .CO(n49146));
    SB_LUT4 position_2041_add_4_5_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[3]), .I3(n49144), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_5 (.CI(n49144), .I0(direction_N_3840), 
            .I1(encoder1_position[3]), .CO(n49145));
    SB_LUT4 position_2041_add_4_4_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[2]), .I3(n49143), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_4 (.CI(n49143), .I0(direction_N_3840), 
            .I1(encoder1_position[2]), .CO(n49144));
    SB_LUT4 position_2041_add_4_3_lut (.I0(GND_net), .I1(direction_N_3840), 
            .I2(encoder1_position[1]), .I3(n49142), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_3 (.CI(n49142), .I0(direction_N_3840), 
            .I1(encoder1_position[1]), .CO(n49143));
    SB_LUT4 position_2041_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder1_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2041_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2041_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder1_position[0]), 
            .CO(n49142));
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1795), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF b_new_i1 (.Q(\b_new[1] ), .C(n1795), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF a_prev_40 (.Q(a_prev), .C(n1795), .D(n29064));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_2041__i0 (.Q(encoder1_position[0]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFF b_prev_41 (.Q(b_prev), .C(n1795), .D(n28938));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFF direction_42 (.Q(n1800), .C(n1795), .D(n28937));   // vhdl/quadrature_decoder.vhd(48[3] 72[10])
    SB_DFFE position_2041__i1 (.Q(encoder1_position[1]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i2 (.Q(encoder1_position[2]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i3 (.Q(encoder1_position[3]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i4 (.Q(encoder1_position[4]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i5 (.Q(encoder1_position[5]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i6 (.Q(encoder1_position[6]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i7 (.Q(encoder1_position[7]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i8 (.Q(encoder1_position[8]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i9 (.Q(encoder1_position[9]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i10 (.Q(encoder1_position[10]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i11 (.Q(encoder1_position[11]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i12 (.Q(encoder1_position[12]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i13 (.Q(encoder1_position[13]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i14 (.Q(encoder1_position[14]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i15 (.Q(encoder1_position[15]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i16 (.Q(encoder1_position[16]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i17 (.Q(encoder1_position[17]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i18 (.Q(encoder1_position[18]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i19 (.Q(encoder1_position[19]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i20 (.Q(encoder1_position[20]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i21 (.Q(encoder1_position[21]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i22 (.Q(encoder1_position[22]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i23 (.Q(encoder1_position[23]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i24 (.Q(encoder1_position[24]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i25 (.Q(encoder1_position[25]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i26 (.Q(encoder1_position[26]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i27 (.Q(encoder1_position[27]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i28 (.Q(encoder1_position[28]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i29 (.Q(encoder1_position[29]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i30 (.Q(encoder1_position[30]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_DFFE position_2041__i31 (.Q(encoder1_position[31]), .C(n1795), .E(position_31__N_3836), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(62[4] 70[11])
    SB_LUT4 position_31__I_937_4_lut (.I0(a_prev), .I1(b_prev), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(position_31__N_3836));   // vhdl/quadrature_decoder.vhd(63[11:57])
    defparam position_31__I_937_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 debounce_cnt_I_936_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(\b_new[1] ), .O(debounce_cnt_N_3833));   // vhdl/quadrature_decoder.vhd(53[8:58])
    defparam debounce_cnt_I_936_4_lut.LUT_INIT = 16'h7bde;
    
endmodule
//
// Verilog Description of module coms
//

module coms (n2882, \data_out_frame[18] , clk16MHz, n55292, n29434, 
            VCC_net, \data_in_frame[18] , n55291, n55290, n29431, 
            n55289, n55288, n55242, n55287, \data_out_frame[9] , \FRAME_MATCHER.i_31__N_2509 , 
            encoder1_position_scaled, n8, rx_data, \data_in_frame[2] , 
            \data_in_frame[12] , IntegralLimit, \data_out_frame[19] , 
            n55286, n55285, n55284, n55283, n55282, \data_out_frame[3][1] , 
            n55409, \data_out_frame[8][7] , \encoder0_position_scaled[7] , 
            n55281, n55280, n55279, \data_out_frame[20] , n55278, 
            \data_out_frame[8][6] , \encoder0_position_scaled[6] , \data_out_frame[3][3] , 
            n55408, n29428, \data_out_frame[3][4] , n55407, \data_out_frame[8][5] , 
            \encoder0_position_scaled[5] , n55277, \data_out_frame[3][6] , 
            n55406, n29006, \data_in_frame[6] , \data_out_frame[3][7] , 
            n55405, n55276, \data_out_frame[8][4] , \encoder0_position_scaled[4] , 
            \data_out_frame[8][3] , \encoder0_position_scaled[3] , \data_in_frame[13] , 
            \data_out_frame[8][2] , \encoder0_position_scaled[2] , n55275, 
            n55274, \data_out_frame[7] , \encoder0_position_scaled[15] , 
            n28729, n55273, n55272, \data_out_frame[21] , n55271, 
            n55270, n55269, n55268, \data_out_frame[1][7] , GND_net, 
            n55267, n28721, n55241, n55266, \data_out_frame[1][6] , 
            \data_out_frame[22] , n55265, n55264, n55263, n55262, 
            n55261, n28713, n29424, \data_out_frame[4] , n55404, n55403, 
            \data_out_frame[1][5] , \data_out_frame[1][3] , \data_out_frame[1][1] , 
            n29421, n55260, n28711, \data_out_frame[1][0] , \data_out_frame[0][4] , 
            \data_out_frame[0][3] , \data_out_frame[0][2] , \data_out_frame[23] , 
            n55259, \data_in_frame[21] , n27934, n55419, n55402, displacement, 
            n55401, n29418, n55400, n55399, n55398, n29415, \data_in_frame[17] , 
            \data_out_frame[5] , n55397, n55396, n29409, \data_in_frame[17][5] , 
            n29406, \data_in_frame[17][4] , n55395, n29403, \data_in_frame[17][3] , 
            n55300, n29400, \data_in_frame[17][2] , n55394, n29397, 
            \data_in_frame[17][1] , n55393, n55258, n55257, n55256, 
            n28706, n55392, n55255, n55391, n55254, n29394, \data_in_frame[17][0] , 
            n28703, \data_out_frame[6] , n55390, \data_out_frame[24] , 
            n55301, n29009, n55389, n29392, \data_in_frame[16] , n55388, 
            n29389, n55387, n29384, n55386, deadband, n55253, \data_in_frame[14][6] , 
            n55252, n55251, n29381, n55250, n55249, n28696, n55299, 
            \data_out_frame[25] , n55248, n55247, \data_in_frame[20] , 
            n27932, n29378, n55246, n55245, n55244, n28689, n55385, 
            \encoder0_position_scaled[11] , \data_in_frame[15] , n28688, 
            \encoder0_position_scaled[10] , n55243, \data_out_frame[26] , 
            n55454, n55453, n55384, n55452, n55451, n55450, n55445, 
            byte_transmit_counter, \data_out_frame[17] , \data_out_frame[16] , 
            n28680, n55455, \data_out_frame[27] , n55446, n55447, 
            n55448, n55449, n55443, reset, n55444, n29012, n27898, 
            setpoint, n28672, n29374, \r_SM_Main_2__N_3545[0] , tx_active, 
            n53, n55456, \encoder0_position_scaled[9] , \FRAME_MATCHER.i[3] , 
            \FRAME_MATCHER.i[4] , \encoder0_position_scaled[8] , \FRAME_MATCHER.i[5] , 
            \byte_transmit_counter[5] , \byte_transmit_counter[6] , \byte_transmit_counter[7] , 
            n29371, n55383, n29368, \encoder0_position_scaled[14] , 
            \FRAME_MATCHER.state[3] , n8_adj_4, n56368, n29365, \data_in_frame[19] , 
            n55382, n58202, n29362, n55381, \FRAME_MATCHER.i[0] , 
            \data_in_frame[3][3] , n29359, n29356, n29353, n29015, 
            n29349, n55380, n3484, n29346, n55379, n29343, \data_in_frame[3][5] , 
            \data_in_frame[3][6] , \data_in_frame[1] , \encoder0_position_scaled[23] , 
            \data_in_frame[3][0] , \data_in_frame[19][0] , n29316, n29313, 
            n29309, n29306, n29303, n29300, n29297, n55378, n29294, 
            n29291, n29288, n29285, n29282, \data_in_frame[6][6] , 
            n29278, n29275, n29272, n29269, n29266, \data_in_frame[11] , 
            n29263, n29024, \data_in_frame[6][7] , n29258, n29255, 
            n29252, n55377, n29249, n29246, n29243, n29030, \data_in_frame[7][1] , 
            n29033, \data_in_frame[7][2] , n29042, \data_in_frame[7][4] , 
            \data_in_frame[3][7] , n29045, \data_in_frame[7][5] , n29048, 
            \data_in_frame[7][6] , n29051, \data_in_frame[7][7] , n66714, 
            n55302, n66702, n56366, n56162, n56050, n27906, \data_in_frame[21][1] , 
            n25895, n55418, n55417, n55416, n55415, n55414, n55413, 
            n55412, n55411, n55410, n55376, n55303, n55375, n55374, 
            n55373, n55372, n55371, n55370, n55369, n55368, n55367, 
            n55366, n55365, n55364, n55363, \data_out_frame[10] , 
            n55362, n55361, n55360, n55359, n55358, n55357, n55356, 
            n55355, \data_out_frame[11] , n55354, n55353, n55352, 
            n55351, n55350, n55349, n55348, n55347, \data_out_frame[12] , 
            n55346, n55345, n55344, n55343, n55342, n55341, n55340, 
            n55339, \data_out_frame[13] , n55338, n55337, n55336, 
            n55335, n55334, n55333, n55332, n55331, \data_out_frame[14] , 
            n55330, n55329, n55328, n55327, n55326, n55325, n55305, 
            n55324, \data_out_frame[15] , n55323, n55322, n55321, 
            n55320, n55319, n55318, n55317, n55304, n55316, n55315, 
            n55314, n55313, n55312, n29061, \FRAME_MATCHER.rx_data_ready_prev , 
            n55311, n55310, n55309, n55308, n55307, n55306, n55298, 
            n55297, n55296, n55295, \data_in_frame[5] , LED_c, n56120, 
            n55985, DE_c, n55294, \data_in_frame[0] , n50260, n24804, 
            n25941, n55648, \data_in_frame[6][0] , Kp_23__N_875, n50264, 
            n55624, n55775, \data_in_frame[21][2] , n25705, n32987, 
            \data_in_frame[21][3] , n25490, n55681, \data_in_frame[4] , 
            n56062, n27900, n29437, \encoder0_position_scaled[13] , 
            n29440, n28912, n29468, n29477, n29481, n29484, n29487, 
            n29493, \data_in_frame[21][0] , n29496, n29499, n29506, 
            n29509, \data_in_frame[21][4] , n29512, \data_in_frame[21][5] , 
            \data_in_frame[0][4] , n29546, \data_in_frame[23] , n29549, 
            n29552, n29555, n29558, n54697, n54695, n28940, n28946, 
            n28949, n28952, n54733, n28958, \Kp[1] , \Kp[2] , \Kp[3] , 
            \Kp[4] , \Kp[5] , \Kp[6] , \Kp[7] , \Kp[8] , \Kp[9] , 
            \Kp[10] , \Kp[11] , \Kp[12] , \Kp[13] , \Kp[14] , \Kp[15] , 
            \Ki[1] , \Ki[2] , \Ki[3] , \Ki[4] , \Ki[5] , \Ki[6] , 
            \Ki[7] , \Ki[8] , \Ki[9] , \Ki[10] , \Ki[11] , \Ki[12] , 
            \Ki[13] , \Ki[14] , \Ki[15] , n29677, neopxl_color, n29676, 
            n28961, n29674, n29673, n29671, n29670, n29669, n29668, 
            n29667, n29666, n29665, n29664, n29662, n29661, n29660, 
            n29659, n29658, n29657, n29656, n29655, n29654, control_mode, 
            n29650, n29649, n29648, n29647, n29646, current_limit, 
            n29645, n29644, n29643, n29642, n29640, n29638, n29637, 
            n29636, n29635, n29634, n29633, n29632, PWMLimit, n28964, 
            n28967, n28976, n55293, n28982, ID, n28988, n28991, 
            n28994, n28997, n28923, n28922, n28921, \Ki[0] , \Kp[0] , 
            n29000, n29003, n56059, n63134, n27904, n25933, n55668, 
            pwm_setpoint, \encoder0_position_scaled[12] , n57376, n27513, 
            n66672, n66654, n50946, n56231, n56201, n24633, n56165, 
            n22318, n50377, n66864, n66618, n56183, Kp_23__N_748, 
            \encoder0_position_scaled[22] , n73, rx_data_ready, n51197, 
            n51161, n51296, n37097, n27926, n27902, n55952, n55152, 
            n56109, n22369, n50927, n50183, n25803, n26439, n51232, 
            n55884, n27939, n55989, n63131, n25494, n4, n55181, 
            n105, control_update, n7064, n38328, n24981, n38638, 
            n6, n55149, n10, n15, n27260, n15_adj_5, n15_adj_6, 
            n55766, n56024, n38266, n38695, \encoder0_position_scaled[21] , 
            \encoder0_position_scaled[20] , \encoder0_position_scaled[19] , 
            \encoder0_position_scaled[18] , \encoder0_position_scaled[17] , 
            n50591, \encoder0_position_scaled[16] , n55151, n57943, 
            \current[7] , \current[6] , n55587, \current[5] , \current[4] , 
            \current[3] , \current[2] , \current[1] , \current[0] , 
            \current[15] , n55153, n60056, n60054, \current[11] , 
            \current[10] , \current[9] , \current[8] , \r_SM_Main[1] , 
            r_Clock_Count, n39972, tx_o, n20722, \r_SM_Main[0] , n27315, 
            n23, \o_Rx_DV_N_3488[12] , n5228, \o_Rx_DV_N_3488[24] , 
            n27, n29, n39919, n29589, \r_Bit_Index[0] , n51433, 
            n39937, n57036, n31, n58374, n58502, o_Tx_Serial_N_3598, 
            tx_enable, baudrate, r_SM_Main, r_Rx_Data, RX_N_2, r_Clock_Count_adj_20, 
            n25108, n5225, \o_Rx_DV_N_3488[8] , \o_Rx_DV_N_3488[7] , 
            \o_Rx_DV_N_3488[6] , \o_Rx_DV_N_3488[5] , \o_Rx_DV_N_3488[4] , 
            \o_Rx_DV_N_3488[3] , \o_Rx_DV_N_3488[2] , \o_Rx_DV_N_3488[1] , 
            \o_Rx_DV_N_3488[0] , n27312, n29592, \r_Bit_Index[0]_adj_17 , 
            n51425, n29596, n29582, n29581, n29580, n29578, n29577, 
            n29576, n29575, \r_SM_Main_2__N_3446[1] , n56281, n6_adj_18, 
            n55184, n58618, n4_adj_19, n27308, n58594, n58896, n58898, 
            n58932, n58844, n58970, n58934, n58880, n58952) /* synthesis syn_module_defined=1 */ ;
    input n2882;
    output [7:0]\data_out_frame[18] ;
    input clk16MHz;
    input n55292;
    input n29434;
    input VCC_net;
    output [7:0]\data_in_frame[18] ;
    input n55291;
    input n55290;
    input n29431;
    input n55289;
    input n55288;
    input n55242;
    input n55287;
    output [7:0]\data_out_frame[9] ;
    output \FRAME_MATCHER.i_31__N_2509 ;
    input [23:0]encoder1_position_scaled;
    output n8;
    output [7:0]rx_data;
    output [7:0]\data_in_frame[2] ;
    output [7:0]\data_in_frame[12] ;
    output [23:0]IntegralLimit;
    output [7:0]\data_out_frame[19] ;
    input n55286;
    input n55285;
    input n55284;
    input n55283;
    input n55282;
    output \data_out_frame[3][1] ;
    input n55409;
    output \data_out_frame[8][7] ;
    input \encoder0_position_scaled[7] ;
    input n55281;
    input n55280;
    input n55279;
    output [7:0]\data_out_frame[20] ;
    input n55278;
    output \data_out_frame[8][6] ;
    input \encoder0_position_scaled[6] ;
    output \data_out_frame[3][3] ;
    input n55408;
    input n29428;
    output \data_out_frame[3][4] ;
    input n55407;
    output \data_out_frame[8][5] ;
    input \encoder0_position_scaled[5] ;
    input n55277;
    output \data_out_frame[3][6] ;
    input n55406;
    input n29006;
    output [7:0]\data_in_frame[6] ;
    output \data_out_frame[3][7] ;
    input n55405;
    input n55276;
    output \data_out_frame[8][4] ;
    input \encoder0_position_scaled[4] ;
    output \data_out_frame[8][3] ;
    input \encoder0_position_scaled[3] ;
    output [7:0]\data_in_frame[13] ;
    output \data_out_frame[8][2] ;
    input \encoder0_position_scaled[2] ;
    input n55275;
    input n55274;
    output [7:0]\data_out_frame[7] ;
    input \encoder0_position_scaled[15] ;
    input n28729;
    input n55273;
    input n55272;
    output [7:0]\data_out_frame[21] ;
    input n55271;
    input n55270;
    input n55269;
    input n55268;
    output \data_out_frame[1][7] ;
    input GND_net;
    input n55267;
    input n28721;
    input n55241;
    input n55266;
    output \data_out_frame[1][6] ;
    output [7:0]\data_out_frame[22] ;
    input n55265;
    input n55264;
    input n55263;
    input n55262;
    input n55261;
    input n28713;
    input n29424;
    output [7:0]\data_out_frame[4] ;
    input n55404;
    input n55403;
    output \data_out_frame[1][5] ;
    output \data_out_frame[1][3] ;
    output \data_out_frame[1][1] ;
    input n29421;
    input n55260;
    input n28711;
    output \data_out_frame[1][0] ;
    output \data_out_frame[0][4] ;
    output \data_out_frame[0][3] ;
    output \data_out_frame[0][2] ;
    output [7:0]\data_out_frame[23] ;
    input n55259;
    output [7:0]\data_in_frame[21] ;
    output n27934;
    input n55419;
    input n55402;
    input [23:0]displacement;
    input n55401;
    input n29418;
    input n55400;
    input n55399;
    input n55398;
    input n29415;
    output [7:0]\data_in_frame[17] ;
    output [7:0]\data_out_frame[5] ;
    input n55397;
    input n55396;
    input n29409;
    output \data_in_frame[17][5] ;
    input n29406;
    output \data_in_frame[17][4] ;
    input n55395;
    input n29403;
    output \data_in_frame[17][3] ;
    input n55300;
    input n29400;
    output \data_in_frame[17][2] ;
    input n55394;
    input n29397;
    output \data_in_frame[17][1] ;
    input n55393;
    input n55258;
    input n55257;
    input n55256;
    input n28706;
    input n55392;
    input n55255;
    input n55391;
    input n55254;
    input n29394;
    output \data_in_frame[17][0] ;
    input n28703;
    output [7:0]\data_out_frame[6] ;
    input n55390;
    output [7:0]\data_out_frame[24] ;
    input n55301;
    input n29009;
    input n55389;
    input n29392;
    output [7:0]\data_in_frame[16] ;
    input n55388;
    input n29389;
    input n55387;
    input n29384;
    input n55386;
    output [23:0]deadband;
    input n55253;
    output \data_in_frame[14][6] ;
    input n55252;
    input n55251;
    input n29381;
    input n55250;
    input n55249;
    input n28696;
    input n55299;
    output [7:0]\data_out_frame[25] ;
    input n55248;
    input n55247;
    output [7:0]\data_in_frame[20] ;
    output n27932;
    input n29378;
    input n55246;
    input n55245;
    input n55244;
    input n28689;
    input n55385;
    input \encoder0_position_scaled[11] ;
    output [7:0]\data_in_frame[15] ;
    input n28688;
    input \encoder0_position_scaled[10] ;
    input n55243;
    output [7:0]\data_out_frame[26] ;
    input n55454;
    input n55453;
    input n55384;
    input n55452;
    input n55451;
    input n55450;
    input n55445;
    output [7:0]byte_transmit_counter;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[16] ;
    input n28680;
    input n55455;
    output [7:0]\data_out_frame[27] ;
    input n55446;
    input n55447;
    input n55448;
    input n55449;
    input n55443;
    input reset;
    input n55444;
    input n29012;
    output n27898;
    output [23:0]setpoint;
    input n28672;
    input n29374;
    output \r_SM_Main_2__N_3545[0] ;
    output tx_active;
    input n53;
    input n55456;
    input \encoder0_position_scaled[9] ;
    output \FRAME_MATCHER.i[3] ;
    output \FRAME_MATCHER.i[4] ;
    input \encoder0_position_scaled[8] ;
    output \FRAME_MATCHER.i[5] ;
    output \byte_transmit_counter[5] ;
    output \byte_transmit_counter[6] ;
    output \byte_transmit_counter[7] ;
    input n29371;
    input n55383;
    input n29368;
    input \encoder0_position_scaled[14] ;
    output \FRAME_MATCHER.state[3] ;
    output n8_adj_4;
    input n56368;
    input n29365;
    output [7:0]\data_in_frame[19] ;
    input n55382;
    output n58202;
    input n29362;
    input n55381;
    output \FRAME_MATCHER.i[0] ;
    output \data_in_frame[3][3] ;
    input n29359;
    input n29356;
    input n29353;
    input n29015;
    input n29349;
    input n55380;
    output n3484;
    input n29346;
    input n55379;
    input n29343;
    output \data_in_frame[3][5] ;
    output \data_in_frame[3][6] ;
    output [7:0]\data_in_frame[1] ;
    input \encoder0_position_scaled[23] ;
    output \data_in_frame[3][0] ;
    output \data_in_frame[19][0] ;
    input n29316;
    input n29313;
    input n29309;
    input n29306;
    input n29303;
    input n29300;
    input n29297;
    input n55378;
    input n29294;
    input n29291;
    input n29288;
    input n29285;
    input n29282;
    output \data_in_frame[6][6] ;
    input n29278;
    input n29275;
    input n29272;
    input n29269;
    input n29266;
    output [7:0]\data_in_frame[11] ;
    input n29263;
    input n29024;
    output \data_in_frame[6][7] ;
    input n29258;
    input n29255;
    input n29252;
    input n55377;
    input n29249;
    input n29246;
    input n29243;
    input n29030;
    output \data_in_frame[7][1] ;
    input n29033;
    output \data_in_frame[7][2] ;
    input n29042;
    output \data_in_frame[7][4] ;
    output \data_in_frame[3][7] ;
    input n29045;
    output \data_in_frame[7][5] ;
    input n29048;
    output \data_in_frame[7][6] ;
    input n29051;
    output \data_in_frame[7][7] ;
    output n66714;
    input n55302;
    output n66702;
    output n56366;
    input n56162;
    input n56050;
    output n27906;
    output \data_in_frame[21][1] ;
    output n25895;
    input n55418;
    input n55417;
    input n55416;
    input n55415;
    input n55414;
    input n55413;
    input n55412;
    input n55411;
    input n55410;
    input n55376;
    input n55303;
    input n55375;
    input n55374;
    input n55373;
    input n55372;
    input n55371;
    input n55370;
    input n55369;
    input n55368;
    input n55367;
    input n55366;
    input n55365;
    input n55364;
    input n55363;
    output [7:0]\data_out_frame[10] ;
    input n55362;
    input n55361;
    input n55360;
    input n55359;
    input n55358;
    input n55357;
    input n55356;
    input n55355;
    output [7:0]\data_out_frame[11] ;
    input n55354;
    input n55353;
    input n55352;
    input n55351;
    input n55350;
    input n55349;
    input n55348;
    input n55347;
    output [7:0]\data_out_frame[12] ;
    input n55346;
    input n55345;
    input n55344;
    input n55343;
    input n55342;
    input n55341;
    input n55340;
    input n55339;
    output [7:0]\data_out_frame[13] ;
    input n55338;
    input n55337;
    input n55336;
    input n55335;
    input n55334;
    input n55333;
    input n55332;
    input n55331;
    output [7:0]\data_out_frame[14] ;
    input n55330;
    input n55329;
    input n55328;
    input n55327;
    input n55326;
    input n55325;
    input n55305;
    input n55324;
    output [7:0]\data_out_frame[15] ;
    input n55323;
    input n55322;
    input n55321;
    input n55320;
    input n55319;
    input n55318;
    input n55317;
    input n55304;
    input n55316;
    input n55315;
    input n55314;
    input n55313;
    input n55312;
    input n29061;
    output \FRAME_MATCHER.rx_data_ready_prev ;
    input n55311;
    input n55310;
    input n55309;
    input n55308;
    input n55307;
    input n55306;
    input n55298;
    input n55297;
    input n55296;
    input n55295;
    output [7:0]\data_in_frame[5] ;
    output LED_c;
    input n56120;
    output n55985;
    output DE_c;
    input n55294;
    output [7:0]\data_in_frame[0] ;
    output n50260;
    output n24804;
    output n25941;
    output n55648;
    output \data_in_frame[6][0] ;
    input Kp_23__N_875;
    output n50264;
    output n55624;
    output n55775;
    output \data_in_frame[21][2] ;
    input n25705;
    input n32987;
    output \data_in_frame[21][3] ;
    input n25490;
    input n55681;
    output [7:0]\data_in_frame[4] ;
    output n56062;
    output n27900;
    input n29437;
    input \encoder0_position_scaled[13] ;
    input n29440;
    input n28912;
    input n29468;
    input n29477;
    input n29481;
    input n29484;
    input n29487;
    input n29493;
    output \data_in_frame[21][0] ;
    input n29496;
    input n29499;
    input n29506;
    input n29509;
    output \data_in_frame[21][4] ;
    input n29512;
    output \data_in_frame[21][5] ;
    output \data_in_frame[0][4] ;
    input n29546;
    output [7:0]\data_in_frame[23] ;
    input n29549;
    input n29552;
    input n29555;
    input n29558;
    input n54697;
    input n54695;
    input n28940;
    input n28946;
    input n28949;
    input n28952;
    input n54733;
    input n28958;
    output \Kp[1] ;
    output \Kp[2] ;
    output \Kp[3] ;
    output \Kp[4] ;
    output \Kp[5] ;
    output \Kp[6] ;
    output \Kp[7] ;
    output \Kp[8] ;
    output \Kp[9] ;
    output \Kp[10] ;
    output \Kp[11] ;
    output \Kp[12] ;
    output \Kp[13] ;
    output \Kp[14] ;
    output \Kp[15] ;
    output \Ki[1] ;
    output \Ki[2] ;
    output \Ki[3] ;
    output \Ki[4] ;
    output \Ki[5] ;
    output \Ki[6] ;
    output \Ki[7] ;
    output \Ki[8] ;
    output \Ki[9] ;
    output \Ki[10] ;
    output \Ki[11] ;
    output \Ki[12] ;
    output \Ki[13] ;
    output \Ki[14] ;
    output \Ki[15] ;
    input n29677;
    output [23:0]neopxl_color;
    input n29676;
    input n28961;
    input n29674;
    input n29673;
    input n29671;
    input n29670;
    input n29669;
    input n29668;
    input n29667;
    input n29666;
    input n29665;
    input n29664;
    input n29662;
    input n29661;
    input n29660;
    input n29659;
    input n29658;
    input n29657;
    input n29656;
    input n29655;
    input n29654;
    output [7:0]control_mode;
    input n29650;
    input n29649;
    input n29648;
    input n29647;
    input n29646;
    output [15:0]current_limit;
    input n29645;
    input n29644;
    input n29643;
    input n29642;
    input n29640;
    input n29638;
    input n29637;
    input n29636;
    input n29635;
    input n29634;
    input n29633;
    input n29632;
    output [23:0]PWMLimit;
    input n28964;
    input n28967;
    input n28976;
    input n55293;
    input n28982;
    input [7:0]ID;
    input n28988;
    input n28991;
    input n28994;
    input n28997;
    input n28923;
    input n28922;
    input n28921;
    output \Ki[0] ;
    output \Kp[0] ;
    input n29000;
    input n29003;
    input n56059;
    input n63134;
    output n27904;
    output n25933;
    input n55668;
    input [23:0]pwm_setpoint;
    input \encoder0_position_scaled[12] ;
    input n57376;
    output n27513;
    input n66672;
    input n66654;
    input n50946;
    output n56231;
    output n56201;
    input n24633;
    input n56165;
    output n22318;
    output n50377;
    input n66864;
    input n66618;
    input n56183;
    input Kp_23__N_748;
    input \encoder0_position_scaled[22] ;
    output n73;
    output rx_data_ready;
    output n51197;
    output n51161;
    input n51296;
    output n37097;
    output n27926;
    output n27902;
    input n55952;
    output n55152;
    input n56109;
    output n22369;
    output n50927;
    output n50183;
    output n25803;
    output n26439;
    output n51232;
    output n55884;
    input n27939;
    output n55989;
    input n63131;
    output n25494;
    output n4;
    input n55181;
    input n105;
    input control_update;
    output n7064;
    input n38328;
    output n24981;
    output n38638;
    output n6;
    output n55149;
    output n10;
    output n15;
    output n27260;
    output n15_adj_5;
    output n15_adj_6;
    input n55766;
    output n56024;
    output n38266;
    output n38695;
    input \encoder0_position_scaled[21] ;
    input \encoder0_position_scaled[20] ;
    input \encoder0_position_scaled[19] ;
    input \encoder0_position_scaled[18] ;
    input \encoder0_position_scaled[17] ;
    input n50591;
    input \encoder0_position_scaled[16] ;
    output n55151;
    output n57943;
    input \current[7] ;
    input \current[6] ;
    output n55587;
    input \current[5] ;
    input \current[4] ;
    input \current[3] ;
    input \current[2] ;
    input \current[1] ;
    input \current[0] ;
    input \current[15] ;
    output n55153;
    input n60056;
    input n60054;
    input \current[11] ;
    input \current[10] ;
    input \current[9] ;
    input \current[8] ;
    output \r_SM_Main[1] ;
    output [8:0]r_Clock_Count;
    input n39972;
    output tx_o;
    input n20722;
    output \r_SM_Main[0] ;
    output n27315;
    output n23;
    output \o_Rx_DV_N_3488[12] ;
    input n5228;
    output \o_Rx_DV_N_3488[24] ;
    output n27;
    output n29;
    output n39919;
    input n29589;
    output \r_Bit_Index[0] ;
    input n51433;
    input n39937;
    output n57036;
    output n31;
    output n58374;
    output n58502;
    output o_Tx_Serial_N_3598;
    output tx_enable;
    input [31:0]baudrate;
    output [2:0]r_SM_Main;
    output r_Rx_Data;
    input RX_N_2;
    output [7:0]r_Clock_Count_adj_20;
    output n25108;
    input n5225;
    output \o_Rx_DV_N_3488[8] ;
    output \o_Rx_DV_N_3488[7] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[0] ;
    output n27312;
    input n29592;
    output \r_Bit_Index[0]_adj_17 ;
    input n51425;
    input n29596;
    input n29582;
    input n29581;
    input n29580;
    input n29578;
    input n29577;
    input n29576;
    input n29575;
    input \r_SM_Main_2__N_3446[1] ;
    output n56281;
    output n6_adj_18;
    output n55184;
    input n58618;
    output n4_adj_19;
    output n27308;
    output n58594;
    input n58896;
    output n58898;
    input n58932;
    output n58844;
    output n58970;
    output n58934;
    output n58880;
    output n58952;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(41[6:14])
    
    wire n2, n2_adj_5286, n2_adj_5287, n2_adj_5288, n2_adj_5289, n2_adj_5290, 
        n2_adj_5291;
    wire [31:0]\FRAME_MATCHER.state_31__N_2612 ;
    
    wire n2_adj_5292, n55507, n29872, Kp_23__N_1748, n32097, n29720, 
        n2_adj_5293, n2_adj_5294, n2_adj_5295, n2_adj_5296, n2_adj_5297, 
        n2_adj_5298, n2_adj_5299, n29721, n2_adj_5300, n2_adj_5301, 
        n2_adj_5302, n2_adj_5303, n2_adj_5304, n2_adj_5305, n2_adj_5306, 
        n2_adj_5307, n2_adj_5308, n2_adj_5309, n29722, n2_adj_5310, 
        n2_adj_5311, n2_adj_5312, n2_adj_5313, n29723, n29724, n2_adj_5314, 
        n2_adj_5315, n2_adj_5316, n2_adj_5317, n2_adj_5318, n2_adj_5319, 
        n2_adj_5320, n29725, n2_adj_5321, n2_adj_5322, n2_adj_5323, 
        n2_adj_5324, n2_adj_5325, n2_adj_5326, n2_adj_5327, n2_adj_5328, 
        n2_adj_5329, n2_adj_5330, n2_adj_5331, n2_adj_5332, n2_adj_5333, 
        n2_adj_5334, n2_adj_5335, n2_adj_5336, n2_adj_5337, n2_adj_5338, 
        n2_adj_5339, n2_adj_5340, n29726, n2_adj_5341, n2_adj_5342, 
        n2_adj_5343, n2_adj_5344, n29727, n2_adj_5345, n2_adj_5346, 
        n2_adj_5347, n2_adj_5348, n54583, n2_adj_5349;
    wire [7:0]\data_in_frame[21]_c ;   // verilog/coms.v(99[12:25])
    
    wire n54683, n2_adj_5350, n29728, n2_adj_5351, n29729, n29730, 
        n2_adj_5352, n2_adj_5353, n2_adj_5354, n2_adj_5355, n2_adj_5356, 
        n29414;
    wire [7:0]\data_in_frame[17]_c ;   // verilog/coms.v(99[12:25])
    
    wire n2_adj_5357, n2_adj_5358, n2_adj_5359, n2_adj_5360, n2_adj_5361, 
        n2_adj_5362, n2_adj_5363, n2_adj_5364, n2_adj_5365, n2_adj_5366, 
        n2_adj_5367, n2_adj_5368, n2_adj_5369, n2_adj_5370, n2_adj_5371, 
        n2_adj_5372, n2_adj_5373, n2_adj_5374, n2_adj_5375;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(99[12:25])
    
    wire n29731, n2_adj_5376, n29732, n2_adj_5377, n2_adj_5378, n29733, 
        n2_adj_5379, n2_adj_5380, n2_adj_5381, n2_adj_5382, n2_adj_5383, 
        n2_adj_5384, n29490, n29734, n29735, n29736, n2_adj_5385, 
        n2_adj_5386, n2_adj_5387, n29474, n29911;
    wire [7:0]\data_in_frame[2]_c ;   // verilog/coms.v(99[12:25])
    
    wire n29875, n2_adj_5388, n2_adj_5389, n29737, n29738, n2_adj_5390, 
        n29739, n29740, n2_adj_5391, n29741, n2_adj_5392, n2_adj_5393, 
        n3, n3_adj_5394, n2_adj_5395, n3_adj_5396, n3_adj_5397, n3_adj_5398, 
        n3_adj_5399, n67035, n29742, n67038, n3_adj_5400, n29743, 
        n3_adj_5401, n3_adj_5402, n3_adj_5403, n3_adj_5404, n3_adj_5405, 
        n3_adj_5406, n2076, n3_adj_5407, n66765, n29744, n29745, 
        n29878;
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(99[12:25])
    
    wire n54807;
    wire [23:0]n4940;
    
    wire n27322, n3_adj_5408, n29746, n29747, n10_c, n55512, n161, 
        tx_transmit_N_3416, n3_adj_5409, n2_adj_5410;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(118[11:12])
    
    wire \FRAME_MATCHER.i_31__N_2507 , n63103, n1, n55431, n63080, 
        n63079, n29881, n63058, n66768, n29884, n2_adj_5411, n63056, 
        n29748, n1_adj_5412, n55430, n1_adj_5413;
    wire [7:0]byte_transmit_counter_c;   // verilog/coms.v(105[12:33])
    
    wire n55429, n1_adj_5414, n55432, n63053, n63052, n1_adj_5415, 
        n55434, n1_adj_5416, n55433, n63051, n1_adj_5417, n55435, 
        n2_adj_5418, n29749, n2_adj_5419, n63050, \FRAME_MATCHER.i_31__N_2514 , 
        n1959, n57378, n4452, n20741, n22285, n59705, n26637, 
        n3303, \FRAME_MATCHER.i_31__N_2512 , n2068, n1962, n1965, 
        n59708, n57595, n54455, n63047, n63046, n1963, n25069, 
        n20746, n29750, n2057, n771, \FRAME_MATCHER.i_31__N_2508 , 
        n2056, n63045, n29887, n63043, n27630, n27843, n49203, 
        n62946, n27628, n49202, n62958, n27626, n49201, n62959, 
        n5, n22287, n25087, n24963, n27624, n49200, n62963, n63042, 
        n29751, n9, n55145, n29752, n27622, n49199, n62966, n27620, 
        n49198, n62967, n27618, n49197, n62970, n27616, n49196, 
        n62975, n27614, n49195, n62976, n63041, n27612, n49194, 
        n63023, n29753, n27190, n27610, n49193, n63024, n57971, 
        n63040, n26633, n27608, n49192, n63027, n26634, n27606, 
        n49191, n63033;
    wire [7:0]\data_in[2] ;   // verilog/coms.v(98[12:19])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(98[12:19])
    
    wire n10_adj_5421, n27604, n49190, n63034;
    wire [7:0]\data_in[0] ;   // verilog/coms.v(98[12:19])
    
    wire n14, n25121, n27602, n49189, n63035, n20, n24976;
    wire [7:0]\data_in[1] ;   // verilog/coms.v(98[12:19])
    
    wire n19, n59864, n27600, n49188, n27598, n49187, n27596, 
        n49186, n66753, n66756, n27594, n49185, n25223, n18, n27592, 
        n49184, n27590, n49183, n27588, n49182, n27586, n49181, 
        n32103, n5_adj_5422, n66747, n27584, n49180, n25127, n20_adj_5423, 
        n27582, n49179, n27580, n49178, n15_c, n27578, n49177, 
        n4_c, n27576, n49176, n66750, n27574, n49175, n27572, 
        n49174, n27570, n49173;
    wire [31:0]n133;
    wire [7:0]\data_in_frame[19]_c ;   // verilog/coms.v(99[12:25])
    
    wire n39951, n10_adj_5424, n16, n17, n14_adj_5425, n15_adj_5426, 
        n16_adj_5427, n29340, n17_adj_5428, \FRAME_MATCHER.i_31__N_2513 , 
        n32100, n4_adj_5429, \FRAME_MATCHER.i_31__N_2511 , n6_c, n67128, 
        n8_adj_5430, n29866, n29869, n29890, n29893, n29337, n48382, 
        n55427, n29334, n48381, n29331, n29328, n29325, n29322, 
        n29319, n48380, n29312;
    wire [7:0]\data_in_frame[6]_c ;   // verilog/coms.v(99[12:25])
    
    wire n48379, n2_adj_5431, n29021, n54823;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(99[12:25])
    
    wire n2_adj_5432, n48378, n29240;
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(99[12:25])
    
    wire n29237, n29234, n55844, n29231, n29228;
    wire [7:0]\data_in_frame[1]_c ;   // verilog/coms.v(99[12:25])
    
    wire n29225, n29222, n29219, n29216;
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(99[12:25])
    
    wire n29213, n29210, n29207, n29204, n29201, n29198, n29195, 
        n29192;
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(99[12:25])
    
    wire n29189, n29186, n54827, n66717, n29054, n29057, n66720, 
        n66711, n48377, n66699, n15_adj_5433, n29160, n15_adj_5434, 
        n7, n8_adj_5435, n48376, n59598, n51148, n59602, n50620, 
        n56171, n59608, n51168, n50179, n51243, n59614, n55428, 
        n56246, n55975, n56168, n59620, n55672, n51239, n51173, 
        n59626, n55633, n55815, n59462, n50305, n55946, n55932, 
        n57892, n50370, n50368, n55892, n57445, n51150, n55972, 
        n4_adj_5436, n57531, n59424, n59426, n59428, Kp_23__N_1389, 
        n59434, n26257, n55829, n59438, n56047, Kp_23__N_1067, n59444, 
        n25345, n51414, n55819, n59450, n2_adj_5437, n2_adj_5438, 
        n2_adj_5439, n2_adj_5440, n2_adj_5441, n2_adj_5442, n2_adj_5443, 
        n2_adj_5444, n2_adj_5445, n2_adj_5446, n2_adj_5447, n2_adj_5448, 
        n2_adj_5449, n11, n2_adj_5450, n2_adj_5451, n2_adj_5452, n2_adj_5453, 
        n2_adj_5454, n2_adj_5455, n2_adj_5456, n2_adj_5457, n2_adj_5458, 
        n2_adj_5459, n2_adj_5460, n2_adj_5461, n2_adj_5462, n2_adj_5463, 
        n2_adj_5464, n2_adj_5465, n2_adj_5466, n2_adj_5467, n2_adj_5468, 
        n2_adj_5469, n2_adj_5470, n2_adj_5471, n2_adj_5472, n2_adj_5473, 
        n2_adj_5474, n2_adj_5475, n2_adj_5476, n2_adj_5477, n2_adj_5478, 
        n2_adj_5479, n2_adj_5480, n2_adj_5481, n2_adj_5482, n29095, 
        n2_adj_5483, n29094, n2_adj_5484, n29093, n2_adj_5485, n29092, 
        n2_adj_5486, n29091, n29090, n29089, n29088, n2_adj_5487, 
        n29087, n29086, n29085, n2_adj_5488, n29084, n29083, n29082, 
        n2_adj_5489, n29081, n29080, n29079, n2_adj_5490, n29078, 
        n29077, n29076, n2_adj_5491, n29075, n29074, n29073, n29072, 
        n2_adj_5492, n29071, n29070, n29069, n2_adj_5493, n29068, 
        n29067, n29066, n2_adj_5494, n29065, n2_adj_5495, n2_adj_5496, 
        n2_adj_5497, n2_adj_5498, n2_adj_5499, n2_adj_5500, n2_adj_5501, 
        n2_adj_5502, n2_adj_5503, n2_adj_5504, n56181, n56147, Kp_23__N_1518, 
        n2_adj_5505, n6_adj_5506, n25246, n55606, n55889, n59542, 
        n56159, n59548, n56138, n10_adj_5507, n55695, n27541, n56035, 
        Kp_23__N_843, n25500, n28428, n26277, n24707, n14_adj_5508, 
        n55929, n57567, n58144, n50393, n54275, n56156, n55917, 
        n59470, n51206, n55772, n55613, n58097, n59538, n55911, 
        n26520, n28387, n51247, n50907, n55757, n14_adj_5509, n56174, 
        n55978, n15_adj_5510, n1_adj_5511, n28384, n51228, n55926, 
        n7_adj_5512, n51359, n56144, n55941, n55851, n25428, n2_adj_5513, 
        n55621, n51226, n1_adj_5514, n51256, n50317, n56117, n14_adj_5515, 
        n25607, n10_adj_5516, n55704, n6_adj_5517, n55867, n57764, 
        n25337, n57296, n57981, n26, n8_adj_5518, n56041, n50272, 
        Kp_23__N_1607, n55596, n10_adj_5519, n55599, n14_adj_5520, 
        n51363, Kp_23__N_1080, n58210, n56085, n56264, n56261, n56222, 
        n14_adj_5521, n55665, n55787, n56204, n55698, n13, n58100, 
        n4_adj_5522, n26424, n26055, n25557, n56027, n55938, n58201, 
        n55569, n50310, n55968, n50498, n18_adj_5523, n56075, n56219, 
        n56004, n24, Kp_23__N_699, n22, n26_adj_5524, n51319, Kp_23__N_974, 
        n56237, n56112, n51230, n50366, n10_adj_5525, n56153, n55721, 
        n14_adj_5526, n26001, n25514, n55732, n24777, n55802, n10_adj_5527, 
        n56065, n12, n55754, n55760, n26413, n26406, n55515, n66885, 
        n66888, n25439, n59558, n59564, n59568, n59574, n50744, 
        n59580, n55684, n59586, n55652, n58045;
    wire [7:0]\data_in_frame[0]_c ;   // verilog/coms.v(99[12:25])
    
    wire n22_adj_5528, n25541, n66873, n55644, n55730, n7_adj_5529, 
        n23332, Kp_23__N_767, n26166, n4_adj_5530, n55745, n26031, 
        n51189, n25321, n25282, n25769, n6_adj_5531, n55689, n25839, 
        Kp_23__N_1085, n25572, n55923, n25481, n51250, n23345, n55808, 
        n24683, n59476, n29443, n29446, n54635, n29453, n54599, 
        n29459, n29462, n29465, n54577;
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(99[12:25])
    
    wire n59482, n29863, n29860, n29857, n29854, n29851, n29848, 
        n29845, n29842, n29839, n29836, n29833, n29830, n29827, 
        n29524, n54663, n29530, n29533, n29537, n29540, n29543, 
        n54803, n54687;
    wire [7:0]\data_in_frame[23]_c ;   // verilog/coms.v(99[12:25])
    
    wire n29597, n54743, n29719, n29718, n29717, n29716, n29715, 
        n29714, n29713, n29712, n29711, n29710, n29709, n29708, 
        n29707, n29706, n29705, n29704, n29703, n29702, n29701, 
        n29700, n29699, n29698, n29697, n29696, n29695, n29694, 
        n29693, n29692, n29691, n29690, n29689, n29688, n29687, 
        n29686, n29685, n29684, n29683, n29682, n29681, n29680, 
        n29679, n29678, n66876, n59988, n59989, n66675, n60148, 
        n60147, n66678, n29672, n29663, n29653, n29652, n29651, 
        n29641, n29639, n29631, n29630, n29629, n29628, n29627, 
        n29626, n29625, n29624, n29623, n29622, n29621, n29620, 
        n29619, n29618, n29617, n29616, n29615, n29614, n29613, 
        n29612, n29611, n29610, n29609, n54819, n54747, n26028, 
        n2_adj_5532, n28979, n50169, n24695, n25908, n66279, n12_adj_5533, 
        n28934, n10_adj_5534, n11_adj_5535, n28985, n9_adj_5536, n56072, 
        n28924, n28920, n28919, n28918, n28911, n30, n59532, n25770, 
        n55847, n50417, n59640, n20_adj_5537, n59646, n59652, n59656, 
        n55769, n59660, n59666, n55748, n50165, n56007, n59672, 
        n56078, n51223, n64943, n66867, n66636, n7_adj_5538;
    wire [7:0]tx_data;   // verilog/coms.v(108[13:20])
    
    wire Kp_23__N_709, n51294, n6_adj_5539, n25960, n66267, n55675, 
        n55560, n6_adj_5540, n6_adj_5541, n66277, n7_adj_5542, Kp_23__N_758, 
        n59488, n12_adj_5543, n14_adj_5544, n13_adj_5545, n21, n26_adj_5546, 
        n59868, n28, n32, n59732, LED_N_3408, n10_adj_5547, n56132, 
        n8_adj_5548, n7_adj_5549, n59494, n59496, n57334, n57397, 
        n58102, n8_adj_5550, n59502, n57426, n57950, n57143, n59508, 
        n59510, n10_adj_5551, n60123, n60124, n60082, n60081, n66786, 
        n63125, n60003, n60004, n57436, n60295, n60294, n59512, 
        n12_adj_5552, n62990, n9_adj_5553, n12_adj_5554, n11_adj_5555, 
        n62989, n59516, n4_adj_5556, n9_adj_5557, n57404, n59632, 
        n12_adj_5558, n11_adj_5559, n1_adj_5560, n60039, n60066, n60067, 
        n60085, n60084, n62987, n67347, n62988, n5_adj_5561, n4_adj_5562, 
        n59520, n57780, n60090, n60091, n60130, n60129, n60096, 
        n60097, n60100, n60099, n27553, n60109, n60110, n60108, 
        n63136, n66594, n65355, n63129, n60061, n60062, n60060, 
        n63135, n66582, n65357, n60145, n27637, n60146, n60144, 
        n66774, n63159, n66552, n65359, n65363, n60076, n60077, 
        n60075, n66780, n63112, n66624, n65365, n55959, n10_adj_5563, 
        n14_adj_5564, n58083, n30_adj_5565, n34, n32_adj_5566, n33, 
        n31_c, n55886, n51134, n6_adj_5567, n55896, n51146, n25648, 
        n50221, n56103, n55793, n16_adj_5568, n50685, n56088, n17_adj_5569, 
        n15_adj_5570, n56097, n15_adj_5571, n55707, n14_adj_5572, 
        n50187, n51378, n56249, n55823, n51156, n8_adj_5573, n6_adj_5574, 
        n51282, n56243, n56135, n55878, n10_adj_5575, n6_adj_5576, 
        n23288, n55714, n24672, n27511, n60079, n60080, n60078, 
        n8_adj_5577, n55965, n57163, n55551, n57177, n55902, n58178, 
        n50266, n55855, n10_adj_5578, n51154, n59783, n51265, n56234, 
        n6_adj_5579, n6_adj_5580, n50388, n55572, n6_adj_5581, n55861, 
        n55784, n66855, n50004, n50410, n12_adj_5582, n55799, n57678, 
        n57257, n51376, n51210, n57923, n29_c, n55935, n37, n25239, 
        n36, n42, n56129, n40, n41, n55790, n56177, n39, n51237, 
        n55710, n56150, n58113, n10_adj_5583, n55949, n55920, n51302, 
        n51261, n55717, n12_adj_5584, n56081, n56252, n26368, n51140, 
        n27_c, n66642, n7_adj_5585, n25271, n50298, n6_adj_5586, 
        n50391, n25385, n55763, n42_adj_5587, n50229, n40_adj_5588, 
        n55805, n50372, n41_adj_5589, n55778, n39_adj_5590, n37_adj_5591, 
        n48, n51219, n43, n38, n26337, n25687, n18_adj_5592, n57868, 
        n20_adj_5593, n57829, n7_adj_5594, n15_adj_5595, n25642, n56189, 
        n56030, n55609, n56198, n8_adj_5596, n55543, n1168, n55554, 
        n10_adj_5597, n25964, n50234, n26123, n26397, n17_adj_5598, 
        n55735, n56213, n56126, n50270, n56240, n55738, n56100, 
        n12_adj_5599, n56228, n57849, n55998, n51330, n55908, n49936, 
        n50341, n50331, n56258, n58237, n6_adj_5600, n58122, n56225, 
        n55992, n58154, n56010, n1835, n6_adj_5601, n26012, n56016, 
        n55579, n55727, n50249, n6_adj_5602, n14_adj_5603, n15_adj_5604, 
        n14_adj_5605, n13_adj_5606, n55678, n24677, n25996, n14_adj_5607, 
        n26092, n57840, n13_adj_5608, n26378, n26187, n18_adj_5609, 
        n56195, n17_adj_5610, n25820, n37_adj_5611, n19_adj_5612, 
        n66843, n66606, n7_adj_5613, n55751, n56094, n1516, n56123, 
        n55630, n12_adj_5614, n55995, n56186, n10_adj_5615, n55590, 
        n66837, n50190, n25656, n26267, n66804, n7_adj_5616, n55796, 
        n55498, n56210, n56001, n24_adj_5617, n55781, n22_adj_5618, 
        n26_adj_5619, n55864, n58238, n24_adj_5620, n56091, n22_adj_5621, 
        n18_adj_5622, n56207, n26_adj_5623, n56053, n1699, n1130, 
        n10_adj_5625, n66831, n10_adj_5626, n7_adj_5627, n14_adj_5628, 
        n26960, n56056, n10_adj_5629, n55662, n56019, n1720, n66825, 
        n55873, n6_adj_5630, n55742, n25661, n10_adj_5631, n25915, 
        n12_adj_5632, n33_adj_5633, n55636, n56044, n66798, n7_adj_5635, 
        n10_adj_5636, n1191, n6_adj_5637, n7_adj_5638, n58239, n40_adj_5639, 
        n38_adj_5640, n56192, n39_adj_5641, n26479, n37_adj_5642, 
        n66813, n42_adj_5643, n60040, n46, n41_adj_5644, n58240, 
        n12_adj_5645, n55565, n55575, n10_adj_5646, n10_adj_5647, 
        n30_adj_5648, n4_adj_5649, n47470, n6_adj_5654, n8_adj_5655, 
        n59336, n27862, n66645, n14_adj_5656, n66639, n66807, n60044, 
        n66633, n66588, n66576, n66627, n66630, n66621, n66801, 
        n66795, n66789, n66792, n66783, n23_c, n27_adj_5657, n66777, 
        n29_adj_5658, n31_adj_5659, n66771, n66603, n66591, n66585, 
        n66579, n66573, n27860, n66558, n65305, n65306, n66546, 
        n66561, n66555, n66549, n66543;
    
    SB_DFFESS data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2), .S(n55292));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i150 (.Q(\data_in_frame[18] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29434));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5286), .S(n55291));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5287), .S(n55290));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i149 (.Q(\data_in_frame[18] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29431));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5288), .S(n55289));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5289), .S(n55288));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5290), .S(n55242));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5291), .S(n55287));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_72_i2_4_lut (.I0(\data_out_frame[9] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5292));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_72_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14027_3_lut_4_lut (.I0(n8), .I1(n55507), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n29872));
    defparam i14027_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13875_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[12] [3]), 
            .I3(IntegralLimit[11]), .O(n29720));   // verilog/coms.v(148[4] 304[11])
    defparam i13875_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5293), .S(n55286));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5294), .S(n55285));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5295), .S(n55284));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5296), .S(n55283));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5297), .S(n55282));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i26 (.Q(\data_out_frame[3][1] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5298), .S(n55409));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_71_i2_4_lut (.I0(\data_out_frame[8][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5299));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_71_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13876_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[12] [2]), 
            .I3(IntegralLimit[10]), .O(n29721));   // verilog/coms.v(148[4] 304[11])
    defparam i13876_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5300), .S(n55281));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5301), .S(n55280));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5302), .S(n55279));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5303), .S(n55278));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_70_i2_4_lut (.I0(\data_out_frame[8][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5304));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_70_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i28 (.Q(\data_out_frame[3][3] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5305), .S(n55408));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i148 (.Q(\data_in_frame[18] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29428));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i29 (.Q(\data_out_frame[3][4] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5306), .S(n55407));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_69_i2_4_lut (.I0(\data_out_frame[8][5] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5307));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_69_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5308), .S(n55277));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i31 (.Q(\data_out_frame[3][6] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5309), .S(n55406));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13877_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[12] [1]), 
            .I3(IntegralLimit[9]), .O(n29722));   // verilog/coms.v(148[4] 304[11])
    defparam i13877_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF data_in_frame_0___i50 (.Q(\data_in_frame[6] [1]), .C(clk16MHz), 
           .D(n29006));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i32 (.Q(\data_out_frame[3][7] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5310), .S(n55405));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5311), .S(n55276));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_68_i2_4_lut (.I0(\data_out_frame[8][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[4] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5312));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_68_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_67_i2_4_lut (.I0(\data_out_frame[8][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[3] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5313));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_67_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13878_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[12] [0]), 
            .I3(IntegralLimit[8]), .O(n29723));   // verilog/coms.v(148[4] 304[11])
    defparam i13878_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13879_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[13] [7]), 
            .I3(IntegralLimit[7]), .O(n29724));   // verilog/coms.v(148[4] 304[11])
    defparam i13879_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_4_lut (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[8][2] ), 
            .I2(\encoder0_position_scaled[2] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5314));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_DFFESS data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5315), .S(n55275));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5316), .S(n55274));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_63_i2_4_lut (.I0(\data_out_frame[7] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5317));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_63_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5318), .S(n28729));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5319), .S(n55273));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5320), .S(n55272));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13880_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[13] [6]), 
            .I3(IntegralLimit[6]), .O(n29725));   // verilog/coms.v(148[4] 304[11])
    defparam i13880_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5321), .S(n55271));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5322), .S(n55270));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5323), .S(n55269));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5324), .S(n55268));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_15_i2_3_lut (.I0(\data_out_frame[1][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5325));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_15_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFESS data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5326), .S(n55267));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5327), .S(n28721));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5328), .S(n55241));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5329), .S(n55266));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_14_i2_3_lut (.I0(\data_out_frame[1][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5330));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_14_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFESS data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5331), .S(n55265));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5332), .S(n55264));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5333), .S(n55263));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5334), .S(n55262));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5335), .S(n55261));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5336), .S(n28713));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i147 (.Q(\data_in_frame[18] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29424));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5337), .S(n55404));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5338), .S(n55403));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_13_i2_3_lut (.I0(\data_out_frame[1][5] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5339));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_13_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_787_Select_11_i2_3_lut (.I0(\data_out_frame[1][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5340));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_11_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13881_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[13] [5]), 
            .I3(IntegralLimit[5]), .O(n29726));   // verilog/coms.v(148[4] 304[11])
    defparam i13881_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_9_i2_3_lut (.I0(\data_out_frame[1][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5341));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_9_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFE data_in_frame_0___i146 (.Q(\data_in_frame[18] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29421));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5342), .S(n55260));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5343), .S(n28711));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_8_i2_3_lut (.I0(\data_out_frame[1][0] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5344));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_8_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13882_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[13] [4]), 
            .I3(IntegralLimit[4]), .O(n29727));   // verilog/coms.v(148[4] 304[11])
    defparam i13882_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_4_i2_3_lut (.I0(\data_out_frame[0][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5345));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_4_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_787_Select_3_i2_3_lut (.I0(\data_out_frame[0][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5346));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_3_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 select_787_Select_2_i2_3_lut (.I0(\data_out_frame[0][2] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5347));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_2_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFESS data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5348), .S(n55259));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i49194_3_lut (.I0(rx_data[7]), .I1(\data_in_frame[21] [7]), 
            .I2(n27934), .I3(GND_net), .O(n54583));   // verilog/coms.v(94[13:20])
    defparam i49194_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5349), .S(n55419));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i49196_3_lut (.I0(rx_data[6]), .I1(\data_in_frame[21]_c [6]), 
            .I2(n27934), .I3(GND_net), .O(n54683));   // verilog/coms.v(94[13:20])
    defparam i49196_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5350), .S(n55402));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_157_i2_4_lut (.I0(\data_out_frame[19] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5300));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_157_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13883_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[13] [3]), 
            .I3(IntegralLimit[3]), .O(n29728));   // verilog/coms.v(148[4] 304[11])
    defparam i13883_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5351), .S(n55401));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i145 (.Q(\data_in_frame[18] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29418));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13884_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[13] [2]), 
            .I3(IntegralLimit[2]), .O(n29729));   // verilog/coms.v(148[4] 304[11])
    defparam i13884_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13885_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[13] [1]), 
            .I3(IntegralLimit[1]), .O(n29730));   // verilog/coms.v(148[4] 304[11])
    defparam i13885_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5352), .S(n55400));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5353), .S(n55399));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5354), .S(n55398));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i144 (.Q(\data_in_frame[17] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29415));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5355), .S(n55397));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5356), .S(n55396));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i143 (.Q(\data_in_frame[17]_c [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29414));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i142 (.Q(\data_in_frame[17][5] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29409));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i141 (.Q(\data_in_frame[17][4] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29406));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5357), .S(n55395));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i140 (.Q(\data_in_frame[17][3] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29403));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5358), .S(n55300));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i139 (.Q(\data_in_frame[17][2] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29400));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5359), .S(n55394));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i138 (.Q(\data_in_frame[17][1] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29397));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5360), .S(n55393));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5361), .S(n55258));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5362), .S(n55257));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5363), .S(n55256));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5364), .S(n28706));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5365), .S(n55392));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5366), .S(n55255));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5367), .S(n55391));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5368), .S(n55254));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i137 (.Q(\data_in_frame[17][0] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29394));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5369), .S(n28703));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5370), .S(n55390));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5371), .S(n55301));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i51 (.Q(\data_in_frame[6] [2]), .C(clk16MHz), 
           .D(n29009));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5372), .S(n55389));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i136 (.Q(\data_in_frame[16] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29392));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5373), .S(n55388));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i135 (.Q(\data_in_frame[16] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29389));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5374), .S(n55387));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i134 (.Q(\data_in_frame[16] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29384));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5375), .S(n55386));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13886_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[14] [7]), 
            .I3(deadband[23]), .O(n29731));   // verilog/coms.v(148[4] 304[11])
    defparam i13886_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5376), .S(n55253));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13887_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[14][6] ), 
            .I3(deadband[22]), .O(n29732));   // verilog/coms.v(148[4] 304[11])
    defparam i13887_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5377), .S(n55252));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5378), .S(n55251));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i133 (.Q(\data_in_frame[16] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29381));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13888_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[14] [5]), 
            .I3(deadband[21]), .O(n29733));   // verilog/coms.v(148[4] 304[11])
    defparam i13888_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5379), .S(n55250));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5380), .S(n55249));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5381), .S(n28696));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5382), .S(n55299));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5383), .S(n55248));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5384), .S(n55247));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13645_3_lut (.I0(\data_in_frame[20] [7]), .I1(rx_data[7]), 
            .I2(n27932), .I3(GND_net), .O(n29490));   // verilog/coms.v(130[12] 305[6])
    defparam i13645_3_lut.LUT_INIT = 16'hacac;
    SB_DFFE data_in_frame_0___i132 (.Q(\data_in_frame[16] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29378));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13889_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[14] [4]), 
            .I3(deadband[20]), .O(n29734));   // verilog/coms.v(148[4] 304[11])
    defparam i13889_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13890_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[14] [3]), 
            .I3(deadband[19]), .O(n29735));   // verilog/coms.v(148[4] 304[11])
    defparam i13890_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13891_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[14] [2]), 
            .I3(deadband[18]), .O(n29736));   // verilog/coms.v(148[4] 304[11])
    defparam i13891_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5385), .S(n55246));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5386), .S(n55245));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5387), .S(n55244));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13629_3_lut (.I0(\data_in_frame[20] [2]), .I1(rx_data[2]), 
            .I2(n27932), .I3(GND_net), .O(n29474));   // verilog/coms.v(130[12] 305[6])
    defparam i13629_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19059_3_lut (.I0(n27932), .I1(rx_data[1]), .I2(\data_in_frame[20] [1]), 
            .I3(GND_net), .O(n29911));   // verilog/coms.v(94[13:20])
    defparam i19059_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14030_3_lut_4_lut (.I0(n8), .I1(n55507), .I2(rx_data[1]), 
            .I3(\data_in_frame[2]_c [1]), .O(n29875));
    defparam i14030_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESS data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5388), .S(n28689));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5389), .S(n55385));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13892_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[14] [1]), 
            .I3(deadband[17]), .O(n29737));   // verilog/coms.v(148[4] 304[11])
    defparam i13892_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13893_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[14] [0]), 
            .I3(deadband[16]), .O(n29738));   // verilog/coms.v(148[4] 304[11])
    defparam i13893_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_59_i2_4_lut (.I0(\data_out_frame[7] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[11] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5390));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_59_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13894_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[15] [7]), 
            .I3(deadband[15]), .O(n29739));   // verilog/coms.v(148[4] 304[11])
    defparam i13894_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13895_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[15] [6]), 
            .I3(deadband[14]), .O(n29740));   // verilog/coms.v(148[4] 304[11])
    defparam i13895_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5391), .S(n28688));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13896_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[15] [5]), 
            .I3(deadband[13]), .O(n29741));   // verilog/coms.v(148[4] 304[11])
    defparam i13896_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_58_i2_4_lut (.I0(\data_out_frame[7] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[10] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5392));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_58_i2_4_lut.LUT_INIT = 16'hc088;
    SB_DFFESS data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5393), .S(n55243));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk16MHz), 
            .E(n2882), .D(n3), .S(n55454));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk16MHz), 
            .E(n2882), .D(n3_adj_5394), .S(n55453));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5395), .S(n55384));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk16MHz), 
            .E(n2882), .D(n3_adj_5396), .S(n55452));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk16MHz), 
            .E(n2882), .D(n3_adj_5397), .S(n55451));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk16MHz), 
            .E(n2882), .D(n3_adj_5398), .S(n55450));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk16MHz), 
            .E(n2882), .D(n3_adj_5399), .S(n55445));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(byte_transmit_counter[1]), .O(n67035));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i13897_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[15] [4]), 
            .I3(deadband[12]), .O(n29742));   // verilog/coms.v(148[4] 304[11])
    defparam i13897_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n67035_bdd_4_lut (.I0(n67035), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(byte_transmit_counter[1]), 
            .O(n67038));
    defparam n67035_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESS data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk16MHz), 
            .E(n2882), .D(n3_adj_5400), .S(n28680));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13898_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[15] [3]), 
            .I3(deadband[11]), .O(n29743));   // verilog/coms.v(148[4] 304[11])
    defparam i13898_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk16MHz), 
            .E(n2882), .D(n3_adj_5401), .S(n55455));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk16MHz), 
            .E(n2882), .D(n3_adj_5402), .S(n55446));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk16MHz), 
            .E(n2882), .D(n3_adj_5403), .S(n55447));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk16MHz), 
            .E(n2882), .D(n3_adj_5404), .S(n55448));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk16MHz), 
            .E(n2882), .D(n3_adj_5405), .S(n55449));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk16MHz), 
            .E(n2882), .D(n3_adj_5406), .S(n55443));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR \FRAME_MATCHER.state_FSM_i1  (.Q(Kp_23__N_1748), .C(clk16MHz), 
            .D(n2076), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFESS data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk16MHz), 
            .E(n2882), .D(n3_adj_5407), .S(n55444));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49666 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(byte_transmit_counter[1]), .O(n66765));
    defparam byte_transmit_counter_0__bdd_4_lut_49666.LUT_INIT = 16'he4aa;
    SB_LUT4 i13899_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[15] [2]), 
            .I3(deadband[10]), .O(n29744));   // verilog/coms.v(148[4] 304[11])
    defparam i13899_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13900_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[15] [1]), 
            .I3(deadband[9]), .O(n29745));   // verilog/coms.v(148[4] 304[11])
    defparam i13900_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14033_3_lut_4_lut (.I0(n8), .I1(n55507), .I2(rx_data[2]), 
            .I3(\data_in_frame[2]_c [2]), .O(n29878));
    defparam i14033_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0___i52 (.Q(\data_in_frame[6] [3]), .C(clk16MHz), 
           .D(n29012));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i49200_3_lut (.I0(rx_data[1]), .I1(\data_in_frame[3] [1]), .I2(n27898), 
            .I3(GND_net), .O(n54807));   // verilog/coms.v(94[13:20])
    defparam i49200_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFER setpoint_i0_i0 (.Q(setpoint[0]), .C(clk16MHz), .E(n27322), 
            .D(n4940[0]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk16MHz), 
            .E(n2882), .D(n3_adj_5408), .S(n28672));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i131 (.Q(\data_in_frame[16] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29374));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13901_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[15] [0]), 
            .I3(deadband[8]), .O(n29746));   // verilog/coms.v(148[4] 304[11])
    defparam i13901_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13902_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[16] [7]), 
            .I3(deadband[7]), .O(n29747));   // verilog/coms.v(148[4] 304[11])
    defparam i13902_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i39369_4_lut (.I0(reset), .I1(n10_c), .I2(n55512), .I3(n161), 
            .O(n27898));
    defparam i39369_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i49264_3_lut (.I0(\r_SM_Main_2__N_3545[0] ), .I1(tx_active), 
            .I2(n53), .I3(GND_net), .O(tx_transmit_N_3416));
    defparam i49264_3_lut.LUT_INIT = 16'h0101;
    SB_DFFESS data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk16MHz), 
            .E(n2882), .D(n3_adj_5409), .S(n55456));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 select_787_Select_57_i2_4_lut (.I0(\data_out_frame[7] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[9] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5410));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_57_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i46796_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63103));   // verilog/coms.v(158[12:15])
    defparam i46796_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk16MHz), 
            .E(n2882), .D(n1), .S(n55431));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i46489_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63080));   // verilog/coms.v(158[12:15])
    defparam i46489_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i47062_2_lut (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63079));   // verilog/coms.v(158[12:15])
    defparam i47062_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14036_3_lut_4_lut (.I0(n8), .I1(n55507), .I2(rx_data[3]), 
            .I3(\data_in_frame[2]_c [3]), .O(n29881));
    defparam i14036_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i46421_2_lut (.I0(\FRAME_MATCHER.i[4] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63058));   // verilog/coms.v(158[12:15])
    defparam i46421_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 n66765_bdd_4_lut (.I0(n66765), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(byte_transmit_counter[1]), 
            .O(n66768));
    defparam n66765_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14039_3_lut_4_lut (.I0(n8), .I1(n55507), .I2(rx_data[4]), 
            .I3(\data_in_frame[2]_c [4]), .O(n29884));
    defparam i14039_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_56_i2_4_lut (.I0(\data_out_frame[7] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[8] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5411));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_56_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i46356_2_lut (.I0(\FRAME_MATCHER.i[5] ), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63056));   // verilog/coms.v(158[12:15])
    defparam i46356_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13903_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[16] [6]), 
            .I3(deadband[6]), .O(n29748));   // verilog/coms.v(148[4] 304[11])
    defparam i13903_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFESS byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk16MHz), 
            .E(n2882), .D(n1_adj_5412), .S(n55430));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter_c[3]), 
            .C(clk16MHz), .E(n2882), .D(n1_adj_5413), .S(n55429));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter_c[4]), 
            .C(clk16MHz), .E(n2882), .D(n1_adj_5414), .S(n55432));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i46410_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63053));   // verilog/coms.v(158[12:15])
    defparam i46410_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i46409_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63052));   // verilog/coms.v(158[12:15])
    defparam i46409_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS byte_transmit_counter_i0_i5 (.Q(\byte_transmit_counter[5] ), 
            .C(clk16MHz), .E(n2882), .D(n1_adj_5415), .S(n55434));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS byte_transmit_counter_i0_i6 (.Q(\byte_transmit_counter[6] ), 
            .C(clk16MHz), .E(n2882), .D(n1_adj_5416), .S(n55433));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i46408_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63051));   // verilog/coms.v(158[12:15])
    defparam i46408_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS byte_transmit_counter_i0_i7 (.Q(\byte_transmit_counter[7] ), 
            .C(clk16MHz), .E(n2882), .D(n1_adj_5417), .S(n55435));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i130 (.Q(\data_in_frame[16] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29371));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5418), .S(n55383));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i13904_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[16] [5]), 
            .I3(deadband[5]), .O(n29749));   // verilog/coms.v(148[4] 304[11])
    defparam i13904_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE data_in_frame_0___i129 (.Q(\data_in_frame[16] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29368));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1090 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[7] [6]), 
            .I2(\encoder0_position_scaled[14] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5419));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1090.LUT_INIT = 16'ha088;
    SB_LUT4 i46406_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63050));   // verilog/coms.v(158[12:15])
    defparam i46406_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5246_4_lut (.I0(\FRAME_MATCHER.i_31__N_2514 ), .I1(n1959), 
            .I2(n57378), .I3(n4452), .O(n20741));   // verilog/coms.v(148[4] 304[11])
    defparam i5246_4_lut.LUT_INIT = 16'ha0a2;
    SB_LUT4 i1_4_lut_adj_1091 (.I0(n20741), .I1(n1959), .I2(n22285), .I3(n59705), 
            .O(n26637));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1091.LUT_INIT = 16'hbbba;
    SB_LUT4 i460_2_lut (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), .I2(GND_net), 
            .I3(GND_net), .O(n2068));   // verilog/coms.v(148[4] 304[11])
    defparam i460_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i42661_4_lut (.I0(n1959), .I1(n1962), .I2(n3303), .I3(n1965), 
            .O(n59708));   // verilog/coms.v(139[4] 141[7])
    defparam i42661_4_lut.LUT_INIT = 16'h0a02;
    SB_LUT4 i1_4_lut_adj_1092 (.I0(\FRAME_MATCHER.i_31__N_2512 ), .I1(n1962), 
            .I2(n59708), .I3(n57595), .O(n54455));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1092.LUT_INIT = 16'hb3a0;
    SB_LUT4 i46401_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63047));   // verilog/coms.v(158[12:15])
    defparam i46401_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i46394_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63046));   // verilog/coms.v(158[12:15])
    defparam i46394_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5251_4_lut (.I0(n1963), .I1(\FRAME_MATCHER.state[3] ), .I2(n1965), 
            .I3(n25069), .O(n20746));   // verilog/coms.v(148[4] 304[11])
    defparam i5251_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i13905_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[16] [4]), 
            .I3(deadband[4]), .O(n29750));   // verilog/coms.v(148[4] 304[11])
    defparam i13905_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i449_2_lut (.I0(\FRAME_MATCHER.state_31__N_2612 [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(GND_net), .I3(GND_net), .O(n2057));   // verilog/coms.v(148[4] 304[11])
    defparam i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i448_2_lut (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), .I2(GND_net), 
            .I3(GND_net), .O(n2056));   // verilog/coms.v(148[4] 304[11])
    defparam i448_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46411_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63045));   // verilog/coms.v(158[12:15])
    defparam i46411_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14042_3_lut_4_lut (.I0(n8), .I1(n55507), .I2(rx_data[5]), 
            .I3(\data_in_frame[2]_c [5]), .O(n29887));
    defparam i14042_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i46392_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63043));   // verilog/coms.v(158[12:15])
    defparam i46392_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_33_lut  (.I0(n62946), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [31]), .I3(n49203), .O(n27630)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_33_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_32_lut  (.I0(n62958), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [30]), .I3(n49202), .O(n27628)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_32_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_32  (.CI(n49202), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [30]), .CO(n49203));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_31_lut  (.I0(n62959), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [29]), .I3(n49201), .O(n27626)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_31_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i22648_4_lut (.I0(n5), .I1(\FRAME_MATCHER.i [31]), .I2(\FRAME_MATCHER.i [2]), 
            .I3(\FRAME_MATCHER.i[3] ), .O(n771));   // verilog/coms.v(160[9:60])
    defparam i22648_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i2_2_lut (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), .I2(GND_net), 
            .I3(GND_net), .O(n22287));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut (.I0(\FRAME_MATCHER.i[4] ), .I1(n25087), .I2(GND_net), 
            .I3(GND_net), .O(n24963));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_31  (.CI(n49201), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [29]), .CO(n49202));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_30_lut  (.I0(n62963), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [28]), .I3(n49200), .O(n27624)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_30_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i46391_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63042));   // verilog/coms.v(158[12:15])
    defparam i46391_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13906_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[16] [3]), 
            .I3(deadband[3]), .O(n29751));   // verilog/coms.v(148[4] 304[11])
    defparam i13906_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i22653_4_lut (.I0(n8_adj_4), .I1(\FRAME_MATCHER.i [31]), .I2(n24963), 
            .I3(\FRAME_MATCHER.i[3] ), .O(n3303));   // verilog/coms.v(230[9:54])
    defparam i22653_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i3_4_lut (.I0(n56368), .I1(\FRAME_MATCHER.i[3] ), .I2(reset), 
            .I3(n9), .O(n55145));   // verilog/coms.v(157[7:23])
    defparam i3_4_lut.LUT_INIT = 16'hfff7;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_30  (.CI(n49200), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [28]), .CO(n49201));
    SB_LUT4 i13907_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[16] [2]), 
            .I3(deadband[2]), .O(n29752));   // verilog/coms.v(148[4] 304[11])
    defparam i13907_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_29_lut  (.I0(n62966), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [27]), .I3(n49199), .O(n27622)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_29_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_29  (.CI(n49199), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [27]), .CO(n49200));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_28_lut  (.I0(n62967), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [26]), .I3(n49198), .O(n27620)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_28_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_28  (.CI(n49198), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [26]), .CO(n49199));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_27_lut  (.I0(n62970), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [25]), .I3(n49197), .O(n27618)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_27_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_27  (.CI(n49197), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [25]), .CO(n49198));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_26_lut  (.I0(n62975), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [24]), .I3(n49196), .O(n27616)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_26_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_26  (.CI(n49196), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [24]), .CO(n49197));
    SB_LUT4 i2_2_lut_adj_1093 (.I0(n3303), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(GND_net), .I3(GND_net), .O(n22285));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_adj_1093.LUT_INIT = 16'h4444;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_25_lut  (.I0(n62976), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [23]), .I3(n49195), .O(n27614)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_25_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_25  (.CI(n49195), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [23]), .CO(n49196));
    SB_LUT4 i46390_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63041));   // verilog/coms.v(158[12:15])
    defparam i46390_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_24_lut  (.I0(n63023), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [22]), .I3(n49194), .O(n27612)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_24_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i13908_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[16] [1]), 
            .I3(deadband[1]), .O(n29753));   // verilog/coms.v(148[4] 304[11])
    defparam i13908_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_24  (.CI(n49194), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [22]), .CO(n49195));
    SB_LUT4 i3_2_lut (.I0(n25069), .I1(\FRAME_MATCHER.i_31__N_2507 ), .I2(GND_net), 
            .I3(GND_net), .O(n27190));   // verilog/coms.v(148[4] 304[11])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_23_lut  (.I0(n63024), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [21]), .I3(n49193), .O(n27610)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_23_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i2_4_lut (.I0(n4452), .I1(n27190), .I2(\FRAME_MATCHER.i_31__N_2514 ), 
            .I3(n22285), .O(n57971));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut.LUT_INIT = 16'hffdc;
    SB_LUT4 i46238_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63040));   // verilog/coms.v(158[12:15])
    defparam i46238_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1094 (.I0(n1965), .I1(n1959), .I2(n57971), .I3(n1962), 
            .O(n26633));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1094.LUT_INIT = 16'h4000;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_23  (.CI(n49193), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [21]), .CO(n49194));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_22_lut  (.I0(n63027), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [20]), .I3(n49192), .O(n27608)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_22_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_4_lut_adj_1095 (.I0(n1962), .I1(n26633), .I2(n1959), .I3(n22287), 
            .O(n26634));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1095.LUT_INIT = 16'heccc;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_22  (.CI(n49192), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [20]), .CO(n49193));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_21_lut  (.I0(n63033), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [19]), .I3(n49191), .O(n27606)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_21_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_21  (.CI(n49191), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [19]), .CO(n49192));
    SB_LUT4 i2_2_lut_adj_1096 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5421));
    defparam i2_2_lut_adj_1096.LUT_INIT = 16'heeee;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_20_lut  (.I0(n63034), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [18]), .I3(n49190), .O(n27604)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_20_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_20  (.CI(n49190), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [18]), .CO(n49191));
    SB_LUT4 i6_4_lut (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), .I2(\data_in[3] [1]), 
            .I3(\data_in[0] [7]), .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut (.I0(\data_in[3] [6]), .I1(n14), .I2(n10_adj_5421), 
            .I3(\data_in[2] [1]), .O(n25121));
    defparam i7_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_19_lut  (.I0(n63035), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [17]), .I3(n49189), .O(n27602)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_19_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i46389_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63035));   // verilog/coms.v(158[12:15])
    defparam i46389_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i8_4_lut (.I0(\data_in[2] [6]), .I1(\data_in[2] [0]), .I2(n25121), 
            .I3(\data_in[0] [5]), .O(n20));
    defparam i8_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i46388_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63034));   // verilog/coms.v(158[12:15])
    defparam i46388_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i46232_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63033));   // verilog/coms.v(158[12:15])
    defparam i46232_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i7_4_lut_adj_1097 (.I0(n24976), .I1(\data_in[3] [7]), .I2(\data_in[1] [6]), 
            .I3(\data_in[2] [5]), .O(n19));
    defparam i7_4_lut_adj_1097.LUT_INIT = 16'hfeff;
    SB_LUT4 i42811_4_lut (.I0(\data_in[1] [2]), .I1(\data_in[1] [3]), .I2(\data_in[0] [1]), 
            .I3(\data_in[3] [2]), .O(n59864));
    defparam i42811_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_19  (.CI(n49189), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [17]), .CO(n49190));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_18_lut  (.I0(n63040), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [16]), .I3(n49188), .O(n27600)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_18_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_18  (.CI(n49188), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [16]), .CO(n49189));
    SB_LUT4 i46341_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63027));   // verilog/coms.v(158[12:15])
    defparam i46341_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i11_3_lut (.I0(n59864), .I1(n19), .I2(n20), .I3(GND_net), 
            .O(n1959));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_17_lut  (.I0(n63041), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [15]), .I3(n49187), .O(n27598)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_17_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_17  (.CI(n49187), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [15]), .CO(n49188));
    SB_DFFE data_in_frame_0___i128 (.Q(\data_in_frame[15] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29365));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_16_lut  (.I0(n63042), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [14]), .I3(n49186), .O(n27596)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_16_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_16  (.CI(n49186), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [14]), .CO(n49187));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49661 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n66753));
    defparam byte_transmit_counter_0__bdd_4_lut_49661.LUT_INIT = 16'he4aa;
    SB_LUT4 n66753_bdd_4_lut (.I0(n66753), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n66756));
    defparam n66753_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_15_lut  (.I0(n63043), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [13]), .I3(n49185), .O(n27594)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_15_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_15  (.CI(n49185), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [13]), .CO(n49186));
    SB_LUT4 i7_4_lut_adj_1098 (.I0(\data_in[2] [4]), .I1(n25121), .I2(\data_in[1] [5]), 
            .I3(n25223), .O(n18));
    defparam i7_4_lut_adj_1098.LUT_INIT = 16'hfffd;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_14_lut  (.I0(n63045), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [12]), .I3(n49184), .O(n27592)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_14_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_14  (.CI(n49184), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [12]), .CO(n49185));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_13_lut  (.I0(n63046), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [11]), .I3(n49183), .O(n27590)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_13_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_13  (.CI(n49183), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [11]), .CO(n49184));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_12_lut  (.I0(n63047), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [10]), .I3(n49182), .O(n27588)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_12_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_12  (.CI(n49182), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [10]), .CO(n49183));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_11_lut  (.I0(n63050), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [9]), .I3(n49181), .O(n27586)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_11_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_2_lut_3_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(n32103), 
            .I3(GND_net), .O(n5_adj_5422));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49651 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [3]), .I2(\data_out_frame[19] [3]), 
            .I3(byte_transmit_counter[1]), .O(n66747));
    defparam byte_transmit_counter_0__bdd_4_lut_49651.LUT_INIT = 16'he4aa;
    SB_LUT4 i19166_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[3] [1]), 
            .I3(\data_in_frame[19] [1]), .O(n4940[1]));   // verilog/coms.v(148[4] 304[11])
    defparam i19166_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_11  (.CI(n49181), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [9]), .CO(n49182));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_10_lut  (.I0(n63051), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [8]), .I3(n49180), .O(n27584)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_10_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i9_4_lut (.I0(\data_in[0] [6]), .I1(n18), .I2(\data_in[3] [0]), 
            .I3(n25127), .O(n20_adj_5423));
    defparam i9_4_lut.LUT_INIT = 16'hfffd;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_10  (.CI(n49180), .I0(n27843), 
            .I1(\FRAME_MATCHER.i [8]), .CO(n49181));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_9_lut  (.I0(n63052), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [7]), .I3(n49179), .O(n27582)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_9_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i46376_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63024));   // verilog/coms.v(158[12:15])
    defparam i46376_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_9  (.CI(n49179), .I0(n27843), .I1(\FRAME_MATCHER.i [7]), 
            .CO(n49180));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_8_lut  (.I0(n63053), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [6]), .I3(n49178), .O(n27580)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_8_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i4_2_lut (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n15_c));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i46398_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n63023));   // verilog/coms.v(158[12:15])
    defparam i46398_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_8  (.CI(n49178), .I0(n27843), .I1(\FRAME_MATCHER.i [6]), 
            .CO(n49179));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_7_lut  (.I0(n63056), .I1(n27843), 
            .I2(\FRAME_MATCHER.i[5] ), .I3(n49177), .O(n27578)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_7_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_7  (.CI(n49177), .I0(n27843), .I1(\FRAME_MATCHER.i[5] ), 
            .CO(n49178));
    SB_LUT4 i10_4_lut (.I0(n15_c), .I1(n20_adj_5423), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n1962));
    defparam i10_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_adj_1099 (.I0(byte_transmit_counter_c[4]), .I1(byte_transmit_counter_c[3]), 
            .I2(GND_net), .I3(GND_net), .O(n4_c));   // verilog/coms.v(217[11:56])
    defparam i1_2_lut_adj_1099.LUT_INIT = 16'h8888;
    SB_LUT4 i46290_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n62976));   // verilog/coms.v(158[12:15])
    defparam i46290_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i17174_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[3] [2]), 
            .I3(\data_in_frame[19] [2]), .O(n4940[2]));   // verilog/coms.v(148[4] 304[11])
    defparam i17174_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i46342_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n62975));   // verilog/coms.v(158[12:15])
    defparam i46342_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESS data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5411), .S(n55382));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_6_lut  (.I0(n63058), .I1(n27843), 
            .I2(\FRAME_MATCHER.i[4] ), .I3(n49176), .O(n27576)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_6_lut .LUT_INIT = 16'h8BB8;
    SB_LUT4 i2_4_lut_adj_1100 (.I0(byte_transmit_counter[0]), .I1(n4_c), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n58202));   // verilog/coms.v(217[11:56])
    defparam i2_4_lut_adj_1100.LUT_INIT = 16'hc8c0;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_6  (.CI(n49176), .I0(n27843), .I1(\FRAME_MATCHER.i[4] ), 
            .CO(n49177));
    SB_LUT4 n66747_bdd_4_lut (.I0(n66747), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[16] [3]), .I3(byte_transmit_counter[1]), 
            .O(n66750));
    defparam n66747_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_5_lut  (.I0(n63079), .I1(n27843), 
            .I2(\FRAME_MATCHER.i[3] ), .I3(n49175), .O(n27574)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_5_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_5  (.CI(n49175), .I0(n27843), .I1(\FRAME_MATCHER.i[3] ), 
            .CO(n49176));
    SB_LUT4 i46265_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n62970));   // verilog/coms.v(158[12:15])
    defparam i46265_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_4_lut  (.I0(n63080), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n49174), .O(n27572)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_4_lut .LUT_INIT = 16'h8BB8;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_4  (.CI(n49174), .I0(n27843), .I1(\FRAME_MATCHER.i [2]), 
            .CO(n49175));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_3_lut  (.I0(n63103), .I1(n27843), 
            .I2(\FRAME_MATCHER.i [1]), .I3(n49173), .O(n27570)) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_3_lut .LUT_INIT = 16'h8BB8;
    SB_DFFE data_in_frame_0___i127 (.Q(\data_in_frame[15] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29362));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5410), .S(n55381));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i46291_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n62967));   // verilog/coms.v(158[12:15])
    defparam i46291_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_3  (.CI(n49173), .I0(n27843), .I1(\FRAME_MATCHER.i [1]), 
            .CO(n49174));
    SB_LUT4 \FRAME_MATCHER.i_2043_add_4_2_lut  (.I0(GND_net), .I1(n161), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \FRAME_MATCHER.i_2043_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \FRAME_MATCHER.i_2043_add_4_2  (.CI(GND_net), .I0(n161), .I1(\FRAME_MATCHER.i[0] ), 
            .CO(n49173));
    SB_LUT4 i46345_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n62966));   // verilog/coms.v(158[12:15])
    defparam i46345_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_1087_i4_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[3][3] ), 
            .I3(\data_in_frame[19]_c [3]), .O(n4940[3]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i4_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i2_3_lut (.I0(\r_SM_Main_2__N_3545[0] ), .I1(n53), .I2(tx_active), 
            .I3(GND_net), .O(n39951));
    defparam i2_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i46492_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n62963));   // verilog/coms.v(158[12:15])
    defparam i46492_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i366_2_lut (.I0(n1962), .I1(n1959), .I2(GND_net), .I3(GND_net), 
            .O(n1963));   // verilog/coms.v(142[4] 144[7])
    defparam i366_2_lut.LUT_INIT = 16'h8888;
    SB_DFFE data_in_frame_0___i126 (.Q(\data_in_frame[15] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29359));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), .I2(\data_in[1] [1]), 
            .I3(\data_in[0] [4]), .O(n10_adj_5424));
    defparam i4_4_lut.LUT_INIT = 16'hfdff;
    SB_DFFE data_in_frame_0___i125 (.Q(\data_in_frame[15] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29356));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i124 (.Q(\data_in_frame[15] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29353));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i53 (.Q(\data_in_frame[6] [4]), .C(clk16MHz), 
           .D(n29015));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut (.I0(\data_in[3] [4]), .I1(n10_adj_5424), .I2(\data_in[2] [7]), 
            .I3(GND_net), .O(n25223));
    defparam i5_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1101 (.I0(\data_in[0] [1]), .I1(\data_in[1] [2]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16));
    defparam i6_4_lut_adj_1101.LUT_INIT = 16'hfffe;
    SB_LUT4 i46229_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n62959));   // verilog/coms.v(158[12:15])
    defparam i46229_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i46243_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n62958));   // verilog/coms.v(158[12:15])
    defparam i46243_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i18809_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[3] [4]), 
            .I3(\data_in_frame[19]_c [4]), .O(n4940[4]));   // verilog/coms.v(148[4] 304[11])
    defparam i18809_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 i7_4_lut_adj_1102 (.I0(\data_in[1] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [3]), .O(n17));
    defparam i7_4_lut_adj_1102.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1103 (.I0(n17), .I1(\data_in[3] [7]), .I2(n16), 
            .I3(\data_in[2] [6]), .O(n25127));
    defparam i9_4_lut_adj_1103.LUT_INIT = 16'hfbff;
    SB_LUT4 i5_3_lut_adj_1104 (.I0(\data_in[1] [0]), .I1(\data_in[2] [4]), 
            .I2(\data_in[3] [0]), .I3(GND_net), .O(n14_adj_5425));
    defparam i5_3_lut_adj_1104.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1105 (.I0(\data_in[1] [4]), .I1(\data_in[0] [6]), 
            .I2(n25223), .I3(\data_in[1] [5]), .O(n15_adj_5426));
    defparam i6_4_lut_adj_1105.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_1106 (.I0(n15_adj_5426), .I1(\data_in[2] [2]), 
            .I2(n14_adj_5425), .I3(\data_in[0] [3]), .O(n24976));
    defparam i8_4_lut_adj_1106.LUT_INIT = 16'hfbff;
    SB_DFFE data_in_frame_0___i123 (.Q(\data_in_frame[15] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29349));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1107 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n24976), .O(n16_adj_5427));
    defparam i6_4_lut_adj_1107.LUT_INIT = 16'hffef;
    SB_DFFESS data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5392), .S(n55380));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i46359_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n62946));   // verilog/coms.v(158[12:15])
    defparam i46359_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i11999_1_lut (.I0(n3484), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n27843));   // verilog/coms.v(148[4] 304[11])
    defparam i11999_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE data_in_frame_0___i122 (.Q(\data_in_frame[15] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29346));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5390), .S(n55379));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i121 (.Q(\data_in_frame[15] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29343));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1087_i6_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[3][5] ), 
            .I3(\data_in_frame[19]_c [5]), .O(n4940[5]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i6_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFFE data_in_frame_0___i120 (.Q(\data_in_frame[14] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29340));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i7_4_lut_adj_1108 (.I0(n25127), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [1]), .O(n17_adj_5428));
    defparam i7_4_lut_adj_1108.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1109 (.I0(n17_adj_5428), .I1(\data_in[3] [5]), 
            .I2(n16_adj_5427), .I3(\data_in[3] [3]), .O(n1965));
    defparam i9_4_lut_adj_1109.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_adj_1110 (.I0(\FRAME_MATCHER.i_31__N_2513 ), .I1(Kp_23__N_1748), 
            .I2(GND_net), .I3(GND_net), .O(n32100));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1110.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1111 (.I0(n1965), .I1(\FRAME_MATCHER.i_31__N_2507 ), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5429));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_adj_1111.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1112 (.I0(\FRAME_MATCHER.i_31__N_2511 ), .I1(n1963), 
            .I2(n39951), .I3(n4_adj_5429), .O(n6_c));   // verilog/coms.v(148[4] 304[11])
    defparam i2_4_lut_adj_1112.LUT_INIT = 16'heca0;
    SB_LUT4 i3_4_lut_adj_1113 (.I0(n32100), .I1(n6_c), .I2(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I3(\FRAME_MATCHER.i_31__N_2509 ), .O(n67128));   // verilog/coms.v(148[4] 304[11])
    defparam i3_4_lut_adj_1113.LUT_INIT = 16'hefee;
    SB_LUT4 mux_1087_i7_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[3][6] ), 
            .I3(\data_in_frame[19]_c [6]), .O(n4940[6]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i7_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i21_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[1] [4]), 
            .I3(\data_in_frame[17][4] ), .O(n4940[20]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i21_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_787_Select_55_i2_4_lut (.I0(\data_out_frame[6] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[23] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5418));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_55_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14021_3_lut_4_lut (.I0(n8_adj_5430), .I1(n55507), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n29866));
    defparam i14021_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14024_3_lut_4_lut (.I0(n8_adj_5430), .I1(n55507), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n29869));
    defparam i14024_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14045_3_lut_4_lut (.I0(n8), .I1(n55507), .I2(rx_data[6]), 
            .I3(\data_in_frame[2]_c [6]), .O(n29890));
    defparam i14045_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14048_3_lut_4_lut (.I0(n8), .I1(n55507), .I2(rx_data[7]), 
            .I3(\data_in_frame[2]_c [7]), .O(n29893));
    defparam i14048_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1087_i22_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[1] [5]), 
            .I3(\data_in_frame[17][5] ), .O(n4940[21]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i22_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i23_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[1] [6]), 
            .I3(\data_in_frame[17]_c [6]), .O(n4940[22]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i23_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i24_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[1] [7]), 
            .I3(\data_in_frame[17] [7]), .O(n4940[23]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i24_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i1_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[3][0] ), 
            .I3(\data_in_frame[19][0] ), .O(n4940[0]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i1_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i9_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[2] [0]), 
            .I3(\data_in_frame[18] [0]), .O(n4940[8]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i9_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFFE data_in_frame_0___i119 (.Q(\data_in_frame[14][6] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29337));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 add_1194_9_lut (.I0(n55427), .I1(\byte_transmit_counter[7] ), 
            .I2(GND_net), .I3(n48382), .O(n55435)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_9_lut.LUT_INIT = 16'h8228;
    SB_DFFE data_in_frame_0___i118 (.Q(\data_in_frame[14] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29334));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1087_i10_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[2]_c [1]), 
            .I3(\data_in_frame[18] [1]), .O(n4940[9]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i10_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 add_1194_8_lut (.I0(n55427), .I1(\byte_transmit_counter[6] ), 
            .I2(GND_net), .I3(n48381), .O(n55433)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_8_lut.LUT_INIT = 16'h8228;
    SB_DFFE data_in_frame_0___i117 (.Q(\data_in_frame[14] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29331));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1087_i11_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[2]_c [2]), 
            .I3(\data_in_frame[18] [2]), .O(n4940[10]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i11_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 mux_1087_i12_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[2]_c [3]), 
            .I3(\data_in_frame[18] [3]), .O(n4940[11]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i12_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFFE data_in_frame_0___i116 (.Q(\data_in_frame[14] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29328));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i115 (.Q(\data_in_frame[14] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29325));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i114 (.Q(\data_in_frame[14] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29322));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i113 (.Q(\data_in_frame[14] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29319));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1194_8 (.CI(n48381), .I0(\byte_transmit_counter[6] ), .I1(GND_net), 
            .CO(n48382));
    SB_LUT4 add_1194_7_lut (.I0(n55427), .I1(\byte_transmit_counter[5] ), 
            .I2(GND_net), .I3(n48380), .O(n55434)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1194_7 (.CI(n48380), .I0(\byte_transmit_counter[5] ), .I1(GND_net), 
            .CO(n48381));
    SB_DFFE data_in_frame_0___i112 (.Q(\data_in_frame[13] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29316));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i111 (.Q(\data_in_frame[13] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29313));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i54 (.Q(\data_in_frame[6]_c [5]), .C(clk16MHz), 
           .D(n29312));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i110 (.Q(\data_in_frame[13] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29309));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1087_i13_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[2]_c [4]), 
            .I3(\data_in_frame[18] [4]), .O(n4940[12]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i13_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 add_1194_6_lut (.I0(n55427), .I1(byte_transmit_counter_c[4]), 
            .I2(GND_net), .I3(n48379), .O(n55432)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_6_lut.LUT_INIT = 16'h8228;
    SB_DFFE data_in_frame_0___i109 (.Q(\data_in_frame[13] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29306));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i108 (.Q(\data_in_frame[13] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29303));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i107 (.Q(\data_in_frame[13] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29300));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1194_6 (.CI(n48379), .I0(byte_transmit_counter_c[4]), .I1(GND_net), 
            .CO(n48380));
    SB_DFFE data_in_frame_0___i106 (.Q(\data_in_frame[13] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29297));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5431), .S(n55378));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i105 (.Q(\data_in_frame[13] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29294));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1087_i14_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[2]_c [5]), 
            .I3(\data_in_frame[18] [5]), .O(n4940[13]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i14_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFFE data_in_frame_0___i104 (.Q(\data_in_frame[12] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29291));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i103 (.Q(\data_in_frame[12] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29288));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i102 (.Q(\data_in_frame[12] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29285));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i101 (.Q(\data_in_frame[12] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29282));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i55 (.Q(\data_in_frame[6][6] ), .C(clk16MHz), 
           .D(n29021));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i100 (.Q(\data_in_frame[12] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29278));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i99 (.Q(\data_in_frame[12] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29275));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i98 (.Q(\data_in_frame[12] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29272));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i97 (.Q(\data_in_frame[12] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29269));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i96 (.Q(\data_in_frame[11] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29266));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1087_i15_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[2]_c [6]), 
            .I3(\data_in_frame[18] [6]), .O(n4940[14]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i15_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFFE data_in_frame_0___i95 (.Q(\data_in_frame[11] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29263));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i56 (.Q(\data_in_frame[6][7] ), .C(clk16MHz), 
           .D(n29024));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i57 (.Q(\data_in_frame[7] [0]), .C(clk16MHz), 
           .D(n54823));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i94 (.Q(\data_in_frame[11] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29258));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i93 (.Q(\data_in_frame[11] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29255));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i92 (.Q(\data_in_frame[11] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29252));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5432), .S(n55377));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i91 (.Q(\data_in_frame[11] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29249));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i90 (.Q(\data_in_frame[11] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29246));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 add_1194_5_lut (.I0(n55427), .I1(byte_transmit_counter_c[3]), 
            .I2(GND_net), .I3(n48378), .O(n55429)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mux_1087_i16_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[2]_c [7]), 
            .I3(\data_in_frame[18] [7]), .O(n4940[15]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i16_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFFE data_in_frame_0___i89 (.Q(\data_in_frame[11] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29243));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i88 (.Q(\data_in_frame[10] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29240));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i87 (.Q(\data_in_frame[10] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29237));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i86 (.Q(\data_in_frame[10] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29234));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1087_i17_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[1] [0]), 
            .I3(\data_in_frame[17][0] ), .O(n4940[16]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i17_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_LUT4 select_787_Select_223_i3_4_lut (.I0(\data_out_frame[25] [6]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n55844), .I3(\data_out_frame[25] [5]), 
            .O(n3_adj_5409));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_223_i3_4_lut.LUT_INIT = 16'h4884;
    SB_DFFE data_in_frame_0___i85 (.Q(\data_in_frame[10] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29231));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i84 (.Q(\data_in_frame[10] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29228));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1087_i18_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[1]_c [1]), 
            .I3(\data_in_frame[17][1] ), .O(n4940[17]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i18_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFFE data_in_frame_0___i83 (.Q(\data_in_frame[10] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29225));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i82 (.Q(\data_in_frame[10] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29222));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i81 (.Q(\data_in_frame[10] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29219));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i80 (.Q(\data_in_frame[9] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29216));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i79 (.Q(\data_in_frame[9] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29213));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i78 (.Q(\data_in_frame[9] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29210));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i77 (.Q(\data_in_frame[9] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29207));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i76 (.Q(\data_in_frame[9] [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29204));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i75 (.Q(\data_in_frame[9] [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29201));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i31776_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[1]_c [2]), 
            .I3(\data_in_frame[17][2] ), .O(n4940[18]));   // verilog/coms.v(148[4] 304[11])
    defparam i31776_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFFE data_in_frame_0___i74 (.Q(\data_in_frame[9] [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29198));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i73 (.Q(\data_in_frame[9] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29195));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i72 (.Q(\data_in_frame[8] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29192));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i71 (.Q(\data_in_frame[8] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29189));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i70 (.Q(\data_in_frame[8] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29186));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i58 (.Q(\data_in_frame[7][1] ), .C(clk16MHz), 
           .D(n29030));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1087_i20_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[1]_c [3]), 
            .I3(\data_in_frame[17][3] ), .O(n4940[19]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i20_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFF data_in_frame_0___i59 (.Q(\data_in_frame[7][2] ), .C(clk16MHz), 
           .D(n29033));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i60 (.Q(\data_in_frame[7] [3]), .C(clk16MHz), 
           .D(n54827));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i23 (.Q(setpoint[23]), .C(clk16MHz), .E(n27322), 
            .D(n4940[23]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49646 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n66717));
    defparam byte_transmit_counter_0__bdd_4_lut_49646.LUT_INIT = 16'he4aa;
    SB_DFFER setpoint_i0_i22 (.Q(setpoint[22]), .C(clk16MHz), .E(n27322), 
            .D(n4940[22]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i21 (.Q(setpoint[21]), .C(clk16MHz), .E(n27322), 
            .D(n4940[21]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i20 (.Q(setpoint[20]), .C(clk16MHz), .E(n27322), 
            .D(n4940[20]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i19 (.Q(setpoint[19]), .C(clk16MHz), .E(n27322), 
            .D(n4940[19]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i18 (.Q(setpoint[18]), .C(clk16MHz), .E(n27322), 
            .D(n4940[18]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i17 (.Q(setpoint[17]), .C(clk16MHz), .E(n27322), 
            .D(n4940[17]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i16 (.Q(setpoint[16]), .C(clk16MHz), .E(n27322), 
            .D(n4940[16]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i61 (.Q(\data_in_frame[7][4] ), .C(clk16MHz), 
           .D(n29042));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 mux_1087_i8_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[3][7] ), 
            .I3(\data_in_frame[19]_c [7]), .O(n4940[7]));   // verilog/coms.v(148[4] 304[11])
    defparam mux_1087_i8_3_lut_4_lut.LUT_INIT = 16'hf870;
    SB_DFF data_in_frame_0___i62 (.Q(\data_in_frame[7][5] ), .C(clk16MHz), 
           .D(n29045));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i63 (.Q(\data_in_frame[7][6] ), .C(clk16MHz), 
           .D(n29048));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i15 (.Q(setpoint[15]), .C(clk16MHz), .E(n27322), 
            .D(n4940[15]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i14 (.Q(setpoint[14]), .C(clk16MHz), .E(n27322), 
            .D(n4940[14]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i13 (.Q(setpoint[13]), .C(clk16MHz), .E(n27322), 
            .D(n4940[13]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i12 (.Q(setpoint[12]), .C(clk16MHz), .E(n27322), 
            .D(n4940[12]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i11 (.Q(setpoint[11]), .C(clk16MHz), .E(n27322), 
            .D(n4940[11]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i10 (.Q(setpoint[10]), .C(clk16MHz), .E(n27322), 
            .D(n4940[10]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i9 (.Q(setpoint[9]), .C(clk16MHz), .E(n27322), 
            .D(n4940[9]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i8 (.Q(setpoint[8]), .C(clk16MHz), .E(n27322), 
            .D(n4940[8]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i7 (.Q(setpoint[7]), .C(clk16MHz), .E(n27322), 
            .D(n4940[7]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i6 (.Q(setpoint[6]), .C(clk16MHz), .E(n27322), 
            .D(n4940[6]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i5 (.Q(setpoint[5]), .C(clk16MHz), .E(n27322), 
            .D(n4940[5]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i64 (.Q(\data_in_frame[7][7] ), .C(clk16MHz), 
           .D(n29051));   // verilog/coms.v(130[12] 305[6])
    SB_CARRY add_1194_5 (.CI(n48378), .I0(byte_transmit_counter_c[3]), .I1(GND_net), 
            .CO(n48379));
    SB_DFF data_in_frame_0___i65 (.Q(\data_in_frame[8] [0]), .C(clk16MHz), 
           .D(n29054));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i66 (.Q(\data_in_frame[8] [1]), .C(clk16MHz), 
           .D(n29057));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i4 (.Q(setpoint[4]), .C(clk16MHz), .E(n27322), 
            .D(n4940[4]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i3 (.Q(setpoint[3]), .C(clk16MHz), .E(n27322), 
            .D(n4940[3]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i2 (.Q(setpoint[2]), .C(clk16MHz), .E(n27322), 
            .D(n4940[2]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFER setpoint_i0_i1 (.Q(setpoint[1]), .C(clk16MHz), .E(n27322), 
            .D(n4940[1]), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS \FRAME_MATCHER.state_FSM_i9  (.Q(\FRAME_MATCHER.i_31__N_2507 ), 
            .C(clk16MHz), .D(n67128), .S(reset));   // verilog/coms.v(148[4] 304[11])
    SB_LUT4 n66717_bdd_4_lut (.I0(n66717), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n66720));
    defparam n66717_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_49686 (.I0(byte_transmit_counter[1]), 
            .I1(\data_out_frame[25] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[0]), .O(n66711));
    defparam byte_transmit_counter_1__bdd_4_lut_49686.LUT_INIT = 16'he4aa;
    SB_LUT4 add_1194_4_lut (.I0(n55427), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n48377), .O(n55430)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 n66711_bdd_4_lut (.I0(n66711), .I1(\data_out_frame[26] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[0]), 
            .O(n66714));
    defparam n66711_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFR \FRAME_MATCHER.state_FSM_i8  (.Q(\FRAME_MATCHER.i_31__N_2508 ), 
            .C(clk16MHz), .D(n26634), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i7  (.Q(\FRAME_MATCHER.i_31__N_2509 ), 
            .C(clk16MHz), .D(n2056), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i6  (.Q(\FRAME_MATCHER.state[3] ), .C(clk16MHz), 
            .D(n2057), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i5  (.Q(\FRAME_MATCHER.i_31__N_2511 ), 
            .C(clk16MHz), .D(n20746), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i4  (.Q(\FRAME_MATCHER.i_31__N_2512 ), 
            .C(clk16MHz), .D(n54455), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i3  (.Q(\FRAME_MATCHER.i_31__N_2513 ), 
            .C(clk16MHz), .D(n2068), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFR \FRAME_MATCHER.state_FSM_i2  (.Q(\FRAME_MATCHER.i_31__N_2514 ), 
            .C(clk16MHz), .D(n26637), .R(reset));   // verilog/coms.v(148[4] 304[11])
    SB_DFFESS data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5419), .S(n55302));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49621 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n66699));
    defparam byte_transmit_counter_0__bdd_4_lut_49621.LUT_INIT = 16'he4aa;
    SB_LUT4 n66699_bdd_4_lut (.I0(n66699), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n66702));
    defparam n66699_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0___i67 (.Q(\data_in_frame[8] [2]), .C(clk16MHz), 
           .D(n15_adj_5433));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i68 (.Q(\data_in_frame[8] [3]), .C(clk16MHz), 
           .D(n29160));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i69 (.Q(\data_in_frame[8] [4]), .C(clk16MHz), 
           .D(n15_adj_5434));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i39383_3_lut_4_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(n7), .I2(n56366), 
            .I3(reset), .O(n27934));   // verilog/coms.v(157[7:23])
    defparam i39383_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 select_787_Select_222_i3_4_lut (.I0(\data_out_frame[23] [4]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n8_adj_5435), .I3(n56162), 
            .O(n3_adj_5408));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_222_i3_4_lut.LUT_INIT = 16'h4884;
    SB_CARRY add_1194_4 (.CI(n48377), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n48378));
    SB_LUT4 add_1194_3_lut (.I0(n55427), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n48376), .O(n55431)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1114 (.I0(\data_in_frame[19]_c [7]), .I1(\data_in_frame[15] [6]), 
            .I2(\data_in_frame[20] [0]), .I3(\data_in_frame[20] [1]), .O(n59598));
    defparam i1_4_lut_adj_1114.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1115 (.I0(n51148), .I1(n59598), .I2(\data_in_frame[20] [3]), 
            .I3(\data_in_frame[20] [2]), .O(n59602));
    defparam i1_4_lut_adj_1115.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1116 (.I0(n50620), .I1(n56050), .I2(n56171), 
            .I3(n59602), .O(n59608));
    defparam i1_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1117 (.I0(n51168), .I1(n50179), .I2(n51243), 
            .I3(n59608), .O(n59614));
    defparam i1_4_lut_adj_1117.LUT_INIT = 16'h6996;
    SB_CARRY add_1194_3 (.CI(n48376), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n48377));
    SB_LUT4 add_1194_2_lut (.I0(n55427), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3416), .I3(GND_net), .O(n55428)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1194_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i49202_3_lut (.I0(rx_data[3]), .I1(\data_in_frame[7] [3]), .I2(n27906), 
            .I3(GND_net), .O(n54827));   // verilog/coms.v(94[13:20])
    defparam i49202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1118 (.I0(n56246), .I1(n55975), .I2(n56168), 
            .I3(n59614), .O(n59620));
    defparam i1_4_lut_adj_1118.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1119 (.I0(n55672), .I1(n51239), .I2(n51173), 
            .I3(n59620), .O(n59626));
    defparam i1_4_lut_adj_1119.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1120 (.I0(n55633), .I1(\data_in_frame[21][1] ), 
            .I2(\data_in_frame[21] [7]), .I3(n55815), .O(n59462));
    defparam i1_4_lut_adj_1120.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1121 (.I0(n50305), .I1(n55946), .I2(n55932), 
            .I3(n59626), .O(n57892));
    defparam i1_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1122 (.I0(n50370), .I1(n57892), .I2(n59462), 
            .I3(n50368), .O(n55892));
    defparam i1_4_lut_adj_1122.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1123 (.I0(n57445), .I1(n51150), .I2(GND_net), 
            .I3(GND_net), .O(n51239));
    defparam i1_2_lut_adj_1123.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1124 (.I0(n55972), .I1(\data_in_frame[21]_c [6]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5436));
    defparam i1_2_lut_adj_1124.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1125 (.I0(\data_in_frame[19]_c [5]), .I1(n4_adj_5436), 
            .I2(n51239), .I3(n57531), .O(n55633));
    defparam i2_4_lut_adj_1125.LUT_INIT = 16'h6996;
    SB_CARRY add_1194_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3416), 
            .CO(n48376));
    SB_LUT4 i1_4_lut_adj_1126 (.I0(\data_in_frame[15] [2]), .I1(\data_in_frame[17][0] ), 
            .I2(\data_in_frame[15] [4]), .I3(\data_in_frame[16] [0]), .O(n59424));
    defparam i1_4_lut_adj_1126.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1127 (.I0(\data_in_frame[15] [0]), .I1(\data_in_frame[16] [4]), 
            .I2(\data_in_frame[10] [6]), .I3(\data_in_frame[13] [6]), .O(n59426));
    defparam i1_4_lut_adj_1127.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1128 (.I0(\data_in_frame[16] [6]), .I1(\data_in_frame[14] [7]), 
            .I2(\data_in_frame[15] [6]), .I3(\data_in_frame[12] [7]), .O(n59428));
    defparam i1_4_lut_adj_1128.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut (.I0(n59426), .I1(Kp_23__N_1389), .I2(n59424), .I3(GND_net), 
            .O(n59434));
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1129 (.I0(n26257), .I1(n59434), .I2(n55829), 
            .I3(n59428), .O(n59438));
    defparam i1_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1130 (.I0(n25895), .I1(n56047), .I2(Kp_23__N_1067), 
            .I3(n59438), .O(n59444));
    defparam i1_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1131 (.I0(n25345), .I1(n51414), .I2(n55819), 
            .I3(n59444), .O(n59450));
    defparam i1_4_lut_adj_1131.LUT_INIT = 16'h9669;
    SB_DFFESS data_out_frame_0___i3 (.Q(\data_out_frame[0][2] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5347), .S(n55418));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5346), .S(n55417));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5345), .S(n55416));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i9 (.Q(\data_out_frame[1][0] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5344), .S(n55415));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i10 (.Q(\data_out_frame[1][1] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5341), .S(n55414));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i12 (.Q(\data_out_frame[1][3] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5340), .S(n55413));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i14 (.Q(\data_out_frame[1][5] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5339), .S(n55412));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i15 (.Q(\data_out_frame[1][6] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5330), .S(n55411));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i16 (.Q(\data_out_frame[1][7] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5325), .S(n55410));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5317), .S(n55376));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i67 (.Q(\data_out_frame[8][2] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5314), .S(n55303));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i68 (.Q(\data_out_frame[8][3] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5313), .S(n55375));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i69 (.Q(\data_out_frame[8][4] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5312), .S(n55374));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i70 (.Q(\data_out_frame[8][5] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5307), .S(n55373));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i71 (.Q(\data_out_frame[8][6] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5304), .S(n55372));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i72 (.Q(\data_out_frame[8][7] ), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5299), .S(n55371));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5292), .S(n55370));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5437), .S(n55369));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5438), .S(n55368));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5439), .S(n55367));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5440), .S(n55366));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5441), .S(n55365));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5442), .S(n55364));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5443), .S(n55363));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5444), .S(n55362));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5445), .S(n55361));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5446), .S(n55360));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5447), .S(n55359));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5448), .S(n55358));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5449), .S(n55357));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk16MHz), 
            .E(n2882), .D(n11), .S(n55356));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5450), .S(n55355));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5451), .S(n55354));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5452), .S(n55353));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5453), .S(n55352));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5454), .S(n55351));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5455), .S(n55350));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5456), .S(n55349));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5457), .S(n55348));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5458), .S(n55347));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5459), .S(n55346));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5460), .S(n55345));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5461), .S(n55344));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5462), .S(n55343));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5463), .S(n55342));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5464), .S(n55341));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5465), .S(n55340));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5466), .S(n55339));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5467), .S(n55338));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5468), .S(n55337));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5469), .S(n55336));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5470), .S(n55335));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5471), .S(n55334));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5472), .S(n55333));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5473), .S(n55332));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5474), .S(n55331));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5475), .S(n55330));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5476), .S(n55329));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5477), .S(n55328));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5478), .S(n55327));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5479), .S(n55326));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5480), .S(n55325));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5481), .S(n55305));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5482), .S(n55324));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk16MHz), .D(n29095));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5483), .S(n55323));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk16MHz), .D(n29094));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5484), .S(n55322));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk16MHz), .D(n29093));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5485), .S(n55321));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk16MHz), .D(n29092));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5486), .S(n55320));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk16MHz), .D(n29091));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk16MHz), .D(n29090));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk16MHz), .D(n29089));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk16MHz), .D(n29088));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5487), .S(n55319));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk16MHz), .D(n29087));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk16MHz), .D(n29086));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk16MHz), .D(n29085));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5488), .S(n55318));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk16MHz), .D(n29084));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk16MHz), .D(n29083));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk16MHz), .D(n29082));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5489), .S(n55317));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk16MHz), .D(n29081));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk16MHz), .D(n29080));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk16MHz), .D(n29079));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5490), .S(n55304));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk16MHz), .D(n29078));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk16MHz), .D(n29077));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk16MHz), .D(n29076));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5491), .S(n55316));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk16MHz), .D(n29075));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk16MHz), .D(n29074));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk16MHz), .D(n29073));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk16MHz), .D(n29072));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5492), .S(n55315));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk16MHz), .D(n29071));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk16MHz), .D(n29070));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk16MHz), .D(n29069));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5493), .S(n55314));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk16MHz), .D(n29068));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk16MHz), .D(n29067));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk16MHz), .D(n29066));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5494), .S(n55313));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk16MHz), .D(n29065));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5495), .S(n55312));   // verilog/coms.v(130[12] 305[6])
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_4012  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk16MHz), .D(n29061));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5496), .S(n55311));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5497), .S(n55310));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5498), .S(n55309));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5499), .S(n55308));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5500), .S(n55307));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5501), .S(n55306));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5502), .S(n55298));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5503), .S(n55297));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5504), .S(n55296));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1132 (.I0(n51173), .I1(n56181), .I2(n59450), 
            .I3(n56147), .O(Kp_23__N_1518));
    defparam i1_4_lut_adj_1132.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_25_i2_3_lut (.I0(\data_out_frame[3][1] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5298));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_25_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFFESS data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5505), .S(n55295));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_3_lut_4_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(n6_adj_5506), .I3(n25246), .O(n55606));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1133 (.I0(n50620), .I1(n55889), .I2(n59542), 
            .I3(n56159), .O(n59548));
    defparam i1_4_lut_adj_1133.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1134 (.I0(n50179), .I1(n56138), .I2(Kp_23__N_1518), 
            .I3(n59548), .O(n55946));
    defparam i1_4_lut_adj_1134.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_adj_1135 (.I0(\data_in_frame[18] [5]), .I1(n51243), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5507));
    defparam i2_2_lut_adj_1135.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1136 (.I0(\data_in_frame[3][5] ), .I1(\data_in_frame[5] [7]), 
            .I2(\data_in_frame[1]_c [3]), .I3(GND_net), .O(n55695));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1136.LUT_INIT = 16'h9696;
    SB_DFFR \FRAME_MATCHER.i_2043__i0  (.Q(\FRAME_MATCHER.i[0] ), .C(clk16MHz), 
            .D(n27541), .R(reset));   // verilog/coms.v(158[12:15])
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[3][5] ), .I1(\data_in_frame[5] [7]), 
            .I2(n56035), .I3(Kp_23__N_843), .O(n25500));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFESS LED_4014 (.Q(LED_c), .C(clk16MHz), .E(n2882), .D(n5_adj_5422), 
            .S(n28428));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i6_4_lut_adj_1137 (.I0(n56159), .I1(n26277), .I2(Kp_23__N_1518), 
            .I3(n24707), .O(n14_adj_5508));
    defparam i6_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1138 (.I0(n55946), .I1(n14_adj_5508), .I2(n10_adj_5507), 
            .I3(\data_in_frame[20] [1]), .O(n55929));
    defparam i7_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1139 (.I0(\data_in_frame[16] [3]), .I1(n57567), 
            .I2(n56120), .I3(GND_net), .O(n26277));
    defparam i1_3_lut_adj_1139.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1140 (.I0(\data_in_frame[20] [5]), .I1(n26277), 
            .I2(\data_in_frame[20] [4]), .I3(GND_net), .O(n55672));
    defparam i2_3_lut_adj_1140.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1141 (.I0(n58144), .I1(n55985), .I2(GND_net), 
            .I3(GND_net), .O(n56181));
    defparam i1_2_lut_adj_1141.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1142 (.I0(n50393), .I1(n54275), .I2(n56156), 
            .I3(n55917), .O(n59470));
    defparam i1_4_lut_adj_1142.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1143 (.I0(n51206), .I1(n55772), .I2(n55613), 
            .I3(\data_in_frame[14][6] ), .O(n58097));
    defparam i3_4_lut_adj_1143.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1144 (.I0(n58097), .I1(n59470), .I2(n59538), 
            .I3(n55911), .O(n58144));
    defparam i1_4_lut_adj_1144.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1145 (.I0(n58144), .I1(\data_in_frame[19]_c [4]), 
            .I2(n57445), .I3(GND_net), .O(n57531));
    defparam i2_3_lut_adj_1145.LUT_INIT = 16'h9696;
    SB_DFFESS driver_enable_4015 (.Q(DE_c), .C(clk16MHz), .E(n2882), .D(n26520), 
            .S(n28387));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i5_3_lut_adj_1146 (.I0(n51247), .I1(n50907), .I2(n55757), 
            .I3(GND_net), .O(n14_adj_5509));
    defparam i5_3_lut_adj_1146.LUT_INIT = 16'h6969;
    SB_LUT4 i6_4_lut_adj_1147 (.I0(n56174), .I1(\data_in_frame[16] [1]), 
            .I2(n25895), .I3(n55978), .O(n15_adj_5510));
    defparam i6_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1148 (.I0(n15_adj_5510), .I1(\data_in_frame[13] [5]), 
            .I2(n14_adj_5509), .I3(\data_in_frame[13] [3]), .O(n57567));
    defparam i8_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_DFFESS tx_transmit_4011 (.Q(\r_SM_Main_2__N_3545[0] ), .C(clk16MHz), 
            .E(n2882), .D(n1_adj_5511), .S(n28384));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1149 (.I0(n51228), .I1(n55926), .I2(GND_net), 
            .I3(GND_net), .O(n51148));
    defparam i1_2_lut_adj_1149.LUT_INIT = 16'h9999;
    SB_LUT4 data_in_frame_17__7__I_0_4040_2_lut (.I0(\data_in_frame[17] [7]), 
            .I1(\data_in_frame[17]_c [6]), .I2(GND_net), .I3(GND_net), 
            .O(Kp_23__N_1389));   // verilog/coms.v(73[16:27])
    defparam data_in_frame_17__7__I_0_4040_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1150 (.I0(n7_adj_5512), .I1(n55978), .I2(n51359), 
            .I3(Kp_23__N_1389), .O(n56144));
    defparam i4_4_lut_adj_1150.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1151 (.I0(n55941), .I1(n55851), .I2(n25428), 
            .I3(n26257), .O(n56156));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_1151.LUT_INIT = 16'h6996;
    SB_DFFESS data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5513), .S(n55294));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_3_lut_adj_1152 (.I0(n56156), .I1(\data_in_frame[15] [3]), 
            .I2(n55621), .I3(GND_net), .O(n51414));
    defparam i2_3_lut_adj_1152.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1153 (.I0(n51359), .I1(n51414), .I2(\data_in_frame[17][5] ), 
            .I3(GND_net), .O(n50179));
    defparam i2_3_lut_adj_1153.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1154 (.I0(\data_in_frame[15] [3]), .I1(n51226), 
            .I2(\data_in_frame[17][4] ), .I3(GND_net), .O(n51150));
    defparam i2_3_lut_adj_1154.LUT_INIT = 16'h6969;
    SB_DFFESS byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk16MHz), 
            .E(n2882), .D(n1_adj_5514), .S(n55428));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1155 (.I0(n51256), .I1(n51228), .I2(GND_net), 
            .I3(GND_net), .O(n55917));
    defparam i1_2_lut_adj_1155.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1156 (.I0(\data_in_frame[12] [7]), .I1(n50317), 
            .I2(GND_net), .I3(GND_net), .O(n55851));
    defparam i1_2_lut_adj_1156.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1157 (.I0(n56117), .I1(n25428), .I2(\data_in_frame[13] [0]), 
            .I3(\data_in_frame[13] [2]), .O(n14_adj_5515));
    defparam i6_4_lut_adj_1157.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1158 (.I0(n25607), .I1(n14_adj_5515), .I2(n10_adj_5516), 
            .I3(\data_in_frame[12] [6]), .O(n51226));
    defparam i7_4_lut_adj_1158.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1159 (.I0(n55704), .I1(n50907), .I2(n51256), 
            .I3(\data_in_frame[14] [7]), .O(n55911));
    defparam i1_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1160 (.I0(n51226), .I1(n56147), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5517));
    defparam i1_2_lut_adj_1160.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1161 (.I0(\data_in_frame[17][3] ), .I1(n51168), 
            .I2(n55911), .I3(n6_adj_5517), .O(n57445));
    defparam i4_4_lut_adj_1161.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1162 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1]_c [1]), 
            .I2(n55867), .I3(\data_in_frame[1]_c [2]), .O(n57764));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i15_2_lut (.I0(n50317), .I1(n51228), .I2(GND_net), .I3(GND_net), 
            .O(n54275));
    defparam i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1163 (.I0(\data_in_frame[11] [2]), .I1(n25337), 
            .I2(n57296), .I3(\data_in_frame[8] [6]), .O(n55926));
    defparam i3_4_lut_adj_1163.LUT_INIT = 16'h9669;
    SB_LUT4 i9_3_lut_4_lut (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1]_c [1]), 
            .I2(n57981), .I3(\data_in_frame[1] [6]), .O(n26));   // verilog/coms.v(99[12:25])
    defparam i9_3_lut_4_lut.LUT_INIT = 16'h0900;
    SB_LUT4 i3_3_lut (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [2]), 
            .I2(n56117), .I3(GND_net), .O(n8_adj_5518));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1164 (.I0(\data_in_frame[15] [4]), .I1(n55926), 
            .I2(n8_adj_5518), .I3(n55941), .O(n51359));
    defparam i1_4_lut_adj_1164.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1165 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1]_c [1]), 
            .I2(\data_in_frame[3][3] ), .I3(GND_net), .O(n56041));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_3_lut_adj_1165.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1166 (.I0(\data_in_frame[15] [5]), .I1(n51168), 
            .I2(n51359), .I3(GND_net), .O(n25345));
    defparam i2_3_lut_adj_1166.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1167 (.I0(n50272), .I1(n50260), .I2(GND_net), 
            .I3(GND_net), .O(n24804));
    defparam i1_2_lut_adj_1167.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1168 (.I0(\data_in_frame[18] [5]), .I1(n25941), 
            .I2(\data_in_frame[16] [5]), .I3(n55648), .O(n55889));
    defparam i3_4_lut_adj_1168.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1169 (.I0(\data_in_frame[18] [6]), .I1(n56168), 
            .I2(n55889), .I3(n55819), .O(Kp_23__N_1607));
    defparam i3_4_lut_adj_1169.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1170 (.I0(n55596), .I1(\data_in_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5519));
    defparam i2_2_lut_adj_1170.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1171 (.I0(n55599), .I1(\data_in_frame[6][0] ), 
            .I2(Kp_23__N_875), .I3(\data_in_frame[9] [4]), .O(n14_adj_5520));
    defparam i6_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1172 (.I0(n51363), .I1(n14_adj_5520), .I2(n10_adj_5519), 
            .I3(Kp_23__N_1080), .O(n58210));
    defparam i7_4_lut_adj_1172.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1173 (.I0(n56085), .I1(n56264), .I2(n56261), 
            .I3(n56222), .O(n14_adj_5521));
    defparam i6_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut (.I0(n55665), .I1(n55787), .I2(n56204), .I3(n55698), 
            .O(n13));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1174 (.I0(n13), .I1(\data_in_frame[14] [2]), .I2(n14_adj_5521), 
            .I3(n58210), .O(n50260));
    defparam i2_4_lut_adj_1174.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1175 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n55613));
    defparam i1_2_lut_adj_1175.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1176 (.I0(\data_in_frame[16] [7]), .I1(n55772), 
            .I2(\data_in_frame[12] [5]), .I3(GND_net), .O(n58100));
    defparam i2_3_lut_adj_1176.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1177 (.I0(\data_in_frame[17][1] ), .I1(n55613), 
            .I2(n58100), .I3(n4_adj_5522), .O(n55985));
    defparam i1_4_lut_adj_1177.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1178 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[14] [5]), 
            .I2(n26424), .I3(GND_net), .O(n4_adj_5522));
    defparam i1_3_lut_adj_1178.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_adj_1179 (.I0(n4_adj_5522), .I1(n26055), .I2(\data_in_frame[12] [4]), 
            .I3(GND_net), .O(n50264));
    defparam i3_3_lut_adj_1179.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1180 (.I0(n25557), .I1(\data_in_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n55599));
    defparam i1_2_lut_adj_1180.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1181 (.I0(n56027), .I1(\data_in_frame[10] [1]), 
            .I2(n55599), .I3(GND_net), .O(n26424));
    defparam i2_3_lut_adj_1181.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1182 (.I0(\data_in_frame[14] [4]), .I1(n55938), 
            .I2(\data_in_frame[12] [2]), .I3(n58201), .O(n25941));
    defparam i3_4_lut_adj_1182.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1183 (.I0(n25941), .I1(\data_in_frame[16] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n55624));
    defparam i1_2_lut_adj_1183.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1184 (.I0(\data_in_frame[14] [3]), .I1(n26424), 
            .I2(n55569), .I3(\data_in_frame[9] [6]), .O(n55648));
    defparam i3_4_lut_adj_1184.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1185 (.I0(\data_in_frame[19][0] ), .I1(n50310), 
            .I2(n55775), .I3(GND_net), .O(n55968));
    defparam i1_3_lut_adj_1185.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1186 (.I0(n55968), .I1(\data_in_frame[21][2] ), 
            .I2(n25705), .I3(GND_net), .O(n55815));
    defparam i2_3_lut_adj_1186.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1187 (.I0(n32987), .I1(\data_in_frame[21][3] ), 
            .I2(n25705), .I3(GND_net), .O(n50370));
    defparam i2_3_lut_adj_1187.LUT_INIT = 16'h9696;
    SB_LUT4 i4_2_lut_adj_1188 (.I0(n25557), .I1(n50498), .I2(GND_net), 
            .I3(GND_net), .O(n18_adj_5523));   // verilog/coms.v(99[12:25])
    defparam i4_2_lut_adj_1188.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1189 (.I0(n56075), .I1(n56219), .I2(\data_in_frame[8] [4]), 
            .I3(n56004), .O(n24));   // verilog/coms.v(99[12:25])
    defparam i10_4_lut_adj_1189.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1190 (.I0(\data_in_frame[9] [6]), .I1(\data_in_frame[6] [3]), 
            .I2(Kp_23__N_699), .I3(\data_in_frame[11] [7]), .O(n22));   // verilog/coms.v(99[12:25])
    defparam i8_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut (.I0(\data_in_frame[12] [0]), .I1(n24), .I2(n18_adj_5523), 
            .I3(\data_in_frame[8] [3]), .O(n26_adj_5524));   // verilog/coms.v(99[12:25])
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(n51319), .I1(n26_adj_5524), .I2(n22), .I3(n25490), 
            .O(n56085));   // verilog/coms.v(99[12:25])
    defparam i13_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1191 (.I0(\data_in_frame[9] [0]), .I1(Kp_23__N_974), 
            .I2(\data_in_frame[9] [1]), .I3(GND_net), .O(n25337));
    defparam i2_3_lut_adj_1191.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1192 (.I0(\data_in_frame[8] [7]), .I1(n56237), 
            .I2(n56112), .I3(n51230), .O(n51228));
    defparam i3_4_lut_adj_1192.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_adj_1193 (.I0(n56085), .I1(n50366), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_5525));
    defparam i2_2_lut_adj_1193.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1194 (.I0(n56153), .I1(\data_in_frame[13] [7]), 
            .I2(n55721), .I3(n25337), .O(n14_adj_5526));
    defparam i6_4_lut_adj_1194.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1195 (.I0(\data_in_frame[14] [1]), .I1(n14_adj_5526), 
            .I2(n10_adj_5525), .I3(\data_in_frame[11] [5]), .O(n50272));
    defparam i7_4_lut_adj_1195.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut (.I0(n55681), .I1(\data_in_frame[8] [3]), .I2(n25500), 
            .I3(GND_net), .O(n26001));   // verilog/coms.v(78[16:43])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1196 (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n55829));
    defparam i1_2_lut_adj_1196.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1197 (.I0(n25428), .I1(n25514), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1067));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1197.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1198 (.I0(n51319), .I1(\data_in_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n51363));
    defparam i1_2_lut_adj_1198.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1199 (.I0(\data_in_frame[12] [1]), .I1(\data_in_frame[9] [5]), 
            .I2(\data_in_frame[11] [7]), .I3(GND_net), .O(n56264));
    defparam i2_3_lut_adj_1199.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1200 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n56219));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1200.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_156_i2_4_lut (.I0(\data_out_frame[19] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5297));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_156_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i4_4_lut_adj_1201 (.I0(n55732), .I1(n24777), .I2(\data_in_frame[10] [2]), 
            .I3(n55802), .O(n10_adj_5527));
    defparam i4_4_lut_adj_1201.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1202 (.I0(n56041), .I1(n56065), .I2(\data_in_frame[10] [3]), 
            .I3(n56035), .O(n12));   // verilog/coms.v(78[16:27])
    defparam i5_4_lut_adj_1202.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1203 (.I0(\data_in_frame[1]_c [2]), .I1(n12), .I2(n56219), 
            .I3(n55754), .O(n26055));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_1203.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1204 (.I0(\data_in_frame[10] [4]), .I1(n55760), 
            .I2(GND_net), .I3(GND_net), .O(n25607));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1204.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1205 (.I0(n25557), .I1(n56264), .I2(n26413), 
            .I3(\data_in_frame[12] [2]), .O(n55569));
    defparam i3_4_lut_adj_1205.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n55681), .I1(\data_in_frame[8] [3]), 
            .I2(\data_in_frame[8] [2]), .I3(n26406), .O(n55760));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1206 (.I0(n26055), .I1(n58201), .I2(GND_net), 
            .I3(GND_net), .O(n51206));
    defparam i1_2_lut_adj_1206.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_4_lut_adj_1207 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[4] [0]), 
            .I2(\data_in_frame[6] [1]), .I3(n25490), .O(n56035));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1208 (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n56204));
    defparam i1_2_lut_adj_1208.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_155_i2_4_lut (.I0(\data_out_frame[19] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5296));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_155_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1209 (.I0(\data_in_frame[10] [6]), .I1(n25514), 
            .I2(GND_net), .I3(GND_net), .O(n55941));
    defparam i1_2_lut_adj_1209.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1210 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[4] [0]), 
            .I2(\data_in_frame[4] [1]), .I3(\data_in_frame[3][6] ), .O(n56062));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1210.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_154_i2_4_lut (.I0(\data_out_frame[19] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5295));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_154_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i39375_3_lut_4_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(n7), .I2(n55515), 
            .I3(reset), .O(n27900));   // verilog/coms.v(157[7:23])
    defparam i39375_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1211 (.I0(n25514), .I1(n26001), .I2(\data_in_frame[10] [5]), 
            .I3(GND_net), .O(n26257));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1211.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49884 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(byte_transmit_counter[1]), .O(n66885));
    defparam byte_transmit_counter_0__bdd_4_lut_49884.LUT_INIT = 16'he4aa;
    SB_LUT4 n66885_bdd_4_lut (.I0(n66885), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(byte_transmit_counter[1]), 
            .O(n66888));
    defparam n66885_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1212 (.I0(\data_in_frame[12] [4]), .I1(n26257), 
            .I2(GND_net), .I3(GND_net), .O(n25439));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1212.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1213 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n59558));
    defparam i1_2_lut_adj_1213.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1214 (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[11] [4]), 
            .I2(\data_in_frame[12] [0]), .I3(\data_in_frame[11] [2]), .O(n59564));
    defparam i1_4_lut_adj_1214.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1215 (.I0(n59564), .I1(n56204), .I2(n59558), 
            .I3(\data_in_frame[12] [6]), .O(n59568));
    defparam i1_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1216 (.I0(n56027), .I1(n55941), .I2(n56237), 
            .I3(n59568), .O(n59574));
    defparam i1_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1217 (.I0(n59574), .I1(n50744), .I2(n25439), 
            .I3(n56112), .O(n59580));
    defparam i1_4_lut_adj_1217.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1218 (.I0(n51206), .I1(n55569), .I2(n59580), 
            .I3(n55684), .O(n59586));
    defparam i1_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1219 (.I0(n50498), .I1(n55652), .I2(n59586), 
            .I3(n55938), .O(n58045));
    defparam i1_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 i12088_3_lut_4_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(n7), .I2(n56366), 
            .I3(reset), .O(n27932));   // verilog/coms.v(157[7:23])
    defparam i12088_3_lut_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[0]_c [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[0] [7]), .I3(\data_in_frame[1] [4]), .O(n22_adj_5528));   // verilog/coms.v(73[16:27])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h9600;
    SB_LUT4 i1_2_lut_adj_1220 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n25541));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1220.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1221 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[13] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n55621));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1221.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49761 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(byte_transmit_counter[1]), .O(n66873));
    defparam byte_transmit_counter_0__bdd_4_lut_49761.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_adj_1222 (.I0(n55684), .I1(\data_in_frame[13] [0]), 
            .I2(n26055), .I3(GND_net), .O(n55644));
    defparam i2_3_lut_adj_1222.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1223 (.I0(n55621), .I1(n55730), .I2(n25541), 
            .I3(\data_in_frame[13] [5]), .O(n50393));   // verilog/coms.v(88[17:63])
    defparam i1_4_lut_adj_1223.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1224 (.I0(n7_adj_5529), .I1(\data_in_frame[11] [5]), 
            .I2(\data_in_frame[9] [4]), .I3(n56112), .O(n55704));
    defparam i4_4_lut_adj_1224.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1225 (.I0(\data_in_frame[0]_c [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[1]_c [1]), .I3(GND_net), .O(n23332));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1225.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1226 (.I0(\data_in_frame[0]_c [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[3][0] ), .I3(Kp_23__N_767), .O(n26166));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1227 (.I0(n56047), .I1(n58045), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5530));
    defparam i1_2_lut_adj_1227.LUT_INIT = 16'h9999;
    SB_LUT4 i2_4_lut_adj_1228 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [2]), 
            .I2(\data_in_frame[13] [1]), .I3(n4_adj_5530), .O(n55745));
    defparam i2_4_lut_adj_1228.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1229 (.I0(n55704), .I1(n50393), .I2(n55644), 
            .I3(GND_net), .O(n50907));   // verilog/coms.v(79[16:43])
    defparam i1_3_lut_adj_1229.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1230 (.I0(n57296), .I1(n26031), .I2(GND_net), 
            .I3(GND_net), .O(n51189));
    defparam i1_2_lut_adj_1230.LUT_INIT = 16'h9999;
    SB_DFF data_in_frame_0___i151 (.Q(\data_in_frame[18] [6]), .C(clk16MHz), 
           .D(n29437));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_3_lut_4_lut (.I0(\data_in_frame[3] [2]), .I1(n23332), .I2(\data_in_frame[5] [4]), 
            .I3(\data_in_frame[5] [5]), .O(n25321));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1231 (.I0(\data_in_frame[11] [6]), .I1(n50744), 
            .I2(n25282), .I3(n26031), .O(n55757));
    defparam i3_4_lut_adj_1231.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1232 (.I0(\data_in_frame[9] [3]), .I1(n55721), 
            .I2(\data_in_frame[11] [4]), .I3(GND_net), .O(n51256));
    defparam i2_3_lut_adj_1232.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_153_i2_4_lut (.I0(\data_out_frame[19] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5294));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_153_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1233 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n25282));
    defparam i1_2_lut_adj_1233.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1234 (.I0(\data_in_frame[3] [2]), .I1(n23332), 
            .I2(n25769), .I3(GND_net), .O(n6_adj_5531));
    defparam i1_2_lut_3_lut_adj_1234.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1235 (.I0(Kp_23__N_875), .I1(\data_in_frame[6] [4]), 
            .I2(n55689), .I3(GND_net), .O(Kp_23__N_974));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1235.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1236 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n25839));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_adj_1236.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_9__7__I_0_2_lut (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1085));   // verilog/coms.v(88[17:28])
    defparam data_in_frame_9__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1237 (.I0(Kp_23__N_843), .I1(n50366), .I2(\data_in_frame[3][5] ), 
            .I3(\data_in_frame[5] [6]), .O(n55802));
    defparam i1_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1238 (.I0(n50744), .I1(n25572), .I2(GND_net), 
            .I3(GND_net), .O(n55923));
    defparam i1_2_lut_adj_1238.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1239 (.I0(n25481), .I1(n55802), .I2(GND_net), 
            .I3(GND_net), .O(n51250));
    defparam i1_2_lut_adj_1239.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1240 (.I0(\data_in_frame[7][7] ), .I1(\data_in_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n55754));
    defparam i1_2_lut_adj_1240.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1241 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[1] [5]), 
            .I2(n55754), .I3(n23345), .O(n56075));
    defparam i3_4_lut_adj_1241.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_8__7__I_0_4031_2_lut (.I0(\data_in_frame[8] [7]), 
            .I1(\data_in_frame[8] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_699));   // verilog/coms.v(74[16:27])
    defparam data_in_frame_8__7__I_0_4031_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_152_i2_4_lut (.I0(\data_out_frame[19] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5293));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_152_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1242 (.I0(Kp_23__N_875), .I1(\data_in_frame[6] [4]), 
            .I2(\data_in_frame[8] [5]), .I3(n55808), .O(n25428));   // verilog/coms.v(78[16:43])
    defparam i2_3_lut_4_lut_adj_1242.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_61_i2_4_lut (.I0(\data_out_frame[7] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[13] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5432));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_61_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1243 (.I0(n25428), .I1(n24683), .I2(Kp_23__N_1080), 
            .I3(\data_in_frame[9] [0]), .O(n50498));
    defparam i1_4_lut_adj_1243.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1244 (.I0(n55732), .I1(Kp_23__N_974), .I2(n55760), 
            .I3(Kp_23__N_699), .O(n59476));
    defparam i1_4_lut_adj_1244.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i152 (.Q(\data_in_frame[18] [7]), .C(clk16MHz), 
           .D(n29440));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i153 (.Q(\data_in_frame[19][0] ), .C(clk16MHz), 
           .D(n29443));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i154 (.Q(\data_in_frame[19] [1]), .C(clk16MHz), 
           .D(n29446));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i25 (.Q(\data_in_frame[3][0] ), .C(clk16MHz), 
           .D(n28912));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i26 (.Q(\data_in_frame[3] [1]), .C(clk16MHz), 
           .D(n54807));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i155 (.Q(\data_in_frame[19] [2]), .C(clk16MHz), 
           .D(n54635));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i156 (.Q(\data_in_frame[19]_c [3]), .C(clk16MHz), 
           .D(n29453));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i157 (.Q(\data_in_frame[19]_c [4]), .C(clk16MHz), 
           .D(n54599));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i158 (.Q(\data_in_frame[19]_c [5]), .C(clk16MHz), 
           .D(n29459));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i159 (.Q(\data_in_frame[19]_c [6]), .C(clk16MHz), 
           .D(n29462));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i160 (.Q(\data_in_frame[19]_c [7]), .C(clk16MHz), 
           .D(n29465));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i161 (.Q(\data_in_frame[20] [0]), .C(clk16MHz), 
           .D(n29468));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i162 (.Q(\data_in_frame[20] [1]), .C(clk16MHz), 
           .D(n29911));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i163 (.Q(\data_in_frame[20] [2]), .C(clk16MHz), 
           .D(n29474));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i164 (.Q(\data_in_frame[20] [3]), .C(clk16MHz), 
           .D(n29477));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i165 (.Q(\data_in_frame[20] [4]), .C(clk16MHz), 
           .D(n29481));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i166 (.Q(\data_in_frame[20] [5]), .C(clk16MHz), 
           .D(n29484));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i167 (.Q(\data_in_frame[20] [6]), .C(clk16MHz), 
           .D(n29487));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i168 (.Q(\data_in_frame[20] [7]), .C(clk16MHz), 
           .D(n29490));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i169 (.Q(\data_in_frame[21][0] ), .C(clk16MHz), 
           .D(n29493));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i170 (.Q(\data_in_frame[21][1] ), .C(clk16MHz), 
           .D(n29496));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i171 (.Q(\data_in_frame[21][2] ), .C(clk16MHz), 
           .D(n29499));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i172 (.Q(\data_in_frame[21][3] ), .C(clk16MHz), 
           .D(n29506));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i173 (.Q(\data_in_frame[21][4] ), .C(clk16MHz), 
           .D(n29509));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i174 (.Q(\data_in_frame[21][5] ), .C(clk16MHz), 
           .D(n29512));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i175 (.Q(\data_in_frame[21]_c [6]), .C(clk16MHz), 
           .D(n54683));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i176 (.Q(\data_in_frame[21] [7]), .C(clk16MHz), 
           .D(n54583));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i177 (.Q(\data_in_frame[22] [0]), .C(clk16MHz), 
           .D(n54577));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i24 (.Q(\data_in_frame[2]_c [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29893));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i23 (.Q(\data_in_frame[2]_c [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29890));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i22 (.Q(\data_in_frame[2]_c [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29887));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i21 (.Q(\data_in_frame[2]_c [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29884));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i20 (.Q(\data_in_frame[2]_c [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29881));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i19 (.Q(\data_in_frame[2]_c [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29878));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i18 (.Q(\data_in_frame[2]_c [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29875));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i17 (.Q(\data_in_frame[2] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29872));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i16 (.Q(\data_in_frame[1] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29869));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i15 (.Q(\data_in_frame[1] [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29866));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1245 (.I0(n51189), .I1(n56112), .I2(n59476), 
            .I3(Kp_23__N_1067), .O(n59482));
    defparam i1_4_lut_adj_1245.LUT_INIT = 16'h9669;
    SB_DFFE data_in_frame_0___i14 (.Q(\data_in_frame[1] [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29863));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i13 (.Q(\data_in_frame[1] [4]), .C(clk16MHz), 
            .E(VCC_net), .D(n29860));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i12 (.Q(\data_in_frame[1]_c [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29857));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i11 (.Q(\data_in_frame[1]_c [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29854));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i10 (.Q(\data_in_frame[1]_c [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29851));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i9 (.Q(\data_in_frame[1] [0]), .C(clk16MHz), 
            .E(VCC_net), .D(n29848));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i8 (.Q(\data_in_frame[0] [7]), .C(clk16MHz), 
            .E(VCC_net), .D(n29845));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i7 (.Q(\data_in_frame[0]_c [6]), .C(clk16MHz), 
            .E(VCC_net), .D(n29842));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1246 (.I0(n51250), .I1(n56153), .I2(n55923), 
            .I3(n59482), .O(n24683));
    defparam i1_4_lut_adj_1246.LUT_INIT = 16'h6996;
    SB_DFFE data_in_frame_0___i6 (.Q(\data_in_frame[0]_c [5]), .C(clk16MHz), 
            .E(VCC_net), .D(n29839));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i5 (.Q(\data_in_frame[0][4] ), .C(clk16MHz), 
            .E(VCC_net), .D(n29836));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i4 (.Q(\data_in_frame[0]_c [3]), .C(clk16MHz), 
            .E(VCC_net), .D(n29833));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i3 (.Q(\data_in_frame[0]_c [2]), .C(clk16MHz), 
            .E(VCC_net), .D(n29830));   // verilog/coms.v(130[12] 305[6])
    SB_DFFE data_in_frame_0___i2 (.Q(\data_in_frame[0]_c [1]), .C(clk16MHz), 
            .E(VCC_net), .D(n29827));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i178 (.Q(\data_in_frame[22] [1]), .C(clk16MHz), 
           .D(n29524));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i179 (.Q(\data_in_frame[22] [2]), .C(clk16MHz), 
           .D(n54663));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i180 (.Q(\data_in_frame[22] [3]), .C(clk16MHz), 
           .D(n29530));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i181 (.Q(\data_in_frame[22] [4]), .C(clk16MHz), 
           .D(n29533));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i182 (.Q(\data_in_frame[22] [5]), .C(clk16MHz), 
           .D(n29537));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i183 (.Q(\data_in_frame[22] [6]), .C(clk16MHz), 
           .D(n29540));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i184 (.Q(\data_in_frame[22] [7]), .C(clk16MHz), 
           .D(n29543));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i185 (.Q(\data_in_frame[23] [0]), .C(clk16MHz), 
           .D(n29546));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i186 (.Q(\data_in_frame[23] [1]), .C(clk16MHz), 
           .D(n29549));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i187 (.Q(\data_in_frame[23] [2]), .C(clk16MHz), 
           .D(n29552));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i27 (.Q(\data_in_frame[3] [2]), .C(clk16MHz), 
           .D(n54803));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i188 (.Q(\data_in_frame[23] [3]), .C(clk16MHz), 
           .D(n29555));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i189 (.Q(\data_in_frame[23] [4]), .C(clk16MHz), 
           .D(n29558));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i190 (.Q(\data_in_frame[23] [5]), .C(clk16MHz), 
           .D(n54697));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i191 (.Q(\data_in_frame[23] [6]), .C(clk16MHz), 
           .D(n54695));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i192 (.Q(\data_in_frame[23]_c [7]), .C(clk16MHz), 
           .D(n54687));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i1 (.Q(\data_in_frame[0]_c [0]), .C(clk16MHz), 
           .D(n29597));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i28 (.Q(\data_in_frame[3][3] ), .C(clk16MHz), 
           .D(n28940));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i29 (.Q(\data_in_frame[3] [4]), .C(clk16MHz), 
           .D(n54743));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i30 (.Q(\data_in_frame[3][5] ), .C(clk16MHz), 
           .D(n28946));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i31 (.Q(\data_in_frame[3][6] ), .C(clk16MHz), 
           .D(n28949));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i32 (.Q(\data_in_frame[3][7] ), .C(clk16MHz), 
           .D(n28952));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i33 (.Q(\data_in_frame[4] [0]), .C(clk16MHz), 
           .D(n54733));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i34 (.Q(\data_in_frame[4] [1]), .C(clk16MHz), 
           .D(n28958));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i1 (.Q(deadband[1]), .C(clk16MHz), .D(n29753), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i2 (.Q(deadband[2]), .C(clk16MHz), .D(n29752), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i3 (.Q(deadband[3]), .C(clk16MHz), .D(n29751), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i4 (.Q(deadband[4]), .C(clk16MHz), .D(n29750), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i5 (.Q(deadband[5]), .C(clk16MHz), .D(n29749), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i6 (.Q(deadband[6]), .C(clk16MHz), .D(n29748), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i7 (.Q(deadband[7]), .C(clk16MHz), .D(n29747), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i8 (.Q(deadband[8]), .C(clk16MHz), .D(n29746), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i9 (.Q(deadband[9]), .C(clk16MHz), .D(n29745), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i10 (.Q(deadband[10]), .C(clk16MHz), .D(n29744), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i11 (.Q(deadband[11]), .C(clk16MHz), .D(n29743), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i12 (.Q(deadband[12]), .C(clk16MHz), .D(n29742), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i13 (.Q(deadband[13]), .C(clk16MHz), .D(n29741), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i14 (.Q(deadband[14]), .C(clk16MHz), .D(n29740), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i15 (.Q(deadband[15]), .C(clk16MHz), .D(n29739), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i16 (.Q(deadband[16]), .C(clk16MHz), .D(n29738), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i17 (.Q(deadband[17]), .C(clk16MHz), .D(n29737), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i18 (.Q(deadband[18]), .C(clk16MHz), .D(n29736), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i19 (.Q(deadband[19]), .C(clk16MHz), .D(n29735), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i20 (.Q(deadband[20]), .C(clk16MHz), .D(n29734), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i21 (.Q(deadband[21]), .C(clk16MHz), .D(n29733), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i22 (.Q(deadband[22]), .C(clk16MHz), .D(n29732), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i23 (.Q(deadband[23]), .C(clk16MHz), .D(n29731), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk16MHz), .D(n29730), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk16MHz), .D(n29729), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk16MHz), .D(n29728), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk16MHz), .D(n29727), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk16MHz), .D(n29726), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk16MHz), .D(n29725), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk16MHz), .D(n29724), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk16MHz), .D(n29723), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk16MHz), .D(n29722), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk16MHz), .D(n29721), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk16MHz), .D(n29720), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk16MHz), .D(n29719), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk16MHz), .D(n29718), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk16MHz), .D(n29717), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk16MHz), .D(n29716), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk16MHz), .D(n29715), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk16MHz), .D(n29714), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk16MHz), .D(n29713), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk16MHz), .D(n29712), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk16MHz), .D(n29711), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk16MHz), .D(n29710), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk16MHz), .D(n29709), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk16MHz), .D(n29708), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i1 (.Q(\Kp[1] ), .C(clk16MHz), .D(n29707), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i2 (.Q(\Kp[2] ), .C(clk16MHz), .D(n29706), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS Kp_i3 (.Q(\Kp[3] ), .C(clk16MHz), .D(n29705), .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i4 (.Q(\Kp[4] ), .C(clk16MHz), .D(n29704), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i5 (.Q(\Kp[5] ), .C(clk16MHz), .D(n29703), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i6 (.Q(\Kp[6] ), .C(clk16MHz), .D(n29702), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i7 (.Q(\Kp[7] ), .C(clk16MHz), .D(n29701), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i8 (.Q(\Kp[8] ), .C(clk16MHz), .D(n29700), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i9 (.Q(\Kp[9] ), .C(clk16MHz), .D(n29699), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i10 (.Q(\Kp[10] ), .C(clk16MHz), .D(n29698), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i11 (.Q(\Kp[11] ), .C(clk16MHz), .D(n29697), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i12 (.Q(\Kp[12] ), .C(clk16MHz), .D(n29696), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i13 (.Q(\Kp[13] ), .C(clk16MHz), .D(n29695), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i14 (.Q(\Kp[14] ), .C(clk16MHz), .D(n29694), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i15 (.Q(\Kp[15] ), .C(clk16MHz), .D(n29693), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i1 (.Q(\Ki[1] ), .C(clk16MHz), .D(n29692), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i2 (.Q(\Ki[2] ), .C(clk16MHz), .D(n29691), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i3 (.Q(\Ki[3] ), .C(clk16MHz), .D(n29690), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i4 (.Q(\Ki[4] ), .C(clk16MHz), .D(n29689), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i5 (.Q(\Ki[5] ), .C(clk16MHz), .D(n29688), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i6 (.Q(\Ki[6] ), .C(clk16MHz), .D(n29687), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i7 (.Q(\Ki[7] ), .C(clk16MHz), .D(n29686), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i8 (.Q(\Ki[8] ), .C(clk16MHz), .D(n29685), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i9 (.Q(\Ki[9] ), .C(clk16MHz), .D(n29684), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i10 (.Q(\Ki[10] ), .C(clk16MHz), .D(n29683), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i11 (.Q(\Ki[11] ), .C(clk16MHz), .D(n29682), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i12 (.Q(\Ki[12] ), .C(clk16MHz), .D(n29681), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i13 (.Q(\Ki[13] ), .C(clk16MHz), .D(n29680), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i14 (.Q(\Ki[14] ), .C(clk16MHz), .D(n29679), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i15 (.Q(\Ki[15] ), .C(clk16MHz), .D(n29678), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk16MHz), .D(n29677));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1247 (.I0(\data_in_frame[10] [7]), .I1(n24683), 
            .I2(\data_in_frame[11] [1]), .I3(n50498), .O(n55652));
    defparam i1_4_lut_adj_1247.LUT_INIT = 16'h9669;
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk16MHz), .D(n29676));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 n66873_bdd_4_lut (.I0(n66873), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(byte_transmit_counter[1]), 
            .O(n66876));
    defparam n66873_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_49616 (.I0(byte_transmit_counter[1]), 
            .I1(n59988), .I2(n59989), .I3(byte_transmit_counter[2]), .O(n66675));
    defparam byte_transmit_counter_1__bdd_4_lut_49616.LUT_INIT = 16'he4aa;
    SB_LUT4 n66675_bdd_4_lut (.I0(n66675), .I1(n60148), .I2(n60147), .I3(byte_transmit_counter[2]), 
            .O(n66678));
    defparam n66675_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0___i35 (.Q(\data_in_frame[4] [2]), .C(clk16MHz), 
           .D(n28961));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk16MHz), .D(n29674));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk16MHz), .D(n29673));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk16MHz), .D(n29672));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk16MHz), .D(n29671));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk16MHz), .D(n29670));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk16MHz), .D(n29669));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk16MHz), .D(n29668));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk16MHz), .D(n29667));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk16MHz), .D(n29666));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk16MHz), .D(n29665));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk16MHz), .D(n29664));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk16MHz), .D(n29663));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk16MHz), .D(n29662));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk16MHz), .D(n29661));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk16MHz), .D(n29660));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk16MHz), .D(n29659));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk16MHz), .D(n29658));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk16MHz), .D(n29657));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk16MHz), .D(n29656));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk16MHz), .D(n29655));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk16MHz), .D(n29654));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk16MHz), .D(n29653));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk16MHz), .D(n29652));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk16MHz), .D(n29651));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk16MHz), .D(n29650));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk16MHz), .D(n29649));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk16MHz), .D(n29648));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk16MHz), .D(n29647));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i1 (.Q(current_limit[1]), .C(clk16MHz), .D(n29646));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i2 (.Q(current_limit[2]), .C(clk16MHz), .D(n29645));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i3 (.Q(current_limit[3]), .C(clk16MHz), .D(n29644));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i4 (.Q(current_limit[4]), .C(clk16MHz), .D(n29643));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i5 (.Q(current_limit[5]), .C(clk16MHz), .D(n29642));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i6 (.Q(current_limit[6]), .C(clk16MHz), .D(n29641));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i7 (.Q(current_limit[7]), .C(clk16MHz), .D(n29640));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i8 (.Q(current_limit[8]), .C(clk16MHz), .D(n29639));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i9 (.Q(current_limit[9]), .C(clk16MHz), .D(n29638));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i10 (.Q(current_limit[10]), .C(clk16MHz), .D(n29637));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i11 (.Q(current_limit[11]), .C(clk16MHz), .D(n29636));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i12 (.Q(current_limit[12]), .C(clk16MHz), .D(n29635));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i13 (.Q(current_limit[13]), .C(clk16MHz), .D(n29634));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i14 (.Q(current_limit[14]), .C(clk16MHz), .D(n29633));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1248 (.I0(Kp_23__N_1085), .I1(n25839), .I2(n25282), 
            .I3(\data_in_frame[9] [3]), .O(Kp_23__N_1080));   // verilog/coms.v(88[17:63])
    defparam i3_4_lut_adj_1248.LUT_INIT = 16'h6996;
    SB_DFF current_limit_i0_i15 (.Q(current_limit[15]), .C(clk16MHz), .D(n29632));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk16MHz), .D(n29631), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk16MHz), .D(n29630), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk16MHz), .D(n29629), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk16MHz), .D(n29628), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk16MHz), .D(n29627), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk16MHz), .D(n29626), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk16MHz), .D(n29625), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFS PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk16MHz), .D(n29624), 
            .S(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk16MHz), .D(n29623), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk16MHz), .D(n29622), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk16MHz), .D(n29621), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk16MHz), .D(n29620), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk16MHz), .D(n29619), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk16MHz), .D(n29618), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk16MHz), .D(n29617), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk16MHz), .D(n29616), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk16MHz), .D(n29615), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk16MHz), .D(n29614), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk16MHz), .D(n29613), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk16MHz), .D(n29612), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk16MHz), .D(n29611), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk16MHz), .D(n29610), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk16MHz), .D(n29609), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i36 (.Q(\data_in_frame[4] [3]), .C(clk16MHz), 
           .D(n28964));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i37 (.Q(\data_in_frame[4] [4]), .C(clk16MHz), 
           .D(n28967));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i38 (.Q(\data_in_frame[4] [5]), .C(clk16MHz), 
           .D(n54819));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i39 (.Q(\data_in_frame[4] [6]), .C(clk16MHz), 
           .D(n54747));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1249 (.I0(\data_in_frame[16] [0]), .I1(n50907), 
            .I2(n55745), .I3(n26028), .O(n56174));
    defparam i3_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1250 (.I0(n51256), .I1(n55757), .I2(GND_net), 
            .I3(GND_net), .O(n26028));
    defparam i1_2_lut_adj_1250.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0___i40 (.Q(\data_in_frame[4] [7]), .C(clk16MHz), 
           .D(n28976));   // verilog/coms.v(130[12] 305[6])
    SB_DFFESS data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk16MHz), 
            .E(n2882), .D(n2_adj_5532), .S(n55293));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1251 (.I0(n50907), .I1(n55829), .I2(n50272), 
            .I3(n51247), .O(n24707));
    defparam i3_4_lut_adj_1251.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0___i41 (.Q(\data_in_frame[5] [0]), .C(clk16MHz), 
           .D(n28979));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_2_lut_adj_1252 (.I0(\data_in_frame[18] [3]), .I1(n24707), 
            .I2(GND_net), .I3(GND_net), .O(n50169));
    defparam i1_2_lut_adj_1252.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1253 (.I0(\data_in_frame[15] [5]), .I1(n55975), 
            .I2(\data_in_frame[17] [7]), .I3(GND_net), .O(n24695));
    defparam i2_3_lut_adj_1253.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1254 (.I0(\data_in_frame[7] [0]), .I1(\data_in_frame[4] [6]), 
            .I2(n25908), .I3(GND_net), .O(n55787));
    defparam i2_3_lut_adj_1254.LUT_INIT = 16'h9696;
    SB_LUT4 i49217_3_lut (.I0(\data_in_frame[0][4] ), .I1(\data_in_frame[2]_c [5]), 
            .I2(\data_in_frame[0]_c [3]), .I3(GND_net), .O(n66279));   // verilog/coms.v(99[12:25])
    defparam i49217_3_lut.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0___i42 (.Q(\data_in_frame[5] [1]), .C(clk16MHz), 
           .D(n28982));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i4_4_lut_adj_1255 (.I0(\data_in_frame[0][4] ), .I1(\data_in_frame[0]_c [6]), 
            .I2(ID[4]), .I3(ID[6]), .O(n12_adj_5533));   // verilog/coms.v(241[12:32])
    defparam i4_4_lut_adj_1255.LUT_INIT = 16'h7bde;
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk16MHz), .D(n28934));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i2_4_lut_adj_1256 (.I0(\data_in_frame[0]_c [1]), .I1(\data_in_frame[0]_c [2]), 
            .I2(ID[1]), .I3(ID[2]), .O(n10_adj_5534));   // verilog/coms.v(241[12:32])
    defparam i2_4_lut_adj_1256.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_1257 (.I0(ID[7]), .I1(\data_in_frame[0]_c [5]), 
            .I2(\data_in_frame[0] [7]), .I3(ID[5]), .O(n11_adj_5535));   // verilog/coms.v(241[12:32])
    defparam i3_4_lut_adj_1257.LUT_INIT = 16'h7bde;
    SB_DFF data_in_frame_0___i43 (.Q(\data_in_frame[5] [2]), .C(clk16MHz), 
           .D(n28985));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i49201_3_lut (.I0(rx_data[0]), .I1(\data_in_frame[7] [0]), .I2(n27906), 
            .I3(GND_net), .O(n54823));   // verilog/coms.v(94[13:20])
    defparam i49201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1258 (.I0(\data_in_frame[0]_c [0]), .I1(\data_in_frame[0]_c [3]), 
            .I2(ID[0]), .I3(ID[3]), .O(n9_adj_5536));   // verilog/coms.v(241[12:32])
    defparam i1_4_lut_adj_1258.LUT_INIT = 16'h7bde;
    SB_DFFR \FRAME_MATCHER.i_2043__i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk16MHz), 
            .D(n27570), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk16MHz), 
            .D(n27572), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i3  (.Q(\FRAME_MATCHER.i[3] ), .C(clk16MHz), 
            .D(n27574), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i4  (.Q(\FRAME_MATCHER.i[4] ), .C(clk16MHz), 
            .D(n27576), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i5  (.Q(\FRAME_MATCHER.i[5] ), .C(clk16MHz), 
            .D(n27578), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk16MHz), 
            .D(n27580), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk16MHz), 
            .D(n27582), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk16MHz), 
            .D(n27584), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk16MHz), 
            .D(n27586), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk16MHz), 
            .D(n27588), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk16MHz), 
            .D(n27590), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk16MHz), 
            .D(n27592), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk16MHz), 
            .D(n27594), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk16MHz), 
            .D(n27596), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk16MHz), 
            .D(n27598), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk16MHz), 
            .D(n27600), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk16MHz), 
            .D(n27602), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk16MHz), 
            .D(n27604), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk16MHz), 
            .D(n27606), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk16MHz), 
            .D(n27608), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk16MHz), 
            .D(n27610), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk16MHz), 
            .D(n27612), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk16MHz), 
            .D(n27614), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk16MHz), 
            .D(n27616), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk16MHz), 
            .D(n27618), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk16MHz), 
            .D(n27620), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk16MHz), 
            .D(n27622), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk16MHz), 
            .D(n27624), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk16MHz), 
            .D(n27626), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk16MHz), 
            .D(n27628), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFFR \FRAME_MATCHER.i_2043__i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk16MHz), 
            .D(n27630), .R(reset));   // verilog/coms.v(158[12:15])
    SB_DFF data_in_frame_0___i44 (.Q(\data_in_frame[5] [3]), .C(clk16MHz), 
           .D(n28988));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i7_4_lut_adj_1259 (.I0(n9_adj_5536), .I1(n11_adj_5535), .I2(n10_adj_5534), 
            .I3(n12_adj_5533), .O(n57981));   // verilog/coms.v(241[12:32])
    defparam i7_4_lut_adj_1259.LUT_INIT = 16'hfffe;
    SB_DFF data_in_frame_0___i45 (.Q(\data_in_frame[5] [4]), .C(clk16MHz), 
           .D(n28991));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i46 (.Q(\data_in_frame[5] [5]), .C(clk16MHz), 
           .D(n28994));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i47 (.Q(\data_in_frame[5] [6]), .C(clk16MHz), 
           .D(n28997));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i3_4_lut_adj_1260 (.I0(n66279), .I1(n56072), .I2(n55787), 
            .I3(\data_in_frame[6][7] ), .O(n57296));
    defparam i3_4_lut_adj_1260.LUT_INIT = 16'h9669;
    SB_DFFR PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk16MHz), .D(n28924), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF current_limit_i0_i0 (.Q(current_limit[0]), .C(clk16MHz), .D(n28923));   // verilog/coms.v(130[12] 305[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk16MHz), .D(n28922));   // verilog/coms.v(130[12] 305[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk16MHz), .D(n28921));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Ki_i0 (.Q(\Ki[0] ), .C(clk16MHz), .D(n28920), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR Kp_i0 (.Q(\Kp[0] ), .C(clk16MHz), .D(n28919), .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk16MHz), .D(n28918), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i48 (.Q(\data_in_frame[5] [7]), .C(clk16MHz), 
           .D(n29000));   // verilog/coms.v(130[12] 305[6])
    SB_DFF data_in_frame_0___i49 (.Q(\data_in_frame[6][0] ), .C(clk16MHz), 
           .D(n29003));   // verilog/coms.v(130[12] 305[6])
    SB_DFFR deadband_i0_i0 (.Q(deadband[0]), .C(clk16MHz), .D(n28911), 
            .R(reset));   // verilog/coms.v(130[12] 305[6])
    SB_LUT4 i1_4_lut_adj_1261 (.I0(n30), .I1(\data_in_frame[5] [1]), .I2(\data_in_frame[3] [1]), 
            .I3(\data_in_frame[7] [3]), .O(n59532));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1262 (.I0(n59532), .I1(n25770), .I2(\data_in_frame[4] [7]), 
            .I3(\data_in_frame[2]_c [6]), .O(n55665));   // verilog/coms.v(99[12:25])
    defparam i1_4_lut_adj_1262.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1263 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[7][1] ), 
            .I2(\data_in_frame[6][7] ), .I3(GND_net), .O(n56261));   // verilog/coms.v(73[16:27])
    defparam i2_3_lut_adj_1263.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1264 (.I0(\data_in_frame[5] [2]), .I1(n55665), 
            .I2(GND_net), .I3(GND_net), .O(n26413));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1264.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1265 (.I0(n55847), .I1(n56261), .I2(n50417), 
            .I3(GND_net), .O(n56112));
    defparam i2_3_lut_adj_1265.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1266 (.I0(n55689), .I1(n56072), .I2(\data_in_frame[4] [5]), 
            .I3(GND_net), .O(n51230));
    defparam i2_3_lut_adj_1266.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1267 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[4] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n59640));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_adj_1267.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_4_lut (.I0(n26406), .I1(\data_in_frame[8] [2]), .I2(n25500), 
            .I3(n25572), .O(n20_adj_5537));   // verilog/coms.v(79[16:43])
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6900;
    SB_LUT4 i1_3_lut_adj_1268 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[2]_c [6]), 
            .I2(\data_in_frame[3][0] ), .I3(GND_net), .O(n59646));   // verilog/coms.v(81[16:27])
    defparam i1_3_lut_adj_1268.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1269 (.I0(n56059), .I1(\data_in_frame[4] [4]), 
            .I2(n59640), .I3(\data_in_frame[3][7] ), .O(n59652));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1269.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1270 (.I0(n25321), .I1(\data_in_frame[7][6] ), 
            .I2(n25481), .I3(GND_net), .O(n25572));
    defparam i1_2_lut_3_lut_adj_1270.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1271 (.I0(n55867), .I1(n59646), .I2(\data_in_frame[5] [0]), 
            .I3(\data_in_frame[3][5] ), .O(n59656));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1272 (.I0(n25321), .I1(\data_in_frame[7][6] ), 
            .I2(\data_in_frame[7][7] ), .I3(n10_adj_5527), .O(n58201));
    defparam i5_3_lut_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1273 (.I0(n56065), .I1(n59656), .I2(n59652), 
            .I3(n55769), .O(n59660));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1273.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1274 (.I0(n56062), .I1(n59660), .I2(n30), .I3(n23332), 
            .O(n59666));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1274.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1275 (.I0(n55748), .I1(n50165), .I2(n56007), 
            .I3(n59666), .O(n59672));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1276 (.I0(n59672), .I1(n25769), .I2(n25321), 
            .I3(n56078), .O(n51223));   // verilog/coms.v(81[16:27])
    defparam i1_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter_c[3]), 
            .I1(n64943), .I2(n63134), .I3(byte_transmit_counter_c[4]), 
            .O(n66867));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i13176_3_lut (.I0(\data_in_frame[6][6] ), .I1(rx_data[6]), .I2(n27904), 
            .I3(GND_net), .O(n29021));   // verilog/coms.v(130[12] 305[6])
    defparam i13176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 n66867_bdd_4_lut (.I0(n66867), .I1(n66636), .I2(n7_adj_5538), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[6]));
    defparam n66867_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1277 (.I0(n50417), .I1(n51223), .I2(Kp_23__N_709), 
            .I3(\data_in_frame[6][0] ), .O(n50366));   // verilog/coms.v(88[17:70])
    defparam i1_4_lut_adj_1277.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1278 (.I0(\data_in_frame[8] [7]), .I1(n51230), 
            .I2(GND_net), .I3(GND_net), .O(n51294));
    defparam i1_2_lut_adj_1278.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1279 (.I0(n23345), .I1(n50366), .I2(\data_in_frame[5] [5]), 
            .I3(GND_net), .O(n24777));
    defparam i2_3_lut_adj_1279.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1280 (.I0(\data_in_frame[6]_c [5]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5539));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1280.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1281 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [1]), 
            .I2(\data_in_frame[6][6] ), .I3(n6_adj_5539), .O(n55596));   // verilog/coms.v(88[17:28])
    defparam i4_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1282 (.I0(\data_in_frame[6][7] ), .I1(n55596), 
            .I2(\data_in_frame[6] [4]), .I3(GND_net), .O(Kp_23__N_709));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_adj_1282.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1283 (.I0(\data_in_frame[3][6] ), .I1(\data_in_frame[6][0] ), 
            .I2(GND_net), .I3(GND_net), .O(n25960));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1283.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1284 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n56065));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1284.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1285 (.I0(\data_in_frame[1]_c [3]), .I1(\data_in_frame[3] [4]), 
            .I2(n56041), .I3(GND_net), .O(n23345));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1285.LUT_INIT = 16'h9696;
    SB_LUT4 i14003_3_lut_4_lut (.I0(n8_adj_5430), .I1(n55507), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n29848));
    defparam i14003_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1286 (.I0(\data_in_frame[1]_c [3]), .I1(\data_in_frame[3] [4]), 
            .I2(\data_in_frame[1]_c [2]), .I3(GND_net), .O(n25481));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1286.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1287 (.I0(n66267), .I1(n25933), .I2(\data_in_frame[1] [5]), 
            .I3(GND_net), .O(n56078));
    defparam i1_2_lut_3_lut_adj_1287.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1288 (.I0(n25481), .I1(n56065), .I2(n55675), 
            .I3(n25960), .O(n26406));   // verilog/coms.v(79[16:43])
    defparam i3_4_lut_adj_1288.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1289 (.I0(\data_in_frame[4] [1]), .I1(n55560), 
            .I2(\data_in_frame[2]_c [1]), .I3(\data_in_frame[4] [2]), .O(n56004));   // verilog/coms.v(99[12:25])
    defparam i3_4_lut_adj_1289.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1290 (.I0(n66267), .I1(n25933), .I2(\data_in_frame[4] [4]), 
            .I3(\data_in_frame[6][6] ), .O(n56072));
    defparam i2_3_lut_4_lut_adj_1290.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1291 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[3][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5540));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1291.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1292 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [5]), 
            .I2(n56004), .I3(n6_adj_5540), .O(n55808));   // verilog/coms.v(73[16:69])
    defparam i4_4_lut_adj_1292.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1293 (.I0(n25908), .I1(\data_in_frame[2]_c [1]), 
            .I2(GND_net), .I3(GND_net), .O(n56007));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1293.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1294 (.I0(\data_in_frame[6]_c [5]), .I1(\data_in_frame[4] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5541));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1294.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1295 (.I0(n55560), .I1(\data_in_frame[4] [4]), 
            .I2(n56007), .I3(n6_adj_5541), .O(n55689));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1295.LUT_INIT = 16'h6996;
    SB_LUT4 i49215_3_lut (.I0(\data_in_frame[0]_c [5]), .I1(\data_in_frame[2]_c [6]), 
            .I2(\data_in_frame[0][4] ), .I3(GND_net), .O(n66277));   // verilog/coms.v(99[12:25])
    defparam i49215_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1296 (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[7][4] ), 
            .I2(n26166), .I3(n6_adj_5531), .O(n55698));
    defparam i4_4_lut_adj_1296.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1297 (.I0(\data_in_frame[5] [2]), .I1(n55698), 
            .I2(n66277), .I3(GND_net), .O(n50744));
    defparam i2_3_lut_adj_1297.LUT_INIT = 16'h6969;
    SB_LUT4 equal_2036_i7_2_lut (.I0(Kp_23__N_974), .I1(\data_in_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5542));   // verilog/coms.v(239[9:81])
    defparam equal_2036_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1298 (.I0(n55681), .I1(n55808), .I2(\data_in_frame[8] [4]), 
            .I3(GND_net), .O(n25514));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_adj_1298.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_0__3__I_0_2_lut (.I0(\data_in_frame[0]_c [3]), .I1(\data_in_frame[0]_c [2]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_758));   // verilog/coms.v(77[16:27])
    defparam data_in_frame_0__3__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1299 (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[2]_c [7]), 
            .I2(Kp_23__N_767), .I3(\data_in_frame[0]_c [5]), .O(n25769));
    defparam i1_4_lut_adj_1299.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1300 (.I0(Kp_23__N_767), .I1(n25769), .I2(\data_in_frame[0] [7]), 
            .I3(GND_net), .O(n25770));   // verilog/coms.v(74[16:69])
    defparam i1_3_lut_adj_1300.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1301 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n55675));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1301.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1302 (.I0(\data_in_frame[1]_c [3]), .I1(\data_in_frame[1]_c [1]), 
            .I2(GND_net), .I3(GND_net), .O(n59488));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1302.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1303 (.I0(n55668), .I1(n55675), .I2(n59488), 
            .I3(\data_in_frame[1]_c [2]), .O(Kp_23__N_767));   // verilog/coms.v(73[16:69])
    defparam i1_4_lut_adj_1303.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1304 (.I0(\data_in_frame[2]_c [5]), .I1(\data_in_frame[0]_c [3]), 
            .I2(\data_in_frame[0]_c [5]), .I3(GND_net), .O(n30));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1304.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1305 (.I0(\data_in_frame[5] [0]), .I1(\data_in_frame[2]_c [6]), 
            .I2(n30), .I3(GND_net), .O(n55847));   // verilog/coms.v(99[12:25])
    defparam i2_3_lut_adj_1305.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1306 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n55769));
    defparam i1_2_lut_adj_1306.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_1__4__I_0_2_lut (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1]_c [3]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_843));   // verilog/coms.v(78[16:27])
    defparam data_in_frame_1__4__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_143_i2_4_lut (.I0(\data_out_frame[17] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5513));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_143_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1307 (.I0(\data_in_frame[3][3] ), .I1(\data_in_frame[3] [1]), 
            .I2(\data_in_frame[5] [3]), .I3(GND_net), .O(n55867));
    defparam i2_3_lut_adj_1307.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_60_i2_4_lut (.I0(\data_out_frame[7] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[12] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5431));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_60_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_4_lut_adj_1308 (.I0(n25770), .I1(\data_in_frame[5] [4]), 
            .I2(n57764), .I3(\data_in_frame[7][5] ), .O(n25557));
    defparam i2_4_lut_adj_1308.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1309 (.I0(n55769), .I1(n55847), .I2(\data_in_frame[7][2] ), 
            .I3(n26166), .O(n12_adj_5543));
    defparam i5_4_lut_adj_1309.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1310 (.I0(Kp_23__N_758), .I1(n12_adj_5543), .I2(n25769), 
            .I3(\data_in_frame[2]_c [4]), .O(n26031));
    defparam i6_4_lut_adj_1310.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1311 (.I0(\data_in_frame[4] [5]), .I1(n51223), 
            .I2(GND_net), .I3(GND_net), .O(n56222));
    defparam i1_2_lut_adj_1311.LUT_INIT = 16'h9999;
    SB_LUT4 i6_4_lut_adj_1312 (.I0(n56222), .I1(n25908), .I2(n55695), 
            .I3(\data_in_frame[8] [1]), .O(n14_adj_5544));
    defparam i6_4_lut_adj_1312.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1313 (.I0(Kp_23__N_709), .I1(n56078), .I2(n25933), 
            .I3(\data_in_frame[3][6] ), .O(n13_adj_5545));
    defparam i5_4_lut_adj_1313.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1314 (.I0(n13_adj_5545), .I1(n51250), .I2(n14_adj_5544), 
            .I3(\data_in_frame[8] [0]), .O(n21));
    defparam i4_4_lut_adj_1314.LUT_INIT = 16'h2184;
    SB_LUT4 i9_3_lut (.I0(n26031), .I1(n25557), .I2(n26001), .I3(GND_net), 
            .O(n26_adj_5546));
    defparam i9_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i42815_4_lut (.I0(n25514), .I1(n7_adj_5542), .I2(n25428), 
            .I3(n50744), .O(n59868));
    defparam i42815_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n21), .I1(n24777), .I2(n51294), .I3(\data_in_frame[7][7] ), 
            .O(n28));
    defparam i11_4_lut.LUT_INIT = 16'h8020;
    SB_LUT4 i15_4_lut (.I0(n59868), .I1(n56112), .I2(n26_adj_5546), .I3(n26413), 
            .O(n32));
    defparam i15_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i42683_2_lut (.I0(n57296), .I1(n57981), .I2(GND_net), .I3(GND_net), 
            .O(n59732));
    defparam i42683_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut (.I0(n55695), .I1(n56075), .I2(n25960), .I3(n26406), 
            .O(n56027));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut (.I0(n59732), .I1(n32), .I2(n28), .I3(n20_adj_5537), 
            .O(LED_N_3408));
    defparam i16_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i4_4_lut_adj_1315 (.I0(\data_in_frame[18] [1]), .I1(n24695), 
            .I2(n50169), .I3(\data_in_frame[20] [4]), .O(n10_adj_5547));
    defparam i4_4_lut_adj_1315.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1316 (.I0(\data_in_frame[22] [1]), .I1(n56132), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5548));
    defparam i2_2_lut_adj_1316.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1317 (.I0(\data_in_frame[19]_c [7]), .I1(\data_in_frame[21] [7]), 
            .I2(\data_in_frame[20] [0]), .I3(GND_net), .O(n7_adj_5549));
    defparam i1_3_lut_adj_1317.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1318 (.I0(\data_in_frame[21][1] ), .I1(n57981), 
            .I2(\data_in_frame[23] [2]), .I3(n57376), .O(n59494));
    defparam i1_4_lut_adj_1318.LUT_INIT = 16'h1221;
    SB_LUT4 i1_4_lut_adj_1319 (.I0(n50370), .I1(n59494), .I2(n55815), 
            .I3(\data_in_frame[23] [4]), .O(n59496));
    defparam i1_4_lut_adj_1319.LUT_INIT = 16'h8448;
    SB_LUT4 i2_4_lut_adj_1320 (.I0(Kp_23__N_1607), .I1(\data_in_frame[21][1] ), 
            .I2(\data_in_frame[23] [3]), .I3(n55815), .O(n57334));
    defparam i2_4_lut_adj_1320.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1321 (.I0(n51173), .I1(n7_adj_5549), .I2(\data_in_frame[19]_c [5]), 
            .I3(n8_adj_5548), .O(n57397));
    defparam i5_4_lut_adj_1321.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1322 (.I0(\data_in_frame[20] [3]), .I1(n10_adj_5547), 
            .I2(\data_in_frame[22] [5]), .I3(GND_net), .O(n58102));
    defparam i5_3_lut_adj_1322.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_adj_1323 (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[22] [4]), 
            .I2(n56144), .I3(GND_net), .O(n8_adj_5550));
    defparam i3_3_lut_adj_1323.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1324 (.I0(n58102), .I1(n57397), .I2(n57334), 
            .I3(n59496), .O(n59502));
    defparam i1_4_lut_adj_1324.LUT_INIT = 16'h0400;
    SB_LUT4 i4_4_lut_adj_1325 (.I0(n57567), .I1(n8_adj_5550), .I2(\data_in_frame[20] [3]), 
            .I3(\data_in_frame[20] [2]), .O(n57426));
    defparam i4_4_lut_adj_1325.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1326 (.I0(\data_in_frame[22] [0]), .I1(n55932), 
            .I2(\data_in_frame[21] [7]), .I3(\data_in_frame[21]_c [6]), 
            .O(n57950));
    defparam i3_4_lut_adj_1326.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1327 (.I0(n55695), .I1(n56075), .I2(n25960), 
            .I3(\data_in_frame[8] [1]), .O(n55732));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_4_lut_adj_1327.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1328 (.I0(n57950), .I1(n57143), .I2(n57426), 
            .I3(n59502), .O(n59508));
    defparam i1_4_lut_adj_1328.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1329 (.I0(n50368), .I1(n59508), .I2(n55972), 
            .I3(\data_in_frame[23] [6]), .O(n59510));
    defparam i1_4_lut_adj_1329.LUT_INIT = 16'h8448;
    SB_LUT4 i4_4_lut_adj_1330 (.I0(n55929), .I1(\data_in_frame[19]_c [7]), 
            .I2(\data_in_frame[22] [3]), .I3(n56144), .O(n10_adj_5551));
    defparam i4_4_lut_adj_1330.LUT_INIT = 16'h6996;
    SB_LUT4 i43061_3_lut (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[17] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60123));
    defparam i43061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43062_3_lut (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[19] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60124));
    defparam i43062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43020_3_lut (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[23] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60082));
    defparam i43020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43019_3_lut (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[21] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60081));
    defparam i43019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47050_2_lut (.I0(n66786), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n63125));
    defparam i47050_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i42941_3_lut (.I0(\data_out_frame[8][7] ), .I1(\data_out_frame[9] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60003));
    defparam i42941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42942_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60004));
    defparam i42942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_adj_1331 (.I0(\data_in_frame[20] [2]), .I1(n10_adj_5551), 
            .I2(\data_in_frame[18] [1]), .I3(GND_net), .O(n57436));
    defparam i5_3_lut_adj_1331.LUT_INIT = 16'h9696;
    SB_LUT4 i43233_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60295));
    defparam i43233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43232_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60294));
    defparam i43232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1332 (.I0(\data_in_frame[23] [5]), .I1(n59510), 
            .I2(n50370), .I3(n50368), .O(n59512));
    defparam i1_4_lut_adj_1332.LUT_INIT = 16'h8448;
    SB_LUT4 i5_4_lut_adj_1333 (.I0(\data_in_frame[20] [0]), .I1(n55929), 
            .I2(\data_in_frame[19]_c [6]), .I3(\data_in_frame[22] [2]), 
            .O(n12_adj_5552));
    defparam i5_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 i46463_2_lut (.I0(\data_out_frame[9] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n62990));
    defparam i46463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i9_3_lut (.I0(\data_out_frame[10] [1]), 
            .I1(\data_out_frame[11] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n9_adj_5553));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i12_3_lut (.I0(\data_out_frame[14] [1]), 
            .I1(\data_out_frame[15] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n12_adj_5554));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i11_3_lut (.I0(\data_out_frame[12] [1]), 
            .I1(\data_out_frame[13] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n11_adj_5555));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46312_2_lut (.I0(\data_out_frame[9] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n62989));
    defparam i46312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1334 (.I0(n59512), .I1(n57436), .I2(\data_in_frame[23]_c [7]), 
            .I3(n55633), .O(n59516));
    defparam i1_4_lut_adj_1334.LUT_INIT = 16'h8008;
    SB_LUT4 i1_2_lut_adj_1335 (.I0(n55892), .I1(\data_in_frame[23] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5556));
    defparam i1_2_lut_adj_1335.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i9_3_lut (.I0(\data_out_frame[10] [0]), 
            .I1(\data_out_frame[11] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n9_adj_5557));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1336 (.I0(n24695), .I1(n12_adj_5552), .I2(n56132), 
            .I3(n51150), .O(n57404));
    defparam i6_4_lut_adj_1336.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1337 (.I0(n51243), .I1(\data_in_frame[20] [5]), 
            .I2(\data_in_frame[22] [7]), .I3(\data_in_frame[18] [5]), .O(n59632));
    defparam i1_4_lut_adj_1337.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i12_3_lut (.I0(\data_out_frame[14] [0]), 
            .I1(\data_out_frame[15] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n12_adj_5558));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i11_3_lut (.I0(\data_out_frame[12] [0]), 
            .I1(\data_out_frame[13] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n11_adj_5559));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i1_3_lut (.I0(\data_out_frame[0][3] ), 
            .I1(\data_out_frame[1][3] ), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n1_adj_5560));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42977_4_lut (.I0(n1_adj_5560), .I1(\data_out_frame[3][3] ), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n60039));
    defparam i42977_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i43004_3_lut (.I0(\data_out_frame[8][6] ), .I1(\data_out_frame[9] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60066));
    defparam i43004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43005_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60067));
    defparam i43005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43023_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60085));
    defparam i43023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43022_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60084));
    defparam i43022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46314_2_lut (.I0(\data_out_frame[0][4] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n62987));
    defparam i46314_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_rep_201_2_lut (.I0(n57376), .I1(n55892), .I2(GND_net), 
            .I3(GND_net), .O(n67347));
    defparam i1_rep_201_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i46276_2_lut (.I0(\data_out_frame[3][4] ), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n62988));
    defparam i46276_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_5561));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i4_3_lut (.I0(\data_out_frame[4] [4]), 
            .I1(\data_out_frame[5] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n4_adj_5562));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1338 (.I0(Kp_23__N_1607), .I1(n57404), .I2(n4_adj_5556), 
            .I3(n59516), .O(n59520));
    defparam i1_4_lut_adj_1338.LUT_INIT = 16'h1200;
    SB_LUT4 i1_4_lut_adj_1339 (.I0(n56246), .I1(n57376), .I2(n59632), 
            .I3(n55892), .O(n57780));
    defparam i1_4_lut_adj_1339.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1340 (.I0(\data_in_frame[23] [0]), .I1(n57780), 
            .I2(n59520), .I3(n67347), .O(n32097));
    defparam i1_4_lut_adj_1340.LUT_INIT = 16'h2010;
    SB_LUT4 i43028_3_lut (.I0(\data_out_frame[8][5] ), .I1(\data_out_frame[9] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60090));
    defparam i43028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43029_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60091));
    defparam i43029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43068_3_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[15] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60130));
    defparam i43068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43067_3_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[13] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60129));
    defparam i43067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43034_3_lut (.I0(\data_out_frame[8][4] ), .I1(\data_out_frame[9] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60096));
    defparam i43034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43035_3_lut (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[11] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60097));
    defparam i43035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43038_3_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[15] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60100));
    defparam i43038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43037_3_lut (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[13] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60099));
    defparam i43037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11709_3_lut (.I0(\data_out_frame[1][1] ), .I1(\data_out_frame[3][1] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n27553));   // verilog/coms.v(109[34:55])
    defparam i11709_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43047_3_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[7] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60109));
    defparam i43047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43048_4_lut (.I0(n60109), .I1(n27553), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n60110));
    defparam i43048_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i43046_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60108));
    defparam i43046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46471_2_lut (.I0(n66720), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n63136));
    defparam i46471_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48293_3_lut (.I0(n67038), .I1(n66594), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n65355));
    defparam i48293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47081_2_lut (.I0(byte_transmit_counter[0]), .I1(\data_out_frame[0][2] ), 
            .I2(GND_net), .I3(GND_net), .O(n63129));
    defparam i47081_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i18342_3_lut (.I0(n27904), .I1(rx_data[5]), .I2(\data_in_frame[6]_c [5]), 
            .I3(GND_net), .O(n29312));   // verilog/coms.v(94[13:20])
    defparam i18342_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i42999_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60061));
    defparam i42999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43000_4_lut (.I0(n60061), .I1(n63129), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n60062));
    defparam i43000_4_lut.LUT_INIT = 16'ha0ac;
    SB_LUT4 i42998_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60060));
    defparam i42998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46503_2_lut (.I0(n66756), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n63135));
    defparam i46503_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48295_3_lut (.I0(n66876), .I1(n66582), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n65357));
    defparam i48295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43083_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60145));
    defparam i43083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_301_i7_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/coms.v(157[7:23])
    defparam equal_301_i7_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i43084_4_lut (.I0(n60145), .I1(n27637), .I2(byte_transmit_counter[2]), 
            .I3(\data_out_frame[1][0] ), .O(n60146));
    defparam i43084_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i43082_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60144));
    defparam i43082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14006_3_lut_4_lut (.I0(n8_adj_5430), .I1(n55507), .I2(rx_data[1]), 
            .I3(\data_in_frame[1]_c [1]), .O(n29851));
    defparam i14006_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16264_4_lut (.I0(Kp_23__N_1748), .I1(\FRAME_MATCHER.i_31__N_2513 ), 
            .I2(n32097), .I3(LED_N_3408), .O(n27322));   // verilog/coms.v(118[11:12])
    defparam i16264_4_lut.LUT_INIT = 16'he420;
    SB_LUT4 i2_3_lut_4_lut_adj_1341 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(n26028), .I3(\data_in_frame[14] [0]), .O(n25895));   // verilog/coms.v(88[17:28])
    defparam i2_3_lut_4_lut_adj_1341.LUT_INIT = 16'h6996;
    SB_LUT4 i47040_2_lut (.I0(n66774), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n63159));
    defparam i47040_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48297_3_lut (.I0(n66888), .I1(n66552), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n65359));
    defparam i48297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11670_3_lut (.I0(\data_out_frame[1][7] ), .I1(\data_out_frame[3][7] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n27513));   // verilog/coms.v(109[34:55])
    defparam i11670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48301_3_lut (.I0(n66672), .I1(n66654), .I2(byte_transmit_counter[1]), 
            .I3(GND_net), .O(n65363));
    defparam i48301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11793_2_lut (.I0(byte_transmit_counter[1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n27637));   // verilog/coms.v(109[34:55])
    defparam i11793_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i43014_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60076));
    defparam i43014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43015_4_lut (.I0(n60076), .I1(n27637), .I2(byte_transmit_counter[2]), 
            .I3(\data_out_frame[1][5] ), .O(n60077));
    defparam i43015_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i43013_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60075));
    defparam i43013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1342 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(n58045), .I3(GND_net), .O(n55730));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_3_lut_adj_1342.LUT_INIT = 16'h6969;
    SB_LUT4 i46355_2_lut (.I0(n66780), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n63112));
    defparam i46355_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i48303_3_lut (.I0(n66768), .I1(n66624), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n65365));
    defparam i48303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_787_Select_221_i3_4_lut (.I0(\data_out_frame[25] [3]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n55959), .I3(\data_out_frame[25] [4]), 
            .O(n3_adj_5407));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_221_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i2_2_lut_adj_1343 (.I0(\FRAME_MATCHER.i [23]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5563));   // verilog/coms.v(157[7:23])
    defparam i2_2_lut_adj_1343.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1344 (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i[5] ), 
            .I2(\FRAME_MATCHER.i [6]), .I3(\FRAME_MATCHER.i [8]), .O(n14_adj_5564));   // verilog/coms.v(157[7:23])
    defparam i6_4_lut_adj_1344.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1345 (.I0(\FRAME_MATCHER.i [10]), .I1(n14_adj_5564), 
            .I2(n10_adj_5563), .I3(\FRAME_MATCHER.i [26]), .O(n58083));   // verilog/coms.v(157[7:23])
    defparam i7_4_lut_adj_1345.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1346 (.I0(\FRAME_MATCHER.i [15]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [28]), .I3(\FRAME_MATCHER.i [16]), .O(n30_adj_5565));   // verilog/coms.v(157[7:23])
    defparam i11_4_lut_adj_1346.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1347 (.I0(\FRAME_MATCHER.i [17]), .I1(n30_adj_5565), 
            .I2(\FRAME_MATCHER.i [13]), .I3(n58083), .O(n34));   // verilog/coms.v(157[7:23])
    defparam i15_4_lut_adj_1347.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1348 (.I0(\FRAME_MATCHER.i [20]), .I1(\FRAME_MATCHER.i [22]), 
            .I2(\FRAME_MATCHER.i [14]), .I3(\FRAME_MATCHER.i [29]), .O(n32_adj_5566));   // verilog/coms.v(157[7:23])
    defparam i13_4_lut_adj_1348.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(\FRAME_MATCHER.i [18]), .I1(\FRAME_MATCHER.i [24]), 
            .I2(\FRAME_MATCHER.i [30]), .I3(\FRAME_MATCHER.i [21]), .O(n33));   // verilog/coms.v(157[7:23])
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1349 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(\FRAME_MATCHER.i [9]), .I3(\FRAME_MATCHER.i [12]), .O(n31_c));   // verilog/coms.v(157[7:23])
    defparam i12_4_lut_adj_1349.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(n31_c), .I1(n33), .I2(n32_adj_5566), .I3(n34), 
            .O(n25087));   // verilog/coms.v(157[7:23])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22654_4_lut (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n25087), .I3(\FRAME_MATCHER.i[4] ), .O(n4452));   // verilog/coms.v(262[9:58])
    defparam i22654_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i468_2_lut (.I0(n4452), .I1(\FRAME_MATCHER.i_31__N_2514 ), .I2(GND_net), 
            .I3(GND_net), .O(n2076));   // verilog/coms.v(148[4] 304[11])
    defparam i468_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13374_3_lut_4_lut (.I0(n8), .I1(n55145), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n29219));
    defparam i13374_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13377_3_lut_4_lut (.I0(n8), .I1(n55145), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n29222));
    defparam i13377_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13380_3_lut_4_lut (.I0(n8), .I1(n55145), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n29225));
    defparam i13380_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_220_i3_4_lut (.I0(n50946), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n55886), .I3(n51134), .O(n3_adj_5406));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_220_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 select_787_Select_219_i3_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n6_adj_5567), .I3(\data_out_frame[25] [2]), 
            .O(n3_adj_5405));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_219_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 select_787_Select_218_i3_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n55896), .I3(n51146), .O(n3_adj_5404));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_218_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i6_4_lut_adj_1350 (.I0(n25648), .I1(n50221), .I2(n56103), 
            .I3(n55793), .O(n16_adj_5568));
    defparam i6_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1351 (.I0(n50685), .I1(n56088), .I2(n56231), 
            .I3(\data_out_frame[22] [6]), .O(n17_adj_5569));
    defparam i7_4_lut_adj_1351.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1352 (.I0(\data_out_frame[23] [0]), .I1(n17_adj_5569), 
            .I2(n15_adj_5570), .I3(n16_adj_5568), .O(n51146));
    defparam i1_4_lut_adj_1352.LUT_INIT = 16'h9669;
    SB_LUT4 i13383_3_lut_4_lut (.I0(n8), .I1(n55145), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n29228));
    defparam i13383_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1353 (.I0(n56201), .I1(n50685), .I2(n24633), 
            .I3(n56097), .O(n15_adj_5571));
    defparam i6_4_lut_adj_1353.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1354 (.I0(n15_adj_5571), .I1(n55707), .I2(n14_adj_5572), 
            .I3(n50187), .O(n51134));
    defparam i8_4_lut_adj_1354.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1355 (.I0(n50946), .I1(n51378), .I2(n56162), 
            .I3(GND_net), .O(n55959));
    defparam i1_3_lut_adj_1355.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1356 (.I0(n51134), .I1(n56249), .I2(n56165), 
            .I3(n51146), .O(n55823));
    defparam i3_4_lut_adj_1356.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_3_lut_3_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(reset), 
            .I3(GND_net), .O(n22318));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_3_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 select_787_Select_217_i3_4_lut (.I0(n51156), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n8_adj_5573), .I3(n55844), .O(n3_adj_5403));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_217_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i2_2_lut_adj_1357 (.I0(n50377), .I1(\data_out_frame[22] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5574));
    defparam i2_2_lut_adj_1357.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1358 (.I0(\data_out_frame[25] [0]), .I1(\data_out_frame[24] [6]), 
            .I2(n6_adj_5574), .I3(n51282), .O(n55896));
    defparam i2_4_lut_adj_1358.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1359 (.I0(\data_out_frame[25] [4]), .I1(\data_out_frame[25] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n56243));
    defparam i1_2_lut_adj_1359.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1360 (.I0(\data_out_frame[25] [2]), .I1(\data_out_frame[25] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n55886));
    defparam i1_2_lut_adj_1360.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1361 (.I0(n56135), .I1(n55878), .I2(n50377), 
            .I3(n56243), .O(n10_adj_5575));
    defparam i4_4_lut_adj_1361.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_215_i3_4_lut (.I0(\data_out_frame[25] [0]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n6_adj_5576), .I3(n23288), 
            .O(n3_adj_5401));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_215_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 select_787_Select_214_i3_4_lut (.I0(n23288), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n55714), .I3(n24672), .O(n3_adj_5400));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_214_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i13386_3_lut_4_lut (.I0(n8), .I1(n55145), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n29231));
    defparam i13386_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11668_3_lut (.I0(\data_out_frame[1][6] ), .I1(\data_out_frame[3][6] ), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n27511));   // verilog/coms.v(109[34:55])
    defparam i11668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43017_3_lut (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[7] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60079));
    defparam i43017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43018_4_lut (.I0(n60079), .I1(n27511), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n60080));
    defparam i43018_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i43016_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60078));
    defparam i43016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13389_3_lut_4_lut (.I0(n8), .I1(n55145), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n29234));
    defparam i13389_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13392_3_lut_4_lut (.I0(n8), .I1(n55145), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n29237));
    defparam i13392_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13395_3_lut_4_lut (.I0(n8), .I1(n55145), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n29240));
    defparam i13395_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i47881_3_lut (.I0(n66864), .I1(n66618), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n64943));
    defparam i47881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1362 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(\data_in_frame[18] [3]), .I3(GND_net), .O(n56138));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1362.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1363 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(n50264), .I3(n56183), .O(n55775));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1363.LUT_INIT = 16'h6996;
    SB_LUT4 i14009_3_lut_4_lut (.I0(n8_adj_5430), .I1(n55507), .I2(rx_data[2]), 
            .I3(\data_in_frame[1]_c [2]), .O(n29854));
    defparam i14009_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12060_3_lut_4_lut (.I0(n8_adj_5577), .I1(reset), .I2(n10_c), 
            .I3(n56368), .O(n27904));
    defparam i12060_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 equal_307_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(GND_net), .O(n8_adj_5577));   // verilog/coms.v(157[7:23])
    defparam equal_307_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i1_2_lut_3_lut_adj_1364 (.I0(\data_in_frame[16] [4]), .I1(n50260), 
            .I2(n55648), .I3(GND_net), .O(n50310));
    defparam i1_2_lut_3_lut_adj_1364.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_213_i3_4_lut (.I0(\data_out_frame[24] [3]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n55965), .I3(\data_out_frame[24] [4]), 
            .O(n3_adj_5399));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_213_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 equal_314_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i[3] ), .I1(\FRAME_MATCHER.i[4] ), 
            .I2(\FRAME_MATCHER.i[5] ), .I3(GND_net), .O(n10_c));   // verilog/coms.v(157[7:23])
    defparam equal_314_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 select_787_Select_212_i3_4_lut (.I0(n57163), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n55551), .I3(n57177), .O(n3_adj_5398));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_212_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i14012_3_lut_4_lut (.I0(n8_adj_5430), .I1(n55507), .I2(rx_data[3]), 
            .I3(\data_in_frame[1]_c [3]), .O(n29857));
    defparam i14012_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_1745_Select_0_i1_2_lut (.I0(tx_transmit_N_3416), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5511));   // verilog/coms.v(148[4] 304[11])
    defparam select_1745_Select_0_i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_787_Select_211_i3_4_lut (.I0(\data_out_frame[24] [2]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n55902), .I3(\data_out_frame[24] [1]), 
            .O(n3_adj_5397));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_211_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i4_4_lut_adj_1365 (.I0(n58178), .I1(\data_out_frame[21] [6]), 
            .I2(n50266), .I3(n55855), .O(n10_adj_5578));
    defparam i4_4_lut_adj_1365.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_210_i3_4_lut (.I0(n51154), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n10_adj_5578), .I3(\data_out_frame[24] [0]), .O(n3_adj_5396));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_210_i3_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i42732_3_lut_4_lut (.I0(n25933), .I1(\data_in_frame[0]_c [0]), 
            .I2(\data_in_frame[2] [0]), .I3(Kp_23__N_748), .O(n59783));
    defparam i42732_3_lut_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 select_787_Select_54_i2_4_lut (.I0(\data_out_frame[6] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[22] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5395));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_54_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i39359_2_lut_3_lut (.I0(n3484), .I1(\FRAME_MATCHER.i[5] ), .I2(n73), 
            .I3(GND_net), .O(n56366));
    defparam i39359_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[20] [4]), 
            .I2(n51265), .I3(n55823), .O(n6_adj_5567));
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1366 (.I0(n57163), .I1(n24672), .I2(GND_net), 
            .I3(GND_net), .O(n55965));
    defparam i1_2_lut_adj_1366.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1367 (.I0(\data_out_frame[22] [2]), .I1(n56234), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5579));
    defparam i1_2_lut_adj_1367.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1368 (.I0(\FRAME_MATCHER.i[4] ), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(\FRAME_MATCHER.i[3] ), 
            .O(n73));   // verilog/coms.v(156[9:50])
    defparam i2_3_lut_4_lut_adj_1368.LUT_INIT = 16'h0008;
    SB_LUT4 i1_4_lut_adj_1369 (.I0(DE_c), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(n6_adj_5580), .I3(\FRAME_MATCHER.i_31__N_2512 ), .O(n26520));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1369.LUT_INIT = 16'haaa8;
    SB_LUT4 i4_4_lut_adj_1370 (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[17] [6]), 
            .I2(n50388), .I3(n6_adj_5579), .O(n55572));
    defparam i4_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1371 (.I0(\data_out_frame[21] [7]), .I1(\data_out_frame[22] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5581));
    defparam i1_2_lut_adj_1371.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1372 (.I0(n55572), .I1(n55861), .I2(n51282), 
            .I3(n6_adj_5581), .O(n55784));
    defparam i4_4_lut_adj_1372.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_49746 (.I0(byte_transmit_counter_c[3]), 
            .I1(n65365), .I2(n63112), .I3(byte_transmit_counter_c[4]), 
            .O(n66855));
    defparam byte_transmit_counter_3__bdd_4_lut_49746.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_adj_1373 (.I0(\data_out_frame[23] [7]), .I1(\data_out_frame[23] [6]), 
            .I2(\data_out_frame[24] [1]), .I3(GND_net), .O(n55855));
    defparam i2_3_lut_adj_1373.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1374 (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[22] [3]), 
            .I2(n50004), .I3(GND_net), .O(n50410));
    defparam i2_3_lut_adj_1374.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1375 (.I0(\data_out_frame[20] [7]), .I1(n51197), 
            .I2(n51378), .I3(n51161), .O(n12_adj_5582));
    defparam i5_4_lut_adj_1375.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1376 (.I0(\data_in_frame[0]_c [3]), .I1(\data_in_frame[0]_c [2]), 
            .I2(\data_in_frame[2]_c [4]), .I3(n25908), .O(n50165));
    defparam i1_2_lut_3_lut_4_lut_adj_1376.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1377 (.I0(\data_out_frame[21] [1]), .I1(n12_adj_5582), 
            .I2(n55799), .I3(n51296), .O(n57678));
    defparam i6_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1378 (.I0(\data_out_frame[22] [6]), .I1(n57257), 
            .I2(GND_net), .I3(GND_net), .O(n56249));
    defparam i1_2_lut_adj_1378.LUT_INIT = 16'h9999;
    SB_LUT4 i12082_3_lut_4_lut (.I0(n8_adj_5430), .I1(reset), .I2(n3484), 
            .I3(n37097), .O(n27926));
    defparam i12082_3_lut_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_adj_1379 (.I0(\data_out_frame[24] [2]), .I1(\data_out_frame[24] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n55551));
    defparam i1_2_lut_adj_1379.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1380 (.I0(\data_out_frame[22] [7]), .I1(\data_out_frame[21] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n56097));
    defparam i1_2_lut_adj_1380.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1381 (.I0(n51150), .I1(n50179), .I2(\data_in_frame[19]_c [6]), 
            .I3(n57531), .O(n55932));
    defparam i1_3_lut_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i13140_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n27902), 
            .I3(GND_net), .O(n28985));   // verilog/coms.v(130[12] 305[6])
    defparam i13140_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut_adj_1382 (.I0(n51150), .I1(n50179), .I2(n57445), 
            .I3(GND_net), .O(n51173));
    defparam i1_2_lut_3_lut_adj_1382.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1383 (.I0(\data_in_frame[13] [5]), .I1(n55917), 
            .I2(\data_in_frame[15] [1]), .I3(n55730), .O(n56147));
    defparam i2_3_lut_4_lut_adj_1383.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1384 (.I0(\data_out_frame[24] [5]), .I1(\data_out_frame[24] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n55714));
    defparam i1_2_lut_adj_1384.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1385 (.I0(\data_out_frame[20] [6]), .I1(n24633), 
            .I2(\data_out_frame[20] [5]), .I3(GND_net), .O(n50221));
    defparam i2_3_lut_adj_1385.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1386 (.I0(\data_out_frame[20] [4]), .I1(n51265), 
            .I2(GND_net), .I3(GND_net), .O(n51376));
    defparam i1_2_lut_adj_1386.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1387 (.I0(n51210), .I1(n50266), .I2(\data_out_frame[23] [5]), 
            .I3(GND_net), .O(n57923));
    defparam i2_3_lut_adj_1387.LUT_INIT = 16'h6969;
    SB_LUT4 i6_2_lut (.I0(\data_out_frame[24] [6]), .I1(\data_out_frame[23] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n29_c));
    defparam i6_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14_4_lut_adj_1388 (.I0(n56165), .I1(n55714), .I2(n55935), 
            .I3(\data_out_frame[23] [1]), .O(n37));
    defparam i14_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1389 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[6] [2]), .I3(\data_out_frame[6] [1]), .O(n25239));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1389.LUT_INIT = 16'h6996;
    SB_LUT4 i18276_3_lut (.I0(n27902), .I1(rx_data[0]), .I2(\data_in_frame[5] [0]), 
            .I3(GND_net), .O(n28979));   // verilog/coms.v(94[13:20])
    defparam i18276_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13_4_lut_adj_1390 (.I0(n56097), .I1(n55551), .I2(n55952), 
            .I3(\data_out_frame[23] [5]), .O(n36));
    defparam i13_4_lut_adj_1390.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut (.I0(n37), .I1(n29_c), .I2(n51376), .I3(n50221), 
            .O(n42));
    defparam i19_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i13220_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in[3] [7]), .O(n29065));   // verilog/coms.v(130[12] 305[6])
    defparam i13220_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13089_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [0]), 
            .I3(\data_in[0] [0]), .O(n28934));   // verilog/coms.v(130[12] 305[6])
    defparam i13089_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i17_4_lut (.I0(n56129), .I1(\data_out_frame[20] [1]), .I2(n56249), 
            .I3(n57678), .O(n40));
    defparam i17_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i18_4_lut_adj_1391 (.I0(n50410), .I1(n36), .I2(n55855), .I3(\data_out_frame[23] [4]), 
            .O(n41));
    defparam i18_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 i13221_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in[3] [6]), .O(n29066));   // verilog/coms.v(130[12] 305[6])
    defparam i13221_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13222_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in[3] [5]), .O(n29067));   // verilog/coms.v(130[12] 305[6])
    defparam i13222_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16_4_lut_adj_1392 (.I0(n55784), .I1(n55790), .I2(\data_out_frame[22] [5]), 
            .I3(n56177), .O(n39));
    defparam i16_4_lut_adj_1392.LUT_INIT = 16'h6996;
    SB_LUT4 i13223_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in[3] [4]), .O(n29068));   // verilog/coms.v(130[12] 305[6])
    defparam i13223_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_787_Select_144_i2_4_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5532));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_144_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i22_4_lut (.I0(n39), .I1(n41), .I2(n40), .I3(n42), .O(n51237));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13350_3_lut_4_lut (.I0(n8_adj_5430), .I1(n55145), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n29195));
    defparam i13350_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13224_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in[3] [3]), .O(n29069));   // verilog/coms.v(130[12] 305[6])
    defparam i13224_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13225_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in[3] [2]), .O(n29070));   // verilog/coms.v(130[12] 305[6])
    defparam i13225_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i49199_3_lut (.I0(rx_data[6]), .I1(\data_in_frame[4] [6]), .I2(n27900), 
            .I3(GND_net), .O(n54747));   // verilog/coms.v(94[13:20])
    defparam i49199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1393 (.I0(n55710), .I1(n56150), .I2(n58113), 
            .I3(\data_out_frame[13] [6]), .O(n10_adj_5583));
    defparam i4_4_lut_adj_1393.LUT_INIT = 16'h9669;
    SB_LUT4 i11_3_lut_adj_1394 (.I0(rx_data[5]), .I1(\data_in_frame[4] [5]), 
            .I2(n27900), .I3(GND_net), .O(n54819));   // verilog/coms.v(94[13:20])
    defparam i11_3_lut_adj_1394.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1395 (.I0(n55949), .I1(n55920), .I2(n10_adj_5583), 
            .I3(\data_out_frame[15] [7]), .O(n51302));
    defparam i2_4_lut_adj_1395.LUT_INIT = 16'h6996;
    SB_LUT4 i13226_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in[3] [1]), .O(n29071));   // verilog/coms.v(130[12] 305[6])
    defparam i13226_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13227_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in[3] [0]), .O(n29072));   // verilog/coms.v(130[12] 305[6])
    defparam i13227_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13228_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [7]), 
            .I3(\data_in[2] [7]), .O(n29073));   // verilog/coms.v(130[12] 305[6])
    defparam i13228_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13229_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [6]), 
            .I3(\data_in[2] [6]), .O(n29074));   // verilog/coms.v(130[12] 305[6])
    defparam i13229_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13353_3_lut_4_lut (.I0(n8_adj_5430), .I1(n55145), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n29198));
    defparam i13353_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13230_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [5]), 
            .I3(\data_in[2] [5]), .O(n29075));   // verilog/coms.v(130[12] 305[6])
    defparam i13230_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13231_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [4]), 
            .I3(\data_in[2] [4]), .O(n29076));   // verilog/coms.v(130[12] 305[6])
    defparam i13231_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13232_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [3]), 
            .I3(\data_in[2] [3]), .O(n29077));   // verilog/coms.v(130[12] 305[6])
    defparam i13232_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13233_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [2]), 
            .I3(\data_in[2] [2]), .O(n29078));   // verilog/coms.v(130[12] 305[6])
    defparam i13233_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13234_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [1]), 
            .I3(\data_in[2] [1]), .O(n29079));   // verilog/coms.v(130[12] 305[6])
    defparam i13234_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5_4_lut_adj_1396 (.I0(n51261), .I1(n55717), .I2(\data_out_frame[19] [7]), 
            .I3(\data_out_frame[15] [3]), .O(n12_adj_5584));
    defparam i5_4_lut_adj_1396.LUT_INIT = 16'h6996;
    SB_LUT4 i13235_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[3] [0]), 
            .I3(\data_in[2] [0]), .O(n29080));   // verilog/coms.v(130[12] 305[6])
    defparam i13235_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13236_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [7]), 
            .I3(\data_in[1] [7]), .O(n29081));   // verilog/coms.v(130[12] 305[6])
    defparam i13236_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13356_3_lut_4_lut (.I0(n8_adj_5430), .I1(n55145), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n29201));
    defparam i13356_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13237_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [6]), 
            .I3(\data_in[1] [6]), .O(n29082));   // verilog/coms.v(130[12] 305[6])
    defparam i13237_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13359_3_lut_4_lut (.I0(n8_adj_5430), .I1(n55145), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n29204));
    defparam i13359_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13238_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [5]), 
            .I3(\data_in[1] [5]), .O(n29083));   // verilog/coms.v(130[12] 305[6])
    defparam i13238_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13239_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [4]), .O(n29084));   // verilog/coms.v(130[12] 305[6])
    defparam i13239_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13240_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [3]), 
            .I3(\data_in[1] [3]), .O(n29085));   // verilog/coms.v(130[12] 305[6])
    defparam i13240_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13241_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [2]), .O(n29086));   // verilog/coms.v(130[12] 305[6])
    defparam i13241_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_1397 (.I0(\data_out_frame[17] [5]), .I1(n12_adj_5584), 
            .I2(n56081), .I3(\data_out_frame[18] [0]), .O(n50004));
    defparam i6_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_LUT4 i13242_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [1]), 
            .I3(\data_in[1] [1]), .O(n29087));   // verilog/coms.v(130[12] 305[6])
    defparam i13242_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13243_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[2] [0]), 
            .I3(\data_in[1] [0]), .O(n29088));   // verilog/coms.v(130[12] 305[6])
    defparam i13243_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1398 (.I0(\data_out_frame[21] [6]), .I1(n56252), 
            .I2(GND_net), .I3(GND_net), .O(n55790));
    defparam i1_2_lut_adj_1398.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1399 (.I0(\data_out_frame[17] [7]), .I1(n26368), 
            .I2(GND_net), .I3(GND_net), .O(n56150));
    defparam i2_2_lut_adj_1399.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1400 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n55145), .O(n55152));
    defparam i1_2_lut_3_lut_4_lut_adj_1400.LUT_INIT = 16'hff7f;
    SB_LUT4 i13250_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [1]), 
            .I3(\data_in[0] [1]), .O(n29095));   // verilog/coms.v(130[12] 305[6])
    defparam i13250_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13249_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [2]), 
            .I3(\data_in[0] [2]), .O(n29094));   // verilog/coms.v(130[12] 305[6])
    defparam i13249_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13248_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [3]), 
            .I3(\data_in[0] [3]), .O(n29093));   // verilog/coms.v(130[12] 305[6])
    defparam i13248_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1401 (.I0(\data_out_frame[19] [0]), .I1(n51140), 
            .I2(GND_net), .I3(GND_net), .O(n55799));
    defparam i1_2_lut_adj_1401.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1402 (.I0(LED_c), .I1(LED_N_3408), .I2(GND_net), 
            .I3(GND_net), .O(n27_c));
    defparam i1_2_lut_adj_1402.LUT_INIT = 16'heeee;
    SB_LUT4 i13247_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [4]), 
            .I3(\data_in[0] [4]), .O(n29092));   // verilog/coms.v(130[12] 305[6])
    defparam i13247_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13246_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [5]), 
            .I3(\data_in[0] [5]), .O(n29091));   // verilog/coms.v(130[12] 305[6])
    defparam i13246_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n66855_bdd_4_lut (.I0(n66855), .I1(n66642), .I2(n7_adj_5585), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[5]));
    defparam n66855_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1403 (.I0(\data_out_frame[19] [6]), .I1(n25271), 
            .I2(n50298), .I3(n6_adj_5586), .O(n56234));   // verilog/coms.v(79[16:43])
    defparam i4_4_lut_adj_1403.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1404 (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[18] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n55949));
    defparam i1_2_lut_adj_1404.LUT_INIT = 16'h6666;
    SB_LUT4 i13245_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [6]), 
            .I3(\data_in[0] [6]), .O(n29090));   // verilog/coms.v(130[12] 305[6])
    defparam i13245_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i17_4_lut_adj_1405 (.I0(n50391), .I1(\data_out_frame[14] [3]), 
            .I2(n25385), .I3(n55763), .O(n42_adj_5587));
    defparam i17_4_lut_adj_1405.LUT_INIT = 16'h6996;
    SB_LUT4 i19064_3_lut (.I0(current_limit[8]), .I1(\data_in_frame[20] [0]), 
            .I2(n22318), .I3(GND_net), .O(n29639));
    defparam i19064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16260_4_lut (.I0(Kp_23__N_1748), .I1(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2509 ), .I3(LED_c), .O(n32103));   // verilog/coms.v(118[11:12])
    defparam i16260_4_lut.LUT_INIT = 16'hfac0;
    SB_LUT4 i18944_3_lut (.I0(current_limit[6]), .I1(\data_in_frame[21]_c [6]), 
            .I2(n22318), .I3(GND_net), .O(n29641));
    defparam i18944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13244_3_lut_4_lut_4_lut (.I0(rx_data_ready), .I1(reset), .I2(\data_in[1] [7]), 
            .I3(\data_in[0] [7]), .O(n29089));   // verilog/coms.v(130[12] 305[6])
    defparam i13244_3_lut_4_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13362_3_lut_4_lut (.I0(n8_adj_5430), .I1(n55145), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n29207));
    defparam i13362_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15_4_lut_adj_1406 (.I0(n50229), .I1(\data_out_frame[19] [4]), 
            .I2(\data_out_frame[18] [7]), .I3(n56109), .O(n40_adj_5588));
    defparam i15_4_lut_adj_1406.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1407 (.I0(n55805), .I1(\data_out_frame[14] [4]), 
            .I2(n55710), .I3(n50372), .O(n41_adj_5589));
    defparam i16_4_lut_adj_1407.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1408 (.I0(n55949), .I1(n56234), .I2(\data_out_frame[17] [7]), 
            .I3(n55778), .O(n39_adj_5590));
    defparam i14_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i21026_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1]_c [3]), 
            .I2(n22318), .I3(GND_net), .O(n29651));
    defparam i21026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31782_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1]_c [2]), 
            .I2(n22318), .I3(GND_net), .O(n29652));
    defparam i31782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31777_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1]_c [1]), 
            .I2(n22318), .I3(GND_net), .O(n29653));
    defparam i31777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_2_lut (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5591));
    defparam i12_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i23_4_lut (.I0(n39_adj_5590), .I1(n41_adj_5589), .I2(n40_adj_5588), 
            .I3(n42_adj_5587), .O(n48));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21244_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n22369), .I3(GND_net), .O(n29663));
    defparam i21244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18_4_lut_adj_1409 (.I0(n51219), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [5]), .I3(\data_out_frame[17] [4]), 
            .O(n43));
    defparam i18_4_lut_adj_1409.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut (.I0(n43), .I1(n48), .I2(n37_adj_5591), .I3(n38), 
            .O(n50927));
    defparam i24_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1410 (.I0(n26337), .I1(n50927), .I2(GND_net), 
            .I3(GND_net), .O(n56103));
    defparam i1_2_lut_adj_1410.LUT_INIT = 16'h6666;
    SB_LUT4 i18343_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6]_c [5]), 
            .I2(n22369), .I3(GND_net), .O(n29672));
    defparam i18343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut_adj_1411 (.I0(\data_out_frame[19] [5]), .I1(\data_out_frame[17] [0]), 
            .I2(n25687), .I3(n56103), .O(n18_adj_5592));
    defparam i7_4_lut_adj_1411.LUT_INIT = 16'h6996;
    SB_LUT4 i43085_3_lut (.I0(\data_out_frame[8][2] ), .I1(\data_out_frame[9] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60147));
    defparam i43085_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i43086_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n60148));
    defparam i43086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42927_3_lut (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n59989));
    defparam i42927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42926_3_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n59988));
    defparam i42926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_4_lut_adj_1412 (.I0(n50183), .I1(n18_adj_5592), .I2(n57868), 
            .I3(n55799), .O(n20_adj_5593));
    defparam i9_4_lut_adj_1412.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1413 (.I0(n57829), .I1(n56177), .I2(n51210), 
            .I3(n50266), .O(n56129));
    defparam i2_3_lut_4_lut_adj_1413.LUT_INIT = 16'h6996;
    SB_LUT4 i13365_3_lut_4_lut (.I0(n8_adj_5430), .I1(n55145), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n29210));
    defparam i13365_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_adj_1414 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[16] [4]), .I3(GND_net), .O(n7_adj_5594));   // verilog/coms.v(88[17:28])
    defparam i2_2_lut_3_lut_adj_1414.LUT_INIT = 16'h9696;
    SB_LUT4 i10_4_lut_adj_1415 (.I0(n15_adj_5595), .I1(n20_adj_5593), .I2(n51296), 
            .I3(\data_out_frame[16] [6]), .O(n50187));
    defparam i10_4_lut_adj_1415.LUT_INIT = 16'h9669;
    SB_LUT4 i13368_3_lut_4_lut (.I0(n8_adj_5430), .I1(n55145), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n29213));
    defparam i13368_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1416 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n25803));
    defparam i1_2_lut_adj_1416.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1417 (.I0(\data_out_frame[10] [0]), .I1(n25642), 
            .I2(\data_out_frame[7] [6]), .I3(\data_out_frame[9] [7]), .O(n56189));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_4_lut_adj_1417.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_adj_1418 (.I0(n25246), .I1(n56030), .I2(n55609), 
            .I3(n56198), .O(n8_adj_5596));
    defparam i3_3_lut_4_lut_adj_1418.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n3484), .I3(\FRAME_MATCHER.i[0] ), .O(n55512));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'hdfff;
    SB_LUT4 i1_2_lut_3_lut_adj_1419 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[5] [5]), .I3(GND_net), .O(n55543));   // verilog/coms.v(74[16:62])
    defparam i1_2_lut_3_lut_adj_1419.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1420 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [5]), 
            .I2(\data_out_frame[6] [7]), .I3(n1168), .O(n55609));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_4_lut_adj_1420.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1421 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n25246));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1421.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1422 (.I0(n55554), .I1(\data_out_frame[12] [0]), 
            .I2(n10_adj_5597), .I3(n55543), .O(n50183));   // verilog/coms.v(74[16:27])
    defparam i5_3_lut_4_lut_adj_1422.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1423 (.I0(n50298), .I1(n25964), .I2(n50234), 
            .I3(GND_net), .O(n26123));
    defparam i1_2_lut_3_lut_adj_1423.LUT_INIT = 16'h9696;
    SB_LUT4 i3_2_lut_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(n26397), .I3(GND_net), .O(n17_adj_5598));   // verilog/coms.v(100[12:26])
    defparam i3_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1424 (.I0(\data_out_frame[6] [6]), .I1(n55735), 
            .I2(\data_out_frame[6] [7]), .I3(n1168), .O(n26397));
    defparam i1_2_lut_4_lut_adj_1424.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1425 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[7] [0]), 
            .I2(\data_out_frame[7] [1]), .I3(\data_out_frame[8][7] ), .O(n56213));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_4_lut_adj_1425.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1426 (.I0(\data_out_frame[8][2] ), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[5] [6]), .I3(GND_net), .O(n56126));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_1426.LUT_INIT = 16'h9696;
    SB_LUT4 i13371_3_lut_4_lut (.I0(n8_adj_5430), .I1(n55145), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n29216));
    defparam i13371_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1427 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n25385));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1427.LUT_INIT = 16'h6666;
    SB_LUT4 i11697_4_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(n133[0]), .I2(n3484), 
            .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n27541));   // verilog/coms.v(158[12:15])
    defparam i11697_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i1_2_lut_adj_1428 (.I0(\data_out_frame[16] [3]), .I1(n57868), 
            .I2(GND_net), .I3(GND_net), .O(n51197));
    defparam i1_2_lut_adj_1428.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1429 (.I0(n25648), .I1(n55707), .I2(n50270), 
            .I3(GND_net), .O(n50685));
    defparam i2_3_lut_adj_1429.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1430 (.I0(\data_out_frame[18] [5]), .I1(n51197), 
            .I2(n51140), .I3(\data_out_frame[16] [4]), .O(n25648));
    defparam i3_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1431 (.I0(\data_out_frame[8][3] ), .I1(\data_out_frame[8][4] ), 
            .I2(\data_out_frame[5] [7]), .I3(GND_net), .O(n6_adj_5506));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1431.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1432 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[6] [2]), .I3(\data_out_frame[5] [5]), .O(n56240));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_4_lut_adj_1432.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_142_i2_4_lut (.I0(\data_out_frame[17] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5505));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_142_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1433 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[17] [0]), 
            .I2(n26439), .I3(GND_net), .O(n55738));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1433.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1434 (.I0(\data_out_frame[13] [7]), .I1(n56100), 
            .I2(n25642), .I3(\data_out_frame[5] [4]), .O(n12_adj_5599));
    defparam i5_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1435 (.I0(n26337), .I1(n56228), .I2(\data_out_frame[19] [4]), 
            .I3(n57849), .O(n57829));
    defparam i2_3_lut_4_lut_adj_1435.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_141_i2_4_lut (.I0(\data_out_frame[17] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5504));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_141_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_140_i2_4_lut (.I0(\data_out_frame[17] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5503));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_140_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i6_4_lut_adj_1436 (.I0(n50234), .I1(n12_adj_5599), .I2(\data_out_frame[14] [1]), 
            .I3(n55998), .O(n57868));
    defparam i6_4_lut_adj_1436.LUT_INIT = 16'h6996;
    SB_LUT4 i49198_3_lut (.I0(rx_data[4]), .I1(\data_in_frame[3] [4]), .I2(n27898), 
            .I3(GND_net), .O(n54743));   // verilog/coms.v(94[13:20])
    defparam i49198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1437 (.I0(n51330), .I1(n55908), .I2(n57868), 
            .I3(\data_out_frame[16] [2]), .O(n49936));
    defparam i3_4_lut_adj_1437.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1438 (.I0(\data_out_frame[18] [3]), .I1(n49936), 
            .I2(GND_net), .I3(GND_net), .O(n50341));
    defparam i1_2_lut_adj_1438.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1439 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(n50331), .I3(GND_net), .O(n51232));
    defparam i2_3_lut_adj_1439.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1440 (.I0(n56258), .I1(n56240), .I2(n58237), 
            .I3(n51261), .O(n6_adj_5600));
    defparam i1_2_lut_4_lut_adj_1440.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1441 (.I0(\data_in_frame[19]_c [3]), .I1(n56181), 
            .I2(n57531), .I3(\data_in_frame[21][5] ), .O(n55972));
    defparam i2_3_lut_4_lut_adj_1441.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_139_i2_4_lut (.I0(\data_out_frame[17] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5502));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_139_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1442 (.I0(n55884), .I1(n58122), .I2(GND_net), 
            .I3(GND_net), .O(n55710));
    defparam i1_2_lut_adj_1442.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_1443 (.I0(\data_in_frame[23]_c [7]), .I1(n56366), 
            .I2(n27939), .I3(rx_data[7]), .O(n54687));   // verilog/coms.v(94[13:20])
    defparam i11_4_lut_adj_1443.LUT_INIT = 16'hca0a;
    SB_LUT4 i3_4_lut_adj_1444 (.I0(\data_out_frame[18] [1]), .I1(n56225), 
            .I2(n55992), .I3(n55710), .O(n58154));
    defparam i3_4_lut_adj_1444.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut_adj_1445 (.I0(rx_data[2]), .I1(\data_in_frame[3] [2]), 
            .I2(n27898), .I3(GND_net), .O(n54803));   // verilog/coms.v(94[13:20])
    defparam i11_3_lut_adj_1445.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1446 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[10] [2]), 
            .I2(\data_out_frame[10] [3]), .I3(GND_net), .O(n56010));   // verilog/coms.v(88[17:63])
    defparam i1_2_lut_3_lut_adj_1446.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1447 (.I0(n50341), .I1(\data_out_frame[13] [6]), 
            .I2(n1835), .I3(n6_adj_5601), .O(n51265));
    defparam i4_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1448 (.I0(n57257), .I1(n25648), .I2(n55989), 
            .I3(\data_out_frame[18] [4]), .O(n26012));
    defparam i3_4_lut_adj_1448.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1449 (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[18] [4]), 
            .I2(\data_in_frame[22] [6]), .I3(n55672), .O(n57143));   // verilog/coms.v(81[16:27])
    defparam i2_3_lut_4_lut_adj_1449.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1450 (.I0(n51261), .I1(\data_out_frame[15] [3]), 
            .I2(n25271), .I3(GND_net), .O(n55778));
    defparam i2_3_lut_adj_1450.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1451 (.I0(n50298), .I1(n25964), .I2(n50234), 
            .I3(n55992), .O(n6_adj_5601));
    defparam i1_2_lut_3_lut_4_lut_adj_1451.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1452 (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[18] [4]), 
            .I2(\data_in_frame[18] [1]), .I3(GND_net), .O(n56159));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1452.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_138_i2_4_lut (.I0(\data_out_frame[17] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5501));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_138_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_4_lut_adj_1453 (.I0(\data_out_frame[6] [6]), .I1(n56198), 
            .I2(n56016), .I3(n55579), .O(n25271));   // verilog/coms.v(77[16:43])
    defparam i3_4_lut_adj_1453.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1454 (.I0(\data_out_frame[17] [4]), .I1(n55727), 
            .I2(n25271), .I3(n50249), .O(n50388));
    defparam i3_4_lut_adj_1454.LUT_INIT = 16'h6996;
    SB_LUT4 i23_3_lut_4_lut (.I0(n8_adj_4), .I1(n55145), .I2(\data_in_frame[8] [4]), 
            .I3(rx_data[4]), .O(n15_adj_5434));
    defparam i23_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 i3_4_lut_adj_1455 (.I0(n50229), .I1(n50388), .I2(\data_out_frame[22] [0]), 
            .I3(\data_out_frame[19] [6]), .O(n56252));
    defparam i3_4_lut_adj_1455.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_137_i2_4_lut (.I0(\data_out_frame[17] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5500));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_137_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13315_3_lut_4_lut (.I0(n8_adj_4), .I1(n55145), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n29160));
    defparam i13315_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1456 (.I0(\data_out_frame[21] [7]), .I1(n56252), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5602));
    defparam i1_2_lut_adj_1456.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1457 (.I0(n56177), .I1(n51154), .I2(\data_out_frame[23] [7]), 
            .I3(n6_adj_5602), .O(n58178));
    defparam i4_4_lut_adj_1457.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1458 (.I0(n57829), .I1(n50388), .I2(n57849), 
            .I3(\data_out_frame[19] [5]), .O(n51154));
    defparam i1_2_lut_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1459 (.I0(n26012), .I1(n51265), .I2(n58154), 
            .I3(GND_net), .O(n14_adj_5603));
    defparam i5_3_lut_adj_1459.LUT_INIT = 16'h6969;
    SB_LUT4 i6_4_lut_adj_1460 (.I0(n55790), .I1(n57829), .I2(n50270), 
            .I3(n50004), .O(n15_adj_5604));
    defparam i6_4_lut_adj_1460.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut_adj_1461 (.I0(n15_adj_5604), .I1(n51302), .I2(n14_adj_5603), 
            .I3(\data_out_frame[22] [1]), .O(n57177));
    defparam i8_4_lut_adj_1461.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_136_i2_4_lut (.I0(\data_out_frame[17] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5499));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_136_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1462 (.I0(n57177), .I1(n58178), .I2(GND_net), 
            .I3(GND_net), .O(n55902));
    defparam i1_2_lut_adj_1462.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_135_i2_4_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5498));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_135_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1463 (.I0(n50298), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[17] [7]), .I3(n26368), .O(n56225));
    defparam i1_2_lut_4_lut_adj_1463.LUT_INIT = 16'h6996;
    SB_LUT4 i23_3_lut_4_lut_adj_1464 (.I0(n8_adj_4), .I1(n55145), .I2(\data_in_frame[8] [2]), 
            .I3(rx_data[2]), .O(n15_adj_5433));
    defparam i23_3_lut_4_lut_adj_1464.LUT_INIT = 16'hf1e0;
    SB_LUT4 i13212_3_lut_4_lut (.I0(n8_adj_4), .I1(n55145), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n29057));
    defparam i13212_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1465 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[15] [7]), 
            .I2(\data_out_frame[13] [7]), .I3(n50331), .O(n51330));
    defparam i1_2_lut_4_lut_adj_1465.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_134_i2_4_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5497));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_134_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1466 (.I0(\data_out_frame[24] [0]), .I1(n51237), 
            .I2(n57923), .I3(GND_net), .O(n56135));
    defparam i2_3_lut_adj_1466.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1467 (.I0(n56135), .I1(n23288), .I2(n55902), 
            .I3(n51282), .O(n14_adj_5605));
    defparam i6_4_lut_adj_1467.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1468 (.I0(\data_out_frame[25] [7]), .I1(n55965), 
            .I2(n51237), .I3(\data_out_frame[22] [4]), .O(n13_adj_5606));
    defparam i5_4_lut_adj_1468.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_209_i3_3_lut (.I0(n13_adj_5606), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n14_adj_5605), .I3(GND_net), .O(n3_adj_5394));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_209_i3_3_lut.LUT_INIT = 16'h4848;
    SB_LUT4 select_787_Select_133_i2_4_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5496));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_133_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1469 (.I0(\data_out_frame[25] [7]), .I1(\data_out_frame[25] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n55878));
    defparam i1_2_lut_adj_1469.LUT_INIT = 16'h6666;
    SB_LUT4 i13209_3_lut_4_lut (.I0(n8_adj_4), .I1(n55145), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n29054));
    defparam i13209_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13341_3_lut_4_lut (.I0(n8_adj_4), .I1(n55145), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n29186));
    defparam i13341_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1470 (.I0(\data_out_frame[13] [0]), .I1(n55678), 
            .I2(\data_out_frame[17] [2]), .I3(n24677), .O(n56228));   // verilog/coms.v(79[16:43])
    defparam i3_4_lut_adj_1470.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1471 (.I0(n25996), .I1(n56010), .I2(\data_out_frame[10] [1]), 
            .I3(\data_out_frame[10] [6]), .O(n14_adj_5607));   // verilog/coms.v(88[17:63])
    defparam i6_4_lut_adj_1471.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1472 (.I0(\data_out_frame[10] [5]), .I1(n26092), 
            .I2(n57840), .I3(\data_out_frame[10] [7]), .O(n13_adj_5608));   // verilog/coms.v(88[17:63])
    defparam i5_4_lut_adj_1472.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1473 (.I0(n26378), .I1(n26187), .I2(n55606), 
            .I3(\data_out_frame[12] [7]), .O(n18_adj_5609));
    defparam i7_4_lut_adj_1473.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1474 (.I0(n13_adj_5608), .I1(n25642), .I2(n14_adj_5607), 
            .I3(n56195), .O(n17_adj_5610));
    defparam i6_4_lut_adj_1474.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut_adj_1475 (.I0(n56010), .I1(n25239), .I2(n25820), 
            .I3(n37_adj_5611), .O(n19_adj_5612));
    defparam i8_4_lut_adj_1475.LUT_INIT = 16'h6996;
    SB_LUT4 i10_3_lut (.I0(n19_adj_5612), .I1(n17_adj_5610), .I2(n18_adj_5609), 
            .I3(GND_net), .O(n51261));
    defparam i10_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i13344_3_lut_4_lut (.I0(n8_adj_4), .I1(n55145), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n29189));
    defparam i13344_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_49736 (.I0(byte_transmit_counter_c[3]), 
            .I1(n65363), .I2(n63131), .I3(byte_transmit_counter_c[4]), 
            .O(n66843));
    defparam byte_transmit_counter_3__bdd_4_lut_49736.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut_adj_1476 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(\data_out_frame[15] [1]), .I3(n6_adj_5600), .O(n57849));
    defparam i4_4_lut_adj_1476.LUT_INIT = 16'h6996;
    SB_LUT4 n66843_bdd_4_lut (.I0(n66843), .I1(n66606), .I2(n7_adj_5613), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[7]));
    defparam n66843_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1477 (.I0(n26337), .I1(n56228), .I2(GND_net), 
            .I3(GND_net), .O(n55751));
    defparam i1_2_lut_adj_1477.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1478 (.I0(\data_out_frame[21] [5]), .I1(n55751), 
            .I2(\data_out_frame[19] [3]), .I3(n56094), .O(n56177));
    defparam i3_4_lut_adj_1478.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1479 (.I0(\data_out_frame[17] [0]), .I1(n26439), 
            .I2(GND_net), .I3(GND_net), .O(n55763));
    defparam i1_2_lut_adj_1479.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1480 (.I0(\data_in_frame[19]_c [3]), 
            .I1(n58144), .I2(n55985), .I3(n32987), .O(n50305));
    defparam i1_2_lut_3_lut_4_lut_adj_1480.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1481 (.I0(n1516), .I1(n56123), .I2(n55630), .I3(\data_out_frame[14] [6]), 
            .O(n12_adj_5614));   // verilog/coms.v(88[17:63])
    defparam i5_4_lut_adj_1481.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1482 (.I0(\data_out_frame[12] [4]), .I1(n12_adj_5614), 
            .I2(\data_out_frame[12] [5]), .I3(n56240), .O(n26337));   // verilog/coms.v(88[17:63])
    defparam i6_4_lut_adj_1482.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1483 (.I0(n55995), .I1(\data_out_frame[10] [0]), 
            .I2(\data_out_frame[12] [3]), .I3(n56186), .O(n10_adj_5615));   // verilog/coms.v(77[16:27])
    defparam i4_4_lut_adj_1483.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1484 (.I0(\data_out_frame[9] [7]), .I1(n10_adj_5615), 
            .I2(\data_out_frame[5] [3]), .I3(GND_net), .O(n26439));   // verilog/coms.v(77[16:27])
    defparam i5_3_lut_adj_1484.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1485 (.I0(n26439), .I1(n50183), .I2(GND_net), 
            .I3(GND_net), .O(n51161));
    defparam i1_2_lut_adj_1485.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_132_i2_4_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5495));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_132_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13347_3_lut_4_lut (.I0(n8_adj_4), .I1(n55145), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n29192));
    defparam i13347_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1486 (.I0(\data_out_frame[16] [1]), .I1(n55738), 
            .I2(n55590), .I3(n26337), .O(n25687));   // verilog/coms.v(88[17:28])
    defparam i3_4_lut_adj_1486.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_49726 (.I0(byte_transmit_counter_c[3]), 
            .I1(n65359), .I2(n63159), .I3(byte_transmit_counter_c[4]), 
            .O(n66837));
    defparam byte_transmit_counter_3__bdd_4_lut_49726.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_4_lut_adj_1487 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[7] [7]), 
            .I2(n55606), .I3(n56126), .O(n58237));   // verilog/coms.v(75[16:27])
    defparam i3_4_lut_adj_1487.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1488 (.I0(n56258), .I1(n56240), .I2(n58237), 
            .I3(GND_net), .O(n50190));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1488.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1489 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [5]), 
            .I2(n25656), .I3(\data_out_frame[16] [7]), .O(n25494));   // verilog/coms.v(88[17:28])
    defparam i3_4_lut_adj_1489.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1490 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n55727));
    defparam i1_2_lut_adj_1490.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1491 (.I0(n25964), .I1(n26267), .I2(\data_out_frame[13] [7]), 
            .I3(\data_out_frame[13] [6]), .O(n55908));
    defparam i2_3_lut_4_lut_adj_1491.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1492 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n55678));
    defparam i1_2_lut_adj_1492.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1493 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n55717));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1493.LUT_INIT = 16'h6666;
    SB_LUT4 n66837_bdd_4_lut (.I0(n66837), .I1(n66804), .I2(n7_adj_5616), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[0]));
    defparam n66837_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_789_Select_0_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n1_adj_5514));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_0_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1047_2_lut (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1835));   // verilog/coms.v(74[16:27])
    defparam i1047_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_131_i2_4_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5494));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_131_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_adj_1494 (.I0(n25642), .I1(n55796), .I2(\data_out_frame[14] [0]), 
            .I3(GND_net), .O(n26267));
    defparam i2_3_lut_adj_1494.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1495 (.I0(n26267), .I1(n50234), .I2(n26368), 
            .I3(GND_net), .O(n50331));
    defparam i2_3_lut_adj_1495.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1496 (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[12] [5]), 
            .I2(\data_out_frame[10] [5]), .I3(GND_net), .O(n56258));
    defparam i2_3_lut_adj_1496.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1497 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n55498));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1497.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1498 (.I0(\data_out_frame[8][3] ), .I1(\data_out_frame[8][4] ), 
            .I2(GND_net), .I3(GND_net), .O(n56210));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1498.LUT_INIT = 16'h6666;
    SB_LUT4 select_789_Select_7_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(\byte_transmit_counter[7] ), 
            .I3(GND_net), .O(n1_adj_5417));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_7_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_adj_1499 (.I0(\data_out_frame[8][5] ), .I1(\data_out_frame[8][6] ), 
            .I2(GND_net), .I3(GND_net), .O(n56016));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1499.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1500 (.I0(n26187), .I1(\data_out_frame[4] [6]), 
            .I2(n56001), .I3(\data_out_frame[6] [4]), .O(n24_adj_5617));   // verilog/coms.v(100[12:26])
    defparam i10_4_lut_adj_1500.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_6_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(\byte_transmit_counter[6] ), 
            .I3(GND_net), .O(n1_adj_5416));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_6_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i8_4_lut_adj_1501 (.I0(\data_out_frame[8][2] ), .I1(\data_out_frame[4] [7]), 
            .I2(n55543), .I3(n55781), .O(n22_adj_5618));   // verilog/coms.v(100[12:26])
    defparam i8_4_lut_adj_1501.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1502 (.I0(n17_adj_5598), .I1(n24_adj_5617), .I2(n25239), 
            .I3(\data_out_frame[4] [4]), .O(n26_adj_5619));   // verilog/coms.v(100[12:26])
    defparam i12_4_lut_adj_1502.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_130_i2_4_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5493));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_130_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_789_Select_5_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(\byte_transmit_counter[5] ), 
            .I3(GND_net), .O(n1_adj_5415));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_5_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i13_4_lut_adj_1503 (.I0(n55864), .I1(n26_adj_5619), .I2(n22_adj_5618), 
            .I3(\data_out_frame[4] [5]), .O(n58238));   // verilog/coms.v(100[12:26])
    defparam i13_4_lut_adj_1503.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_2_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n1_adj_5412));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_2_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i10_4_lut_adj_1504 (.I0(\data_out_frame[9] [7]), .I1(n56016), 
            .I2(n25996), .I3(n56210), .O(n24_adj_5620));   // verilog/coms.v(77[16:43])
    defparam i10_4_lut_adj_1504.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1505 (.I0(n58238), .I1(\data_out_frame[9] [1]), 
            .I2(n56091), .I3(\data_out_frame[5] [4]), .O(n22_adj_5621));   // verilog/coms.v(77[16:43])
    defparam i8_4_lut_adj_1505.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1506 (.I0(\data_out_frame[9] [5]), .I1(n24_adj_5620), 
            .I2(n18_adj_5622), .I3(n56207), .O(n26_adj_5623));   // verilog/coms.v(77[16:43])
    defparam i12_4_lut_adj_1506.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_1_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter[1]), 
            .I3(GND_net), .O(n1));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_1_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 select_789_Select_3_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[3]), 
            .I3(GND_net), .O(n1_adj_5413));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_3_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i13_4_lut_adj_1507 (.I0(n56213), .I1(n26_adj_5623), .I2(n22_adj_5621), 
            .I3(n56053), .O(n57840));   // verilog/coms.v(77[16:43])
    defparam i13_4_lut_adj_1507.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1508 (.I0(n25964), .I1(n26267), .I2(n1699), 
            .I3(n25656), .O(n4));
    defparam i1_2_lut_4_lut_adj_1508.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1509 (.I0(\data_out_frame[13] [1]), .I1(n57840), 
            .I2(GND_net), .I3(GND_net), .O(n56195));
    defparam i1_2_lut_adj_1509.LUT_INIT = 16'h9999;
    SB_LUT4 select_787_Select_129_i2_4_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5492));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_129_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1510 (.I0(\data_out_frame[20] [0]), .I1(n50388), 
            .I2(n57849), .I3(\data_out_frame[19] [5]), .O(n55707));
    defparam i1_2_lut_4_lut_adj_1510.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1511 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26378));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1511.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1512 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(n50187), .I3(GND_net), .O(n55861));   // verilog/coms.v(81[16:27])
    defparam i1_2_lut_3_lut_adj_1512.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1513 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[8][4] ), .I3(n1130), .O(n10_adj_5625));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1513.LUT_INIT = 16'h6996;
    SB_LUT4 select_789_Select_4_i1_2_lut_3_lut (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.i_31__N_2511 ), .I2(byte_transmit_counter_c[4]), 
            .I3(GND_net), .O(n1_adj_5414));   // verilog/coms.v(148[4] 304[11])
    defparam select_789_Select_4_i1_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i2_3_lut_3_lut (.I0(\FRAME_MATCHER.i_31__N_2513 ), .I1(reset), 
            .I2(LED_N_3408), .I3(GND_net), .O(n22369));
    defparam i2_3_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i2_3_lut_adj_1514 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n26187));
    defparam i2_3_lut_adj_1514.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_49721 (.I0(byte_transmit_counter_c[3]), 
            .I1(n65357), .I2(n63135), .I3(byte_transmit_counter_c[4]), 
            .O(n66831));
    defparam byte_transmit_counter_3__bdd_4_lut_49721.LUT_INIT = 16'he4aa;
    SB_LUT4 select_787_Select_128_i2_4_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5491));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_128_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1515 (.I0(\data_out_frame[8][3] ), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n56123));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1515.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_151_i2_4_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5291));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_151_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_2_lut_adj_1516 (.I0(n56030), .I1(\data_out_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5626));   // verilog/coms.v(88[17:28])
    defparam i2_2_lut_adj_1516.LUT_INIT = 16'h6666;
    SB_LUT4 n66831_bdd_4_lut (.I0(n66831), .I1(n66678), .I2(n7_adj_5627), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[2]));
    defparam n66831_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1517 (.I0(n56123), .I1(\data_out_frame[10] [6]), 
            .I2(\data_out_frame[8][4] ), .I3(\data_out_frame[12] [6]), .O(n14_adj_5628));   // verilog/coms.v(88[17:28])
    defparam i6_4_lut_adj_1517.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1518 (.I0(n56126), .I1(n14_adj_5628), .I2(n10_adj_5626), 
            .I3(\data_out_frame[6] [0]), .O(n24677));   // verilog/coms.v(88[17:28])
    defparam i7_4_lut_adj_1518.LUT_INIT = 16'h6996;
    SB_LUT4 i12583_4_lut_4_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2513 ), 
            .I2(n26960), .I3(n27_c), .O(n28428));   // verilog/coms.v(130[12] 305[6])
    defparam i12583_4_lut_4_lut.LUT_INIT = 16'h5450;
    SB_LUT4 select_787_Select_127_i2_4_lut (.I0(\data_out_frame[15] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5490));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_127_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1519 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [5]), 
            .I2(\data_out_frame[19] [7]), .I3(GND_net), .O(n6_adj_5586));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1519.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1520 (.I0(n56056), .I1(\data_out_frame[11] [3]), 
            .I2(\data_out_frame[9] [3]), .I3(n56213), .O(n10_adj_5629));   // verilog/coms.v(88[17:28])
    defparam i4_4_lut_adj_1520.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1521 (.I0(\data_out_frame[13] [5]), .I1(n55662), 
            .I2(n10_adj_5629), .I3(\data_out_frame[9] [1]), .O(n26368));
    defparam i1_4_lut_adj_1521.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1522 (.I0(n25246), .I1(n56019), .I2(n55579), 
            .I3(n26397), .O(n1720));
    defparam i3_4_lut_adj_1522.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1523 (.I0(\data_out_frame[13] [0]), .I1(n24677), 
            .I2(GND_net), .I3(GND_net), .O(n50249));
    defparam i1_2_lut_adj_1523.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1524 (.I0(\data_out_frame[11] [4]), .I1(n26187), 
            .I2(GND_net), .I3(GND_net), .O(n56056));   // verilog/coms.v(88[17:28])
    defparam i1_2_lut_adj_1524.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_49716 (.I0(byte_transmit_counter_c[3]), 
            .I1(n65355), .I2(n63136), .I3(byte_transmit_counter_c[4]), 
            .O(n66825));
    defparam byte_transmit_counter_3__bdd_4_lut_49716.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1525 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n55873));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1525.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1526 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n55781));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1526.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1527 (.I0(n55554), .I1(\data_out_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n56100));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1527.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1528 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[17] [7]), 
            .I2(n26368), .I3(GND_net), .O(n56081));
    defparam i1_2_lut_3_lut_adj_1528.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1529 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5630));
    defparam i1_2_lut_adj_1529.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1530 (.I0(n55742), .I1(\data_out_frame[4] [7]), 
            .I2(n25661), .I3(n6_adj_5630), .O(n55796));
    defparam i4_4_lut_adj_1530.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_126_i2_4_lut (.I0(\data_out_frame[15] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5489));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_126_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i342_2_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1130));   // verilog/coms.v(79[16:27])
    defparam i342_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1531 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n56091));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1531.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1532 (.I0(\data_out_frame[11] [5]), .I1(n56091), 
            .I2(n55735), .I3(\data_out_frame[7] [1]), .O(n10_adj_5631));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1532.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1533 (.I0(n55742), .I1(n10_adj_5631), .I2(\data_out_frame[6] [7]), 
            .I3(GND_net), .O(n50234));   // verilog/coms.v(88[17:70])
    defparam i5_3_lut_adj_1533.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1534 (.I0(n25915), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[11] [4]), .I3(n25661), .O(n12_adj_5632));   // verilog/coms.v(88[17:70])
    defparam i5_4_lut_adj_1534.LUT_INIT = 16'h6996;
    SB_LUT4 i6_3_lut (.I0(\data_out_frame[9] [3]), .I1(n12_adj_5632), .I2(n17_adj_5598), 
            .I3(GND_net), .O(n25964));   // verilog/coms.v(88[17:70])
    defparam i6_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1535 (.I0(n25964), .I1(n50234), .I2(GND_net), 
            .I3(GND_net), .O(n55920));
    defparam i1_2_lut_adj_1535.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_125_i2_4_lut (.I0(\data_out_frame[15] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5488));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_125_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i911_2_lut (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1699));   // verilog/coms.v(74[16:27])
    defparam i911_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1536 (.I0(\data_out_frame[14] [2]), .I1(n56189), 
            .I2(n55796), .I3(\data_out_frame[12] [1]), .O(n10_adj_5597));   // verilog/coms.v(74[16:27])
    defparam i4_4_lut_adj_1536.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1537 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n55864));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1537.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1538 (.I0(\data_in_frame[13] [5]), .I1(n51256), 
            .I2(n51228), .I3(\data_in_frame[13] [4]), .O(n56171));
    defparam i1_2_lut_3_lut_4_lut_adj_1538.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_124_i2_4_lut (.I0(\data_out_frame[15] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5487));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_124_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1539 (.I0(n55181), .I1(n33_adj_5633), .I2(n105), 
            .I3(control_update), .O(n7064));
    defparam i2_3_lut_4_lut_adj_1539.LUT_INIT = 16'h2000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1540 (.I0(n55181), .I1(n33_adj_5633), 
            .I2(n38328), .I3(control_update), .O(n24981));
    defparam i1_2_lut_3_lut_4_lut_adj_1540.LUT_INIT = 16'h2fff;
    SB_LUT4 i22895_2_lut_3_lut_4_lut (.I0(n55181), .I1(n33_adj_5633), .I2(n38328), 
            .I3(control_update), .O(n38638));
    defparam i22895_2_lut_3_lut_4_lut.LUT_INIT = 16'hf2ff;
    SB_LUT4 i1_2_lut_adj_1541 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n55735));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1541.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1542 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[8][7] ), 
            .I2(GND_net), .I3(GND_net), .O(n56198));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1542.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1543 (.I0(\data_in_frame[0]_c [2]), .I1(\data_in_frame[0]_c [1]), 
            .I2(\data_in_frame[0]_c [3]), .I3(GND_net), .O(n6));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1543.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1544 (.I0(n25246), .I1(n56030), .I2(GND_net), 
            .I3(GND_net), .O(n25996));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_adj_1544.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1545 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n56207));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1545.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1546 (.I0(\data_in_frame[0]_c [2]), .I1(\data_in_frame[0]_c [1]), 
            .I2(\data_in_frame[2]_c [3]), .I3(GND_net), .O(n25908));   // verilog/coms.v(78[16:43])
    defparam i1_2_lut_3_lut_adj_1546.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1547 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[7] [1]), 
            .I2(\data_out_frame[8][7] ), .I3(GND_net), .O(n55636));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1547.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1548 (.I0(\data_out_frame[11] [2]), .I1(n37_adj_5611), 
            .I2(\data_out_frame[11] [3]), .I3(GND_net), .O(n56044));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_adj_1548.LUT_INIT = 16'h9696;
    SB_LUT4 n66825_bdd_4_lut (.I0(n66825), .I1(n66798), .I2(n7_adj_5635), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[1]));
    defparam n66825_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1549 (.I0(n56044), .I1(n55636), .I2(\data_out_frame[13] [4]), 
            .I3(n56207), .O(n10_adj_5636));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1549.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_123_i2_4_lut (.I0(\data_out_frame[15] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5486));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_123_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(74[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(n32100), .O(n6_adj_5580));   // verilog/coms.v(148[4] 304[11])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 equal_311_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8));   // verilog/coms.v(157[7:23])
    defparam equal_311_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i12542_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(GND_net), .I3(GND_net), .O(n28387));   // verilog/coms.v(130[12] 305[6])
    defparam i12542_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 select_787_Select_122_i2_4_lut (.I0(\data_out_frame[15] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5485));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_122_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1550 (.I0(\data_out_frame[10] [7]), .I1(n25915), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5637));
    defparam i1_2_lut_adj_1550.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1551 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[11] [2]), .I3(n6_adj_5637), .O(n56019));
    defparam i4_4_lut_adj_1551.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1552 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n55145), .I3(\FRAME_MATCHER.i[0] ), .O(n55149));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1552.LUT_INIT = 16'hfdff;
    SB_LUT4 select_787_Select_121_i2_4_lut (.I0(\data_out_frame[15] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5484));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_121_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_3_lut_4_lut_adj_1553 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(n55498), .I3(LED_c), .O(n26960));   // verilog/coms.v(148[4] 304[11])
    defparam i1_3_lut_4_lut_adj_1553.LUT_INIT = 16'hfe00;
    SB_LUT4 i2_2_lut_adj_1554 (.I0(n37_adj_5611), .I1(n56019), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_5638));
    defparam i2_2_lut_adj_1554.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_1555 (.I0(n50298), .I1(n7_adj_5638), .I2(\data_out_frame[15] [5]), 
            .I3(n8_adj_5596), .O(n51219));
    defparam i2_4_lut_adj_1555.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.i_31__N_2511 ), 
            .I2(GND_net), .I3(GND_net), .O(n55427));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i3_4_lut_adj_1556 (.I0(n50183), .I1(n1699), .I2(\data_out_frame[14] [1]), 
            .I3(n26123), .O(n58239));
    defparam i3_4_lut_adj_1556.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_120_i2_4_lut (.I0(\data_out_frame[15] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(pwm_setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5483));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_120_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1557 (.I0(\FRAME_MATCHER.i_31__N_2508 ), .I1(\FRAME_MATCHER.i_31__N_2512 ), 
            .I2(\FRAME_MATCHER.i_31__N_2514 ), .I3(GND_net), .O(n3484));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_3_lut_adj_1557.LUT_INIT = 16'hfefe;
    SB_LUT4 i16_4_lut_adj_1558 (.I0(n56056), .I1(n50249), .I2(n1720), 
            .I3(n26368), .O(n40_adj_5639));
    defparam i16_4_lut_adj_1558.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1559 (.I0(n56258), .I1(\data_out_frame[14] [6]), 
            .I2(n50331), .I3(\data_out_frame[11] [7]), .O(n38_adj_5640));
    defparam i14_4_lut_adj_1559.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1560 (.I0(\data_out_frame[11] [6]), .I1(n56186), 
            .I2(\data_out_frame[11] [5]), .I3(n56192), .O(n39_adj_5641));
    defparam i15_4_lut_adj_1560.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1561 (.I0(n56044), .I1(n56195), .I2(n58239), 
            .I3(n26479), .O(n37_adj_5642));
    defparam i13_4_lut_adj_1561.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49741 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[6] [3]), .I2(\data_out_frame[7] [3]), .I3(byte_transmit_counter[1]), 
            .O(n66813));
    defparam byte_transmit_counter_0__bdd_4_lut_49741.LUT_INIT = 16'he4aa;
    SB_LUT4 i18_4_lut_adj_1562 (.I0(\data_out_frame[8][3] ), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[10] [6]), .I3(\data_out_frame[11] [1]), 
            .O(n42_adj_5643));
    defparam i18_4_lut_adj_1562.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_119_i2_4_lut (.I0(\data_out_frame[14] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5482));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_119_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n66813_bdd_4_lut (.I0(n66813), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[4] [3]), .I3(byte_transmit_counter[1]), 
            .O(n60040));
    defparam n66813_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i22_4_lut_adj_1563 (.I0(n37_adj_5642), .I1(n39_adj_5641), .I2(n38_adj_5640), 
            .I3(n40_adj_5639), .O(n46));
    defparam i22_4_lut_adj_1563.LUT_INIT = 16'h6996;
    SB_LUT4 equal_305_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_adj_4));   // verilog/coms.v(157[7:23])
    defparam equal_305_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i17_4_lut_adj_1564 (.I0(\data_out_frame[10] [2]), .I1(n55781), 
            .I2(\data_out_frame[7] [6]), .I3(n55873), .O(n41_adj_5644));
    defparam i17_4_lut_adj_1564.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1565 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[14] [6]), 
            .I2(setpoint[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5481));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1565.LUT_INIT = 16'ha088;
    SB_LUT4 i23_3_lut (.I0(n41_adj_5644), .I1(n46), .I2(n42_adj_5643), 
            .I3(GND_net), .O(n58240));
    defparam i23_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1566 (.I0(n1835), .I1(n55717), .I2(n58240), .I3(n55678), 
            .O(n12_adj_5645));
    defparam i5_4_lut_adj_1566.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1567 (.I0(n26479), .I1(n12_adj_5645), .I2(n55727), 
            .I3(n26368), .O(n58122));
    defparam i6_4_lut_adj_1567.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1568 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[6] [0]), .I3(GND_net), .O(n55630));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1568.LUT_INIT = 16'h9696;
    SB_LUT4 equal_304_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i[0] ), .I3(GND_net), .O(n8_adj_5430));   // verilog/coms.v(157[7:23])
    defparam equal_304_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_adj_1569 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n55565));
    defparam i1_2_lut_adj_1569.LUT_INIT = 16'h6666;
    SB_LUT4 i12539_2_lut_2_lut (.I0(reset), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n28384));   // verilog/coms.v(130[12] 305[6])
    defparam i12539_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_3_lut_adj_1570 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[10] [2]), 
            .I2(\data_out_frame[6] [0]), .I3(GND_net), .O(n55995));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1570.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1571 (.I0(\data_out_frame[12] [3]), .I1(n55995), 
            .I2(n55575), .I3(\data_out_frame[7] [7]), .O(n10_adj_5646));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1571.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1572 (.I0(n55565), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[8][2] ), .I3(n55630), .O(n10_adj_5647));   // verilog/coms.v(88[17:70])
    defparam i4_4_lut_adj_1572.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1573 (.I0(\data_out_frame[5] [4]), .I1(n10_adj_5647), 
            .I2(\data_out_frame[4] [0]), .I3(GND_net), .O(n1516));   // verilog/coms.v(88[17:70])
    defparam i5_3_lut_adj_1573.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1574 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[7] [4]), .I3(GND_net), .O(n55554));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1574.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1575 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n25820));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1575.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1576 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n56001));
    defparam i1_2_lut_adj_1576.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1577 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[14] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n56192));
    defparam i1_2_lut_adj_1577.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1578 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n55662));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_adj_1578.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1579 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n56053));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_adj_1579.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1580 (.I0(\data_out_frame[9] [5]), .I1(n56053), 
            .I2(n55662), .I3(\data_out_frame[5] [3]), .O(n25642));   // verilog/coms.v(76[16:34])
    defparam i3_4_lut_adj_1580.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1581 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n55575));   // verilog/coms.v(88[17:70])
    defparam i1_2_lut_adj_1581.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1582 (.I0(\data_out_frame[10] [0]), .I1(n25642), 
            .I2(GND_net), .I3(GND_net), .O(n26092));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_adj_1582.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1583 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n30_adj_5648));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_adj_1583.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1584 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n55998));
    defparam i1_2_lut_adj_1584.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_117_i2_4_lut (.I0(\data_out_frame[14] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5480));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_117_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1585 (.I0(\data_out_frame[12] [1]), .I1(n55998), 
            .I2(n56189), .I3(n30_adj_5648), .O(n50391));
    defparam i1_4_lut_adj_1585.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1586 (.I0(n56192), .I1(n56001), .I2(n25820), 
            .I3(n4_adj_5649), .O(n51140));
    defparam i2_4_lut_adj_1586.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1587 (.I0(\data_out_frame[14] [5]), .I1(n1516), 
            .I2(n55805), .I3(\data_out_frame[12] [4]), .O(n26479));
    defparam i1_4_lut_adj_1587.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1588 (.I0(n55884), .I1(n26479), .I2(n51140), 
            .I3(\data_out_frame[16] [6]), .O(n10));
    defparam i4_4_lut_adj_1588.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1589 (.I0(\data_out_frame[16] [4]), .I1(n10), .I2(n25494), 
            .I3(GND_net), .O(n50372));
    defparam i5_3_lut_adj_1589.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1590 (.I0(n58122), .I1(n51219), .I2(\data_out_frame[16] [0]), 
            .I3(GND_net), .O(n55884));
    defparam i2_3_lut_adj_1590.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1591 (.I0(n47470), .I1(control_mode[1]), 
            .I2(control_mode[0]), .I3(GND_net), .O(n15));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_adj_1591.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_adj_1592 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n25656));
    defparam i1_2_lut_adj_1592.LUT_INIT = 16'h6666;
    SB_LUT4 i22452_3_lut_4_lut (.I0(n47470), .I1(control_mode[1]), .I2(control_update), 
            .I3(control_mode[0]), .O(n27260));   // verilog/coms.v(130[12] 305[6])
    defparam i22452_3_lut_4_lut.LUT_INIT = 16'hb0f0;
    SB_LUT4 i1_2_lut_3_lut_adj_1593 (.I0(control_mode[1]), .I1(n47470), 
            .I2(control_mode[0]), .I3(GND_net), .O(n15_adj_5));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_adj_1593.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1594 (.I0(control_mode[1]), .I1(n47470), 
            .I2(control_mode[0]), .I3(GND_net), .O(n15_adj_6));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_3_lut_adj_1594.LUT_INIT = 16'hefef;
    SB_LUT4 i4_4_lut_adj_1595 (.I0(n7_adj_5594), .I1(\data_out_frame[19] [1]), 
            .I2(n55884), .I3(n55766), .O(n55590));   // verilog/coms.v(88[17:28])
    defparam i4_4_lut_adj_1595.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1596 (.I0(\data_in_frame[16] [4]), .I1(n50260), 
            .I2(n25941), .I3(\data_in_frame[16] [5]), .O(n50620));
    defparam i1_2_lut_3_lut_4_lut_adj_1596.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1597 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5654));
    defparam i1_2_lut_adj_1597.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1598 (.I0(n50190), .I1(\data_out_frame[16] [7]), 
            .I2(n26479), .I3(n6_adj_5654), .O(n56094));
    defparam i4_4_lut_adj_1598.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1599 (.I0(\data_out_frame[21] [4]), .I1(n56228), 
            .I2(n56088), .I3(\data_out_frame[19] [3]), .O(n50266));   // verilog/coms.v(79[16:43])
    defparam i3_4_lut_adj_1599.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1600 (.I0(\data_out_frame[21] [3]), .I1(n56094), 
            .I2(n56024), .I3(\data_out_frame[16] [1]), .O(n51210));
    defparam i3_4_lut_adj_1600.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_116_i2_4_lut (.I0(\data_out_frame[14] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5479));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_116_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_115_i2_4_lut (.I0(\data_out_frame[14] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5478));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_115_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1601 (.I0(n57829), .I1(n56177), .I2(GND_net), 
            .I3(GND_net), .O(n55935));
    defparam i1_2_lut_adj_1601.LUT_INIT = 16'h9999;
    SB_LUT4 select_787_Select_114_i2_4_lut (.I0(\data_out_frame[14] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5477));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_114_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i3_3_lut_adj_1602 (.I0(\data_out_frame[23] [6]), .I1(n51378), 
            .I2(n56129), .I3(GND_net), .O(n8_adj_5655));
    defparam i3_3_lut_adj_1602.LUT_INIT = 16'h6969;
    SB_LUT4 select_787_Select_208_i3_4_lut (.I0(\data_out_frame[23] [4]), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n8_adj_5655), .I3(n55878), 
            .O(n3));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_208_i3_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i2_3_lut_4_lut_adj_1603 (.I0(\FRAME_MATCHER.i[0] ), .I1(n38266), 
            .I2(n3484), .I3(n37097), .O(n38695));
    defparam i2_3_lut_4_lut_adj_1603.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_3_lut_adj_1604 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [2]), 
            .I2(n55738), .I3(GND_net), .O(n56088));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1604.LUT_INIT = 16'h9696;
    SB_LUT4 i4_2_lut_3_lut (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [2]), 
            .I2(\data_out_frame[16] [3]), .I3(GND_net), .O(n15_adj_5595));   // verilog/coms.v(79[16:43])
    defparam i4_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_207_i2_4_lut (.I0(\data_out_frame[25] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5393));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_207_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1605 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [2]), 
            .I2(n55590), .I3(GND_net), .O(n56024));   // verilog/coms.v(79[16:43])
    defparam i1_2_lut_3_lut_adj_1605.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1606 (.I0(\data_out_frame[12] [2]), .I1(n55554), 
            .I2(\data_out_frame[5] [6]), .I3(\data_out_frame[14] [4]), .O(n56186));
    defparam i1_2_lut_4_lut_adj_1606.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1607 (.I0(\data_out_frame[12] [2]), .I1(n55554), 
            .I2(\data_out_frame[5] [6]), .I3(n50391), .O(n4_adj_5649));
    defparam i1_2_lut_4_lut_adj_1607.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut_3_lut_adj_1608 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[9] [6]), .I3(GND_net), .O(n18_adj_5622));
    defparam i4_2_lut_3_lut_adj_1608.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1609 (.I0(control_mode[5]), .I1(control_mode[4]), 
            .I2(GND_net), .I3(GND_net), .O(n59336));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_adj_1609.LUT_INIT = 16'heeee;
    SB_LUT4 select_787_Select_113_i2_4_lut (.I0(\data_out_frame[14] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5476));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_113_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i39367_3_lut_4_lut (.I0(\FRAME_MATCHER.i[0] ), .I1(n38266), 
            .I2(n55515), .I3(reset), .O(n27906));
    defparam i39367_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_4_lut_adj_1610 (.I0(control_mode[7]), .I1(n33_adj_5633), 
            .I2(n59336), .I3(control_mode[6]), .O(n47470));   // verilog/coms.v(130[12] 305[6])
    defparam i1_4_lut_adj_1610.LUT_INIT = 16'hfffe;
    SB_LUT4 select_787_Select_112_i2_4_lut (.I0(\data_out_frame[14] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5475));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_112_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_111_i2_4_lut (.I0(\data_out_frame[13] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5474));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_111_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_4_lut_adj_1611 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[10] [1]), .I3(n10_adj_5646), .O(n55805));
    defparam i5_3_lut_4_lut_adj_1611.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_110_i2_4_lut (.I0(\data_out_frame[13] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5473));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_110_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_109_i2_4_lut (.I0(\data_out_frame[13] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5472));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_109_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_206_i2_4_lut (.I0(\data_out_frame[25] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5391));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_206_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_4_lut_adj_1612 (.I0(\data_out_frame[25] [2]), .I1(\data_out_frame[25] [3]), 
            .I2(n10_adj_5575), .I3(\data_out_frame[25] [1]), .O(n51156));
    defparam i5_3_lut_4_lut_adj_1612.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_53_i2_4_lut (.I0(\data_out_frame[6] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[21] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5389));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_53_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_108_i2_4_lut (.I0(\data_out_frame[13] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5471));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_108_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_205_i2_4_lut (.I0(\data_out_frame[25] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5388));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_205_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_204_i2_4_lut (.I0(\data_out_frame[25] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5387));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_204_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_107_i2_4_lut (.I0(\data_out_frame[13] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5470));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_107_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_203_i2_4_lut (.I0(\data_out_frame[25] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5386));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_203_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_106_i2_4_lut (.I0(\data_out_frame[13] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5469));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_106_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1613 (.I0(n1959), .I1(n4452), .I2(n1962), 
            .I3(n1965), .O(n57378));   // verilog/coms.v(145[4] 147[7])
    defparam i2_3_lut_4_lut_adj_1613.LUT_INIT = 16'h2000;
    SB_LUT4 select_787_Select_202_i2_4_lut (.I0(\data_out_frame[25] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5385));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_202_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_4_lut_4_lut (.I0(n1959), .I1(n4452), .I2(n59705), .I3(\FRAME_MATCHER.i_31__N_2514 ), 
            .O(n57595));   // verilog/coms.v(145[4] 147[7])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'ha2a0;
    SB_LUT4 select_787_Select_105_i2_4_lut (.I0(\data_out_frame[13] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5468));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_105_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_201_i2_4_lut (.I0(\data_out_frame[25] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5384));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_201_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13620_3_lut_4_lut (.I0(n27862), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[19]_c [7]), .O(n29465));
    defparam i13620_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_200_i2_4_lut (.I0(\data_out_frame[25] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5383));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_200_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1614 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[18] [6]), 
            .I2(displacement[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5290));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1614.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_199_i2_4_lut (.I0(\data_out_frame[24] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5382));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_199_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1615 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[24] [6]), 
            .I2(neopxl_color[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5381));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1615.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_104_i2_4_lut (.I0(\data_out_frame[13] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5467));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_104_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13617_3_lut_4_lut (.I0(n27862), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[19]_c [6]), .O(n29462));
    defparam i13617_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13614_3_lut_4_lut (.I0(n27862), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[19]_c [5]), .O(n29459));
    defparam i13614_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1616 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[18] [3]), 
            .I2(n49936), .I3(n51146), .O(n14_adj_5572));
    defparam i5_3_lut_4_lut_adj_1616.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_49587 (.I0(byte_transmit_counter[1]), 
            .I1(n60099), .I2(n60100), .I3(byte_transmit_counter[2]), .O(n66645));
    defparam byte_transmit_counter_1__bdd_4_lut_49587.LUT_INIT = 16'he4aa;
    SB_LUT4 select_787_Select_197_i2_4_lut (.I0(\data_out_frame[24] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5380));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_197_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_103_i2_4_lut (.I0(\data_out_frame[12] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5466));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_103_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_196_i2_4_lut (.I0(\data_out_frame[24] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5379));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_196_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i11_3_lut_4_lut (.I0(n27862), .I1(reset), .I2(\data_in_frame[19]_c [4]), 
            .I3(rx_data[4]), .O(n54599));
    defparam i11_3_lut_4_lut.LUT_INIT = 16'hf1e0;
    SB_LUT4 select_787_Select_195_i2_4_lut (.I0(\data_out_frame[24] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5378));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_195_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_102_i2_4_lut (.I0(\data_out_frame[12] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5465));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_102_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_149_i2_4_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5289));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_149_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13608_3_lut_4_lut (.I0(n27862), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[19]_c [3]), .O(n29453));
    defparam i13608_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_4_lut (.I0(n27862), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n54635));
    defparam i11_4_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_194_i2_4_lut (.I0(\data_out_frame[24] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5377));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_194_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_101_i2_4_lut (.I0(\data_out_frame[12] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(setpoint[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5464));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_101_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13601_3_lut_4_lut (.I0(n27862), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n29446));
    defparam i13601_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_148_i2_4_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5288));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_148_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_193_i2_4_lut (.I0(\data_out_frame[24] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5376));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_193_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n66645_bdd_4_lut (.I0(n66645), .I1(n60097), .I2(n60096), .I3(byte_transmit_counter[2]), 
            .O(n14_adj_5656));
    defparam n66645_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13598_3_lut_4_lut (.I0(n27862), .I1(reset), .I2(rx_data[0]), 
            .I3(\data_in_frame[19][0] ), .O(n29443));
    defparam i13598_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_52_i2_4_lut (.I0(\data_out_frame[6] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[20] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5375));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_52_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1617 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[12] [4]), 
            .I2(setpoint[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5463));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1617.LUT_INIT = 16'ha088;
    SB_LUT4 i2_3_lut_4_lut_adj_1618 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [6]), 
            .I2(\data_out_frame[7] [2]), .I3(\data_out_frame[5] [1]), .O(n25661));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_4_lut_adj_1618.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_99_i2_4_lut (.I0(\data_out_frame[12] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5462));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_99_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_3_lut_4_lut_adj_1619 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [6]), 
            .I2(\data_out_frame[4] [7]), .I3(n10_adj_5636), .O(n50298));   // verilog/coms.v(88[17:70])
    defparam i5_3_lut_4_lut_adj_1619.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_51_i2_4_lut (.I0(\data_out_frame[6] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[19] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5374));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_51_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1620 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[12] [2]), 
            .I2(setpoint[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5461));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1620.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_50_i2_4_lut (.I0(\data_out_frame[6] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[18] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5373));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_50_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1621 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[4] [6]), 
            .I2(\data_out_frame[7] [0]), .I3(n1168), .O(n25915));   // verilog/coms.v(88[17:70])
    defparam i2_3_lut_4_lut_adj_1621.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1622 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[7] [3]), .I3(GND_net), .O(n55742));   // verilog/coms.v(76[16:34])
    defparam i1_2_lut_3_lut_adj_1622.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1623 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(n55543), .I3(n1191), .O(n1168));   // verilog/coms.v(76[16:34])
    defparam i2_3_lut_4_lut_adj_1623.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_97_i2_4_lut (.I0(\data_out_frame[12] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5460));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_97_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1624 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[4] [2]), .I3(\data_out_frame[8][5] ), .O(n56030));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_4_lut_adj_1624.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1625 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[4] [2]), .I3(\data_out_frame[8][6] ), .O(n37_adj_5611));   // verilog/coms.v(100[12:26])
    defparam i1_2_lut_4_lut_adj_1625.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1626 (.I0(\data_out_frame[4] [0]), .I1(n55873), 
            .I2(n10_adj_5625), .I3(n26378), .O(n55579));   // verilog/coms.v(77[16:43])
    defparam i5_3_lut_4_lut_adj_1626.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_96_i2_4_lut (.I0(\data_out_frame[12] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(setpoint[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5459));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_96_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_49_i2_4_lut (.I0(\data_out_frame[6] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[17] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5372));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_49_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14015_3_lut_4_lut (.I0(n8_adj_5430), .I1(n55507), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n29860));
    defparam i14015_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1627 (.I0(\data_out_frame[19] [0]), .I1(n25687), 
            .I2(n50591), .I3(\data_out_frame[21] [2]), .O(n51378));
    defparam i1_2_lut_4_lut_adj_1627.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_192_i2_4_lut (.I0(\data_out_frame[24] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5371));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_192_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i5_2_lut_4_lut (.I0(\data_out_frame[19] [0]), .I1(n25687), .I2(n50591), 
            .I3(n51265), .O(n15_adj_5570));
    defparam i5_2_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i13752_3_lut_4_lut (.I0(n8_adj_4), .I1(n55507), .I2(rx_data[0]), 
            .I3(\data_in_frame[0]_c [0]), .O(n29597));
    defparam i13752_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_49562 (.I0(byte_transmit_counter[1]), 
            .I1(n60129), .I2(n60130), .I3(byte_transmit_counter[2]), .O(n66639));
    defparam byte_transmit_counter_1__bdd_4_lut_49562.LUT_INIT = 16'he4aa;
    SB_LUT4 select_787_Select_95_i2_4_lut (.I0(\data_out_frame[11] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5458));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_95_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13982_3_lut_4_lut (.I0(n8_adj_4), .I1(n55507), .I2(rx_data[1]), 
            .I3(\data_in_frame[0]_c [1]), .O(n29827));
    defparam i13982_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13985_3_lut_4_lut (.I0(n8_adj_4), .I1(n55507), .I2(rx_data[2]), 
            .I3(\data_in_frame[0]_c [2]), .O(n29830));
    defparam i13985_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_94_i2_4_lut (.I0(\data_out_frame[11] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5457));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_94_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_48_i2_4_lut (.I0(\data_out_frame[6] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\encoder0_position_scaled[16] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5370));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_48_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_191_i2_4_lut (.I0(\data_out_frame[23] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5369));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_191_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13988_3_lut_4_lut (.I0(n8_adj_4), .I1(n55507), .I2(rx_data[3]), 
            .I3(\data_in_frame[0]_c [3]), .O(n29833));
    defparam i13988_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13991_3_lut_4_lut (.I0(n8_adj_4), .I1(n55507), .I2(rx_data[4]), 
            .I3(\data_in_frame[0][4] ), .O(n29836));
    defparam i13991_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13994_3_lut_4_lut (.I0(n8_adj_4), .I1(n55507), .I2(rx_data[5]), 
            .I3(\data_in_frame[0]_c [5]), .O(n29839));
    defparam i13994_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_93_i2_4_lut (.I0(\data_out_frame[11] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5456));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_93_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13997_3_lut_4_lut (.I0(n8_adj_4), .I1(n55507), .I2(rx_data[6]), 
            .I3(\data_in_frame[0]_c [6]), .O(n29842));
    defparam i13997_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14000_3_lut_4_lut (.I0(n8_adj_4), .I1(n55507), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n29845));
    defparam i14000_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_190_i2_4_lut (.I0(\data_out_frame[23] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5368));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_190_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1628 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[5] [7]), 
            .I2(control_mode[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5367));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1628.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_189_i2_4_lut (.I0(\data_out_frame[23] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5366));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_189_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n66639_bdd_4_lut (.I0(n66639), .I1(n60091), .I2(n60090), .I3(byte_transmit_counter[2]), 
            .O(n66642));
    defparam n66639_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_787_Select_46_i2_4_lut (.I0(\data_out_frame[5] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5365));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_46_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_188_i2_4_lut (.I0(\data_out_frame[23] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5364));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_188_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_187_i2_4_lut (.I0(\data_out_frame[23] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5363));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_187_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_186_i2_4_lut (.I0(\data_out_frame[23] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5362));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_186_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_185_i2_4_lut (.I0(\data_out_frame[23] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(neopxl_color[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5361));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_185_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_45_i2_4_lut (.I0(\data_out_frame[5] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5360));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_45_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_44_i2_4_lut (.I0(\data_out_frame[5] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5359));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_44_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1629 (.I0(n50388), .I1(n57849), .I2(\data_out_frame[20] [0]), 
            .I3(\data_out_frame[22] [7]), .O(n56231));
    defparam i2_3_lut_4_lut_adj_1629.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1630 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[5] [3]), 
            .I2(control_mode[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5358));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1630.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_42_i2_4_lut (.I0(\data_out_frame[5] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5357));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_42_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_3_lut_4_lut_adj_1631 (.I0(\data_out_frame[15] [4]), .I1(n1720), 
            .I2(n55778), .I3(\data_out_frame[17] [5]), .O(n50229));
    defparam i2_3_lut_4_lut_adj_1631.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1632 (.I0(\data_out_frame[15] [4]), .I1(n1720), 
            .I2(\data_out_frame[17] [6]), .I3(n56225), .O(n58113));
    defparam i2_3_lut_4_lut_adj_1632.LUT_INIT = 16'h6996;
    SB_LUT4 i19054_3_lut (.I0(n27926), .I1(rx_data[6]), .I2(\data_in_frame[17]_c [6]), 
            .I3(GND_net), .O(n29414));   // verilog/coms.v(94[13:20])
    defparam i19054_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n4_adj_5562), .I2(n5_adj_5561), .I3(byte_transmit_counter[2]), 
            .O(n66807));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n66807_bdd_4_lut (.I0(n66807), .I1(n62988), .I2(n62987), .I3(byte_transmit_counter[2]), 
            .O(n60044));
    defparam n66807_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1633 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[18] [2]), 
            .I2(n51330), .I3(GND_net), .O(n55992));
    defparam i1_2_lut_3_lut_adj_1633.LUT_INIT = 16'h6969;
    SB_LUT4 i13_3_lut_4_lut (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[18] [2]), 
            .I2(\data_out_frame[19] [3]), .I3(\data_out_frame[17] [6]), 
            .O(n38));
    defparam i13_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_49557 (.I0(byte_transmit_counter[1]), 
            .I1(n60084), .I2(n60085), .I3(byte_transmit_counter[2]), .O(n66633));
    defparam byte_transmit_counter_1__bdd_4_lut_49557.LUT_INIT = 16'he4aa;
    SB_LUT4 n66633_bdd_4_lut (.I0(n66633), .I1(n60067), .I2(n60066), .I3(byte_transmit_counter[2]), 
            .O(n66636));
    defparam n66633_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(n66588), .I2(n66576), .I3(byte_transmit_counter_c[3]), 
            .O(n66627));
    defparam byte_transmit_counter_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n66627_bdd_4_lut (.I0(n66627), .I1(n60040), .I2(n60039), .I3(byte_transmit_counter_c[3]), 
            .O(n66630));
    defparam n66627_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49567 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [5]), .I2(\data_out_frame[23] [5]), 
            .I3(byte_transmit_counter[1]), .O(n66621));
    defparam byte_transmit_counter_0__bdd_4_lut_49567.LUT_INIT = 16'he4aa;
    SB_LUT4 n66621_bdd_4_lut (.I0(n66621), .I1(\data_out_frame[21] [5]), 
            .I2(\data_out_frame[20] [5]), .I3(byte_transmit_counter[1]), 
            .O(n66624));
    defparam n66621_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1634 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[5] [1]), 
            .I2(control_mode[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5356));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1634.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_40_i2_4_lut (.I0(\data_out_frame[5] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(control_mode[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5355));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_40_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1635 (.I0(n50183), .I1(n4), .I2(n50685), 
            .I3(GND_net), .O(n55989));
    defparam i1_2_lut_3_lut_adj_1635.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1636 (.I0(n50183), .I1(n4), .I2(n25385), 
            .I3(n49936), .O(n57257));
    defparam i2_3_lut_4_lut_adj_1636.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1637 (.I0(\data_out_frame[20] [4]), .I1(n55793), 
            .I2(\data_out_frame[23] [1]), .I3(GND_net), .O(n56201));
    defparam i1_2_lut_3_lut_adj_1637.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1638 (.I0(\data_out_frame[20] [4]), .I1(n55793), 
            .I2(\data_out_frame[20] [5]), .I3(n55861), .O(n50270));
    defparam i2_3_lut_4_lut_adj_1638.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1639 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [1]), 
            .I2(n50410), .I3(n58154), .O(n23288));
    defparam i2_3_lut_4_lut_adj_1639.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1640 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [1]), 
            .I2(\data_out_frame[20] [2]), .I3(GND_net), .O(n55793));
    defparam i1_2_lut_3_lut_adj_1640.LUT_INIT = 16'h9696;
    SB_LUT4 i49205_2_lut_3_lut (.I0(\data_in_frame[0]_c [3]), .I1(\data_in_frame[0]_c [2]), 
            .I2(\data_in_frame[2]_c [4]), .I3(GND_net), .O(n66267));   // verilog/coms.v(99[12:25])
    defparam i49205_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_39_i2_4_lut (.I0(\data_out_frame[4] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5354));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_39_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_38_i2_4_lut (.I0(\data_out_frame[4] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5353));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_38_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1641 (.I0(Kp_23__N_758), .I1(\data_in_frame[2]_c [4]), 
            .I2(n25908), .I3(\data_in_frame[4] [5]), .O(n50417));
    defparam i1_2_lut_4_lut_adj_1641.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_4_lut_adj_1642 (.I0(\data_out_frame[20] [3]), .I1(n58154), 
            .I2(n51376), .I3(\data_out_frame[22] [5]), .O(n50377));
    defparam i1_3_lut_4_lut_adj_1642.LUT_INIT = 16'h9669;
    SB_LUT4 select_787_Select_37_i2_4_lut (.I0(\data_out_frame[4] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5352));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_37_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_92_i2_4_lut (.I0(\data_out_frame[11] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5455));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_92_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_36_i2_4_lut (.I0(\data_out_frame[4] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5351));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_36_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1643 (.I0(\data_out_frame[20] [3]), .I1(n58154), 
            .I2(n51302), .I3(\data_out_frame[20] [2]), .O(n51282));
    defparam i1_2_lut_3_lut_4_lut_adj_1643.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1644 (.I0(n51256), .I1(n55757), .I2(n56174), 
            .I3(n50317), .O(n55975));
    defparam i2_3_lut_4_lut_adj_1644.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1645 (.I0(\data_out_frame[20] [2]), .I1(n51302), 
            .I2(\data_out_frame[22] [3]), .I3(n55572), .O(n24672));
    defparam i2_3_lut_4_lut_adj_1645.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1646 (.I0(Kp_23__N_1080), .I1(n55652), .I2(\data_in_frame[8] [7]), 
            .I3(n51230), .O(n50317));
    defparam i2_3_lut_4_lut_adj_1646.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1647 (.I0(\data_in_frame[5] [2]), .I1(n55665), 
            .I2(n51230), .I3(GND_net), .O(n56153));
    defparam i1_2_lut_3_lut_adj_1647.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1648 (.I0(\data_in_frame[9] [2]), .I1(n57296), 
            .I2(n26031), .I3(GND_net), .O(n55721));
    defparam i1_2_lut_3_lut_adj_1648.LUT_INIT = 16'h6969;
    SB_LUT4 select_787_Select_91_i2_4_lut (.I0(\data_out_frame[11] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5454));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_91_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i2_2_lut_3_lut_adj_1649 (.I0(\data_in_frame[5] [2]), .I1(n55665), 
            .I2(\data_in_frame[9] [3]), .I3(GND_net), .O(n7_adj_5529));
    defparam i2_2_lut_3_lut_adj_1649.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1650 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n55145), .O(n55151));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1650.LUT_INIT = 16'hffef;
    SB_LUT4 i1_4_lut_adj_1651 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[11] [2]), 
            .I2(encoder1_position_scaled[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5453));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1651.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_35_i2_4_lut (.I0(\data_out_frame[4] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5350));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_35_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1652 (.I0(\data_in_frame[11] [3]), .I1(\data_in_frame[9] [1]), 
            .I2(\data_in_frame[9] [2]), .I3(GND_net), .O(n56237));
    defparam i1_2_lut_3_lut_adj_1652.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1653 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[4] [2]), 
            .I2(ID[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5349));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1653.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_3_lut_adj_1654 (.I0(\data_in_frame[10] [4]), .I1(n55760), 
            .I2(\data_in_frame[12] [5]), .I3(GND_net), .O(n55684));
    defparam i1_2_lut_3_lut_adj_1654.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1655 (.I0(n51319), .I1(\data_in_frame[10] [0]), 
            .I2(\data_in_frame[12] [3]), .I3(GND_net), .O(n55938));
    defparam i1_2_lut_3_lut_adj_1655.LUT_INIT = 16'h6969;
    SB_LUT4 i1_4_lut_adj_1656 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[23] [0]), 
            .I2(neopxl_color[16]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5348));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1656.LUT_INIT = 16'ha088;
    SB_LUT4 i1_2_lut_4_lut_adj_1657 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n50744), .I3(n25572), .O(n51319));
    defparam i1_2_lut_4_lut_adj_1657.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1658 (.I0(\data_in_frame[15] [7]), .I1(n55684), 
            .I2(\data_in_frame[13] [0]), .I3(n26055), .O(n56047));
    defparam i1_2_lut_4_lut_adj_1658.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1659 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(n55745), .I3(n51228), .O(n51247));
    defparam i2_3_lut_4_lut_adj_1659.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1660 (.I0(n58201), .I1(\data_in_frame[12] [4]), 
            .I2(n25607), .I3(\data_in_frame[12] [5]), .O(n57943));
    defparam i2_3_lut_4_lut_adj_1660.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1661 (.I0(\data_in_frame[15] [0]), .I1(\data_in_frame[12] [4]), 
            .I2(n26257), .I3(GND_net), .O(n55772));
    defparam i1_2_lut_3_lut_adj_1661.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_147_i2_4_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5287));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_147_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_89_i2_4_lut (.I0(\data_out_frame[11] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5452));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_89_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_146_i2_4_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5286));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_146_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1662 (.I0(\data_in_frame[20] [7]), .I1(\data_in_frame[19][0] ), 
            .I2(n50310), .I3(n55775), .O(n56168));
    defparam i1_2_lut_4_lut_adj_1662.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1663 (.I0(\data_in_frame[16] [3]), .I1(n50272), 
            .I2(n50260), .I3(GND_net), .O(n55819));
    defparam i1_2_lut_3_lut_adj_1663.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1664 (.I0(\data_in_frame[15] [5]), .I1(n51168), 
            .I2(n51359), .I3(\data_in_frame[17]_c [6]), .O(n56132));
    defparam i1_2_lut_4_lut_adj_1664.LUT_INIT = 16'h9669;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(156[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_787_Select_183_i2_4_lut (.I0(\data_out_frame[22] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[7] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5343));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_183_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1665 (.I0(\data_in_frame[13] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(n50317), .I3(n51228), .O(n51168));
    defparam i1_2_lut_4_lut_adj_1665.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1666 (.I0(\FRAME_MATCHER.i[5] ), .I1(n73), .I2(GND_net), 
            .I3(GND_net), .O(n37097));   // verilog/coms.v(156[9:50])
    defparam i1_2_lut_adj_1666.LUT_INIT = 16'h4444;
    SB_LUT4 i3_3_lut_4_lut_adj_1667 (.I0(\data_in_frame[10] [7]), .I1(Kp_23__N_974), 
            .I2(\data_in_frame[8] [6]), .I3(\data_in_frame[11] [0]), .O(n56117));   // verilog/coms.v(74[16:27])
    defparam i3_3_lut_4_lut_adj_1667.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_49696 (.I0(byte_transmit_counter[1]), 
            .I1(n11_adj_5559), .I2(n12_adj_5558), .I3(byte_transmit_counter[2]), 
            .O(n66801));
    defparam byte_transmit_counter_1__bdd_4_lut_49696.LUT_INIT = 16'he4aa;
    SB_LUT4 n66801_bdd_4_lut (.I0(n66801), .I1(n9_adj_5557), .I2(n62989), 
            .I3(byte_transmit_counter[2]), .O(n66804));
    defparam n66801_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1668 (.I0(\data_out_frame[20] [5]), .I1(n51376), 
            .I2(n55784), .I3(n26012), .O(n57163));
    defparam i2_3_lut_4_lut_adj_1668.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_3_lut_adj_1669 (.I0(\data_in_frame[12] [7]), .I1(n50317), 
            .I2(\data_in_frame[15] [2]), .I3(GND_net), .O(n10_adj_5516));
    defparam i2_2_lut_3_lut_adj_1669.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut_adj_1670 (.I0(\data_out_frame[20] [5]), .I1(n51376), 
            .I2(n55959), .I3(n55823), .O(n8_adj_5573));
    defparam i3_3_lut_4_lut_adj_1670.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_182_i2_4_lut (.I0(\data_out_frame[22] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[6] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5342));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_182_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_33_i2_4_lut (.I0(\data_out_frame[4] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5338));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_33_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13474_3_lut_4_lut (.I0(n8_adj_5577), .I1(n55145), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n29319));
    defparam i13474_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_4_lut_adj_1671 (.I0(\data_in_frame[13] [5]), .I1(n55917), 
            .I2(\data_in_frame[13] [4]), .I3(\data_in_frame[18] [0]), .O(n7_adj_5512));
    defparam i2_2_lut_4_lut_adj_1671.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1672 (.I0(\data_in_frame[15] [6]), .I1(n51228), 
            .I2(n55926), .I3(GND_net), .O(n55978));
    defparam i1_2_lut_3_lut_adj_1672.LUT_INIT = 16'h6969;
    SB_LUT4 i1_3_lut_4_lut_adj_1673 (.I0(\data_in_frame[10] [4]), .I1(n55760), 
            .I2(\data_in_frame[15] [1]), .I3(\data_in_frame[17][2] ), .O(n59538));
    defparam i1_3_lut_4_lut_adj_1673.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_32_i2_4_lut (.I0(\data_out_frame[4] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(ID[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), .O(n2_adj_5337));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_32_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13477_3_lut_4_lut (.I0(n8_adj_5577), .I1(n55145), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n29322));
    defparam i13477_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1674 (.I0(\data_in_frame[19]_c [3]), .I1(n56181), 
            .I2(n32987), .I3(\data_in_frame[21][4] ), .O(n50368));
    defparam i1_2_lut_4_lut_adj_1674.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1675 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(\data_in_frame[18] [3]), .I3(\data_in_frame[18] [0]), .O(n59542));
    defparam i1_2_lut_4_lut_adj_1675.LUT_INIT = 16'h6996;
    SB_LUT4 select_787_Select_88_i2_4_lut (.I0(\data_out_frame[11] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5451));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_88_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_49691 (.I0(byte_transmit_counter[1]), 
            .I1(n11_adj_5555), .I2(n12_adj_5554), .I3(byte_transmit_counter[2]), 
            .O(n66795));
    defparam byte_transmit_counter_1__bdd_4_lut_49691.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1676 (.I0(\data_in_frame[0]_c [6]), .I1(\data_in_frame[0]_c [5]), 
            .I2(GND_net), .I3(GND_net), .O(n55587));   // verilog/coms.v(80[16:27])
    defparam i1_2_lut_adj_1676.LUT_INIT = 16'h6666;
    SB_LUT4 i13480_3_lut_4_lut (.I0(n8_adj_5577), .I1(n55145), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n29325));
    defparam i13480_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n66795_bdd_4_lut (.I0(n66795), .I1(n9_adj_5553), .I2(n62990), 
            .I3(byte_transmit_counter[2]), .O(n66798));
    defparam n66795_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_787_Select_181_i2_4_lut (.I0(\data_out_frame[22] [5]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[5] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5336));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_181_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_adj_1677 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[0]_c [0]), 
            .I2(GND_net), .I3(GND_net), .O(n55560));   // verilog/coms.v(99[12:25])
    defparam i1_2_lut_adj_1677.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_180_i2_4_lut (.I0(\data_out_frame[22] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[4] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5335));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_180_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_179_i2_4_lut (.I0(\data_out_frame[22] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[3] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5334));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_179_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13483_3_lut_4_lut (.I0(n8_adj_5577), .I1(n55145), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n29328));
    defparam i13483_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1678 (.I0(\data_in_frame[16] [4]), .I1(n50260), 
            .I2(n55648), .I3(n55819), .O(n51243));
    defparam i1_2_lut_4_lut_adj_1678.LUT_INIT = 16'h6996;
    SB_LUT4 i13486_3_lut_4_lut (.I0(n8_adj_5577), .I1(n55145), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n29331));
    defparam i13486_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_178_i2_4_lut (.I0(\data_out_frame[22] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[2] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5333));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_178_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1679 (.I0(\data_in_frame[20] [6]), .I1(\data_in_frame[18] [3]), 
            .I2(n24707), .I3(GND_net), .O(n56246));
    defparam i1_2_lut_3_lut_adj_1679.LUT_INIT = 16'h9696;
    SB_LUT4 select_787_Select_177_i2_4_lut (.I0(\data_out_frame[22] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[1] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5332));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_177_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1680 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[22] [0]), 
            .I2(\current[0] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5331));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1680.LUT_INIT = 16'ha088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49701 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n66789));
    defparam byte_transmit_counter_0__bdd_4_lut_49701.LUT_INIT = 16'he4aa;
    SB_LUT4 select_787_Select_87_i2_4_lut (.I0(\data_out_frame[10] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5450));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_87_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_175_i2_4_lut (.I0(\data_out_frame[21] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5329));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_175_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1681 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n55145), .O(n55153));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1681.LUT_INIT = 16'hffdf;
    SB_LUT4 select_787_Select_174_i2_4_lut (.I0(\data_out_frame[21] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5328));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_174_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1682 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n55507), .O(n27902));   // verilog/coms.v(157[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1682.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_4_lut_adj_1683 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[21] [5]), 
            .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5327));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1683.LUT_INIT = 16'ha088;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n60110), .I3(n60108), .O(n7_adj_5635));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 select_787_Select_172_i2_4_lut (.I0(\data_out_frame[21] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[15] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5326));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_172_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n60062), .I3(n60060), .O(n7_adj_5627));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n60146), .I3(n60144), .O(n7_adj_5616));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n60056), .I3(n60054), .O(n7_adj_5613));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n60080), .I3(n60078), .O(n7_adj_5538));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n60077), .I3(n60075), .O(n7_adj_5585));   // verilog/coms.v(109[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 select_787_Select_216_i3_3_lut_4_lut (.I0(n57923), .I1(n51156), 
            .I2(\FRAME_MATCHER.state[3] ), .I3(n55896), .O(n3_adj_5402));
    defparam select_787_Select_216_i3_3_lut_4_lut.LUT_INIT = 16'h9060;
    SB_LUT4 select_787_Select_171_i2_4_lut (.I0(\data_out_frame[21] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[11] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5324));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_171_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_170_i2_4_lut (.I0(\data_out_frame[21] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[10] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5323));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_170_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n66789_bdd_4_lut (.I0(n66789), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n66792));
    defparam n66789_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49681 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n66783));
    defparam byte_transmit_counter_0__bdd_4_lut_49681.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_2_lut_3_lut_adj_1684 (.I0(n57923), .I1(n51156), .I2(\data_out_frame[24] [5]), 
            .I3(GND_net), .O(n6_adj_5576));
    defparam i2_2_lut_3_lut_adj_1684.LUT_INIT = 16'h6969;
    SB_LUT4 select_787_Select_169_i2_4_lut (.I0(\data_out_frame[21] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[9] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5322));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_169_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_3_lut_adj_1685 (.I0(n57678), .I1(\data_out_frame[23] [3]), 
            .I2(n57923), .I3(GND_net), .O(n55844));
    defparam i1_2_lut_3_lut_adj_1685.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut_adj_1686 (.I0(n57678), .I1(\data_out_frame[23] [3]), 
            .I2(n56243), .I3(n51210), .O(n8_adj_5435));
    defparam i3_3_lut_4_lut_adj_1686.LUT_INIT = 16'h9669;
    SB_LUT4 i13489_3_lut_4_lut (.I0(n8_adj_5577), .I1(n55145), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n29334));
    defparam i13489_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13492_3_lut_4_lut (.I0(n8_adj_5577), .I1(n55145), .I2(rx_data[6]), 
            .I3(\data_in_frame[14][6] ), .O(n29337));
    defparam i13492_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13495_3_lut_4_lut (.I0(n8_adj_5577), .I1(n55145), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n29340));
    defparam i13495_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n66783_bdd_4_lut (.I0(n66783), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n66786));
    defparam n66783_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1687 (.I0(\data_in_frame[2] [0]), .I1(Kp_23__N_748), 
            .I2(GND_net), .I3(GND_net), .O(n55748));   // verilog/coms.v(73[16:69])
    defparam i1_2_lut_adj_1687.LUT_INIT = 16'h6666;
    SB_LUT4 select_787_Select_168_i2_4_lut (.I0(\data_out_frame[21] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(\current[8] ), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5321));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_168_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1688 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[10] [6]), 
            .I2(encoder1_position_scaled[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n11));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1688.LUT_INIT = 16'ha088;
    SB_LUT4 i2_3_lut_adj_1689 (.I0(\data_in_frame[0]_c [1]), .I1(\data_in_frame[0]_c [0]), 
            .I2(\data_in_frame[2]_c [2]), .I3(GND_net), .O(n25933));   // verilog/coms.v(76[16:42])
    defparam i2_3_lut_adj_1689.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1690 (.I0(Kp_23__N_748), .I1(\data_in_frame[2]_c [7]), 
            .I2(\data_in_frame[2]_c [1]), .I3(n55587), .O(n23_c));
    defparam i6_4_lut_adj_1690.LUT_INIT = 16'h4812;
    SB_LUT4 i1_4_lut_adj_1691 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20] [7]), 
            .I2(displacement[7]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5320));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1691.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_166_i2_4_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[6]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5319));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_166_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_4_lut_adj_1692 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[20] [5]), 
            .I2(displacement[5]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5318));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1692.LUT_INIT = 16'ha088;
    SB_LUT4 select_787_Select_164_i2_4_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[4]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5316));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_164_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_163_i2_4_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[3]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5315));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_163_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i10_4_lut_adj_1693 (.I0(n66279), .I1(n66267), .I2(\data_in_frame[1] [5]), 
            .I3(n66277), .O(n27_adj_5657));
    defparam i10_4_lut_adj_1693.LUT_INIT = 16'h0010;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49676 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n66777));
    defparam byte_transmit_counter_0__bdd_4_lut_49676.LUT_INIT = 16'he4aa;
    SB_LUT4 i12_4_lut_adj_1694 (.I0(n23_c), .I1(n25908), .I2(Kp_23__N_748), 
            .I3(n55560), .O(n29_adj_5658));
    defparam i12_4_lut_adj_1694.LUT_INIT = 16'h0220;
    SB_LUT4 n66777_bdd_4_lut (.I0(n66777), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n66780));
    defparam n66777_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_787_Select_85_i2_4_lut (.I0(\data_out_frame[10] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[13]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5449));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_85_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i14_4_lut_adj_1695 (.I0(n27_adj_5657), .I1(\data_in_frame[1]_c [2]), 
            .I2(n22_adj_5528), .I3(\data_in_frame[1]_c [3]), .O(n31_adj_5659));
    defparam i14_4_lut_adj_1695.LUT_INIT = 16'h8000;
    SB_LUT4 select_787_Select_162_i2_4_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[2]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5311));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_162_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 select_787_Select_31_i2_3_lut (.I0(\data_out_frame[3][7] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5310));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_31_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1696 (.I0(\FRAME_MATCHER.i[4] ), .I1(\FRAME_MATCHER.i[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/coms.v(158[12:15])
    defparam i1_2_lut_adj_1696.LUT_INIT = 16'heeee;
    SB_LUT4 i22526_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(GND_net), .I3(GND_net), .O(n38266));
    defparam i22526_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1697 (.I0(n10_c), .I1(n56368), .I2(GND_net), 
            .I3(GND_net), .O(n55515));
    defparam i1_2_lut_adj_1697.LUT_INIT = 16'hbbbb;
    SB_LUT4 select_787_Select_30_i2_3_lut (.I0(\data_out_frame[3][6] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5309));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_30_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_4_lut_adj_1698 (.I0(\FRAME_MATCHER.i[0] ), .I1(\FRAME_MATCHER.i[4] ), 
            .I2(n25087), .I3(\FRAME_MATCHER.i [1]), .O(n5));
    defparam i1_3_lut_4_lut_adj_1698.LUT_INIT = 16'hfefc;
    SB_LUT4 select_787_Select_161_i2_4_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[1]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5308));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_161_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49671 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n66771));
    defparam byte_transmit_counter_0__bdd_4_lut_49671.LUT_INIT = 16'he4aa;
    SB_LUT4 n66771_bdd_4_lut (.I0(n66771), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n66774));
    defparam n66771_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1699 (.I0(\FRAME_MATCHER.i_31__N_2511 ), .I1(\r_SM_Main_2__N_3545[0] ), 
            .I2(n53), .I3(tx_active), .O(n25069));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_4_lut_adj_1699.LUT_INIT = 16'haa8a;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_49552 (.I0(byte_transmit_counter[1]), 
            .I1(n60294), .I2(n60295), .I3(byte_transmit_counter[2]), .O(n66603));
    defparam byte_transmit_counter_1__bdd_4_lut_49552.LUT_INIT = 16'he4aa;
    SB_LUT4 n66603_bdd_4_lut (.I0(n66603), .I1(n60004), .I2(n60003), .I3(byte_transmit_counter[2]), 
            .O(n66606));
    defparam n66603_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13066_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[16] [0]), 
            .I3(deadband[0]), .O(n28911));   // verilog/coms.v(148[4] 304[11])
    defparam i13066_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13073_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[13] [0]), 
            .I3(IntegralLimit[0]), .O(n28918));   // verilog/coms.v(148[4] 304[11])
    defparam i13073_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13074_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[3][0] ), 
            .I3(\Kp[0] ), .O(n28919));   // verilog/coms.v(148[4] 304[11])
    defparam i13074_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_28_i2_3_lut (.I0(\data_out_frame[3][4] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5306));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_28_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13075_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[5] [0]), 
            .I3(\Ki[0] ), .O(n28920));   // verilog/coms.v(148[4] 304[11])
    defparam i13075_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_84_i2_4_lut (.I0(\data_out_frame[10] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[12]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5448));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_84_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i1_2_lut_4_lut_adj_1700 (.I0(n771), .I1(\FRAME_MATCHER.i_31__N_2508 ), 
            .I2(n25069), .I3(\FRAME_MATCHER.i_31__N_2507 ), .O(n59705));   // verilog/coms.v(148[4] 304[11])
    defparam i1_2_lut_4_lut_adj_1700.LUT_INIT = 16'hfff4;
    SB_LUT4 i13079_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[10] [0]), 
            .I3(PWMLimit[0]), .O(n28924));   // verilog/coms.v(148[4] 304[11])
    defparam i13079_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_27_i2_3_lut (.I0(\data_out_frame[3][3] ), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(\FRAME_MATCHER.state_31__N_2612 [3]), .I3(GND_net), .O(n2_adj_5305));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_27_i2_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13764_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[8] [7]), 
            .I3(PWMLimit[23]), .O(n29609));   // verilog/coms.v(148[4] 304[11])
    defparam i13764_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1701 (.I0(control_mode[3]), .I1(control_mode[2]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5633));   // verilog/coms.v(130[12] 305[6])
    defparam i1_2_lut_adj_1701.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1702 (.I0(\FRAME_MATCHER.i_31__N_2509 ), .I1(\data_out_frame[10] [3]), 
            .I2(encoder1_position_scaled[11]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5447));   // verilog/coms.v(148[4] 304[11])
    defparam i1_4_lut_adj_1702.LUT_INIT = 16'ha088;
    SB_LUT4 i13765_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[8] [6]), 
            .I3(PWMLimit[22]), .O(n29610));   // verilog/coms.v(148[4] 304[11])
    defparam i13765_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i16_4_lut_adj_1703 (.I0(n31_adj_5659), .I1(n29_adj_5658), .I2(n59783), 
            .I3(n26), .O(\FRAME_MATCHER.state_31__N_2612 [3]));
    defparam i16_4_lut_adj_1703.LUT_INIT = 16'h0800;
    SB_LUT4 i13766_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[8] [5]), 
            .I3(PWMLimit[21]), .O(n29611));   // verilog/coms.v(148[4] 304[11])
    defparam i13766_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49538 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [1]), .I2(\data_out_frame[23] [1]), 
            .I3(byte_transmit_counter[1]), .O(n66591));
    defparam byte_transmit_counter_0__bdd_4_lut_49538.LUT_INIT = 16'he4aa;
    SB_LUT4 i17966_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[8] [4]), 
            .I3(PWMLimit[20]), .O(n29612));   // verilog/coms.v(148[4] 304[11])
    defparam i17966_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n66591_bdd_4_lut (.I0(n66591), .I1(\data_out_frame[21] [1]), 
            .I2(\data_out_frame[20] [1]), .I3(byte_transmit_counter[1]), 
            .O(n66594));
    defparam n66591_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13768_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[8] [3]), 
            .I3(PWMLimit[19]), .O(n29613));   // verilog/coms.v(148[4] 304[11])
    defparam i13768_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i18009_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[8] [2]), 
            .I3(PWMLimit[18]), .O(n29614));   // verilog/coms.v(148[4] 304[11])
    defparam i18009_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13770_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[8] [1]), 
            .I3(PWMLimit[17]), .O(n29615));   // verilog/coms.v(148[4] 304[11])
    defparam i13770_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_3_lut_adj_1704 (.I0(\FRAME_MATCHER.i[5] ), .I1(n73), 
            .I2(n55512), .I3(GND_net), .O(n27862));
    defparam i1_2_lut_3_lut_adj_1704.LUT_INIT = 16'hfbfb;
    SB_LUT4 select_787_Select_82_i2_4_lut (.I0(\data_out_frame[10] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[10]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5446));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_82_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13771_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[8] [0]), 
            .I3(PWMLimit[16]), .O(n29616));   // verilog/coms.v(148[4] 304[11])
    defparam i13771_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49520 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n66585));
    defparam byte_transmit_counter_0__bdd_4_lut_49520.LUT_INIT = 16'he4aa;
    SB_LUT4 i13772_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[9] [7]), 
            .I3(PWMLimit[15]), .O(n29617));   // verilog/coms.v(148[4] 304[11])
    defparam i13772_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 n66585_bdd_4_lut (.I0(n66585), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8][3] ), .I3(byte_transmit_counter[1]), 
            .O(n66588));
    defparam n66585_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13773_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[9] [6]), 
            .I3(PWMLimit[14]), .O(n29618));   // verilog/coms.v(148[4] 304[11])
    defparam i13773_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49515 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [2]), .I2(\data_out_frame[23] [2]), 
            .I3(byte_transmit_counter[1]), .O(n66579));
    defparam byte_transmit_counter_0__bdd_4_lut_49515.LUT_INIT = 16'he4aa;
    SB_LUT4 i13774_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[9] [5]), 
            .I3(PWMLimit[13]), .O(n29619));   // verilog/coms.v(148[4] 304[11])
    defparam i13774_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_81_i2_4_lut (.I0(\data_out_frame[10] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[9]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5445));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_81_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n66579_bdd_4_lut (.I0(n66579), .I1(\data_out_frame[21] [2]), 
            .I2(\data_out_frame[20] [2]), .I3(byte_transmit_counter[1]), 
            .O(n66582));
    defparam n66579_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14018_3_lut_4_lut (.I0(n8_adj_5430), .I1(n55507), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n29863));
    defparam i14018_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13775_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[9] [4]), 
            .I3(PWMLimit[12]), .O(n29620));   // verilog/coms.v(148[4] 304[11])
    defparam i13775_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13776_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[9] [3]), 
            .I3(PWMLimit[11]), .O(n29621));   // verilog/coms.v(148[4] 304[11])
    defparam i13776_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13777_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[9] [2]), 
            .I3(PWMLimit[10]), .O(n29622));   // verilog/coms.v(148[4] 304[11])
    defparam i13777_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13778_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[9] [1]), 
            .I3(PWMLimit[9]), .O(n29623));   // verilog/coms.v(148[4] 304[11])
    defparam i13778_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49510 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n66573));
    defparam byte_transmit_counter_0__bdd_4_lut_49510.LUT_INIT = 16'he4aa;
    SB_LUT4 n66573_bdd_4_lut (.I0(n66573), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n66576));
    defparam n66573_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13779_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[9] [0]), 
            .I3(PWMLimit[8]), .O(n29624));   // verilog/coms.v(148[4] 304[11])
    defparam i13779_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13780_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[10] [7]), 
            .I3(PWMLimit[7]), .O(n29625));   // verilog/coms.v(148[4] 304[11])
    defparam i13780_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13781_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[10] [6]), 
            .I3(PWMLimit[6]), .O(n29626));   // verilog/coms.v(148[4] 304[11])
    defparam i13781_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13782_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[10] [5]), 
            .I3(PWMLimit[5]), .O(n29627));   // verilog/coms.v(148[4] 304[11])
    defparam i13782_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13783_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[10] [4]), 
            .I3(PWMLimit[4]), .O(n29628));   // verilog/coms.v(148[4] 304[11])
    defparam i13783_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13784_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[10] [3]), 
            .I3(PWMLimit[3]), .O(n29629));   // verilog/coms.v(148[4] 304[11])
    defparam i13784_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_80_i2_4_lut (.I0(\data_out_frame[10] [0]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[8]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5444));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_80_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13785_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[10] [2]), 
            .I3(PWMLimit[2]), .O(n29630));   // verilog/coms.v(148[4] 304[11])
    defparam i13785_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13786_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[10] [1]), 
            .I3(PWMLimit[1]), .O(n29631));   // verilog/coms.v(148[4] 304[11])
    defparam i13786_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13833_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[4] [7]), 
            .I3(\Ki[15] ), .O(n29678));   // verilog/coms.v(148[4] 304[11])
    defparam i13833_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i18620_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[4] [6]), 
            .I3(\Ki[14] ), .O(n29679));   // verilog/coms.v(148[4] 304[11])
    defparam i18620_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13835_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[4] [5]), 
            .I3(\Ki[13] ), .O(n29680));   // verilog/coms.v(148[4] 304[11])
    defparam i13835_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13836_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[4] [4]), 
            .I3(\Ki[12] ), .O(n29681));   // verilog/coms.v(148[4] 304[11])
    defparam i13836_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_79_i2_4_lut (.I0(\data_out_frame[9] [7]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[23]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5443));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_79_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13837_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[4] [3]), 
            .I3(\Ki[11] ), .O(n29682));   // verilog/coms.v(148[4] 304[11])
    defparam i13837_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13698_3_lut_4_lut (.I0(n27860), .I1(reset), .I2(rx_data[7]), 
            .I3(\data_in_frame[22] [7]), .O(n29543));
    defparam i13698_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_787_Select_78_i2_4_lut (.I0(\data_out_frame[9] [6]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[22]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5442));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_78_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13838_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[4] [2]), 
            .I3(\Ki[10] ), .O(n29683));   // verilog/coms.v(148[4] 304[11])
    defparam i13838_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13839_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[4] [1]), 
            .I3(\Ki[9] ), .O(n29684));   // verilog/coms.v(148[4] 304[11])
    defparam i13839_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13840_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[4] [0]), 
            .I3(\Ki[8] ), .O(n29685));   // verilog/coms.v(148[4] 304[11])
    defparam i13840_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13841_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[5] [7]), 
            .I3(\Ki[7] ), .O(n29686));   // verilog/coms.v(148[4] 304[11])
    defparam i13841_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_77_i2_4_lut (.I0(\data_out_frame[9] [5]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[21]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5441));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_77_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13842_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[5] [6]), 
            .I3(\Ki[6] ), .O(n29687));   // verilog/coms.v(148[4] 304[11])
    defparam i13842_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13843_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[5] [5]), 
            .I3(\Ki[5] ), .O(n29688));   // verilog/coms.v(148[4] 304[11])
    defparam i13843_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_160_i2_4_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[0]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5303));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_160_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i48243_3_lut (.I0(n66750), .I1(n66558), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n65305));
    defparam i48243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13844_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[5] [4]), 
            .I3(\Ki[4] ), .O(n29689));   // verilog/coms.v(148[4] 304[11])
    defparam i13844_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13845_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[5] [3]), 
            .I3(\Ki[3] ), .O(n29690));   // verilog/coms.v(148[4] 304[11])
    defparam i13845_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i48244_4_lut (.I0(n65305), .I1(n66792), .I2(byte_transmit_counter_c[3]), 
            .I3(byte_transmit_counter[2]), .O(n65306));
    defparam i48244_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13695_3_lut_4_lut (.I0(n27860), .I1(reset), .I2(rx_data[6]), 
            .I3(\data_in_frame[22] [6]), .O(n29540));
    defparam i13695_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_49711 (.I0(byte_transmit_counter_c[3]), 
            .I1(n66546), .I2(n63125), .I3(byte_transmit_counter_c[4]), 
            .O(n66561));
    defparam byte_transmit_counter_3__bdd_4_lut_49711.LUT_INIT = 16'he4aa;
    SB_LUT4 n66561_bdd_4_lut (.I0(n66561), .I1(n14_adj_5656), .I2(n60044), 
            .I3(byte_transmit_counter_c[4]), .O(tx_data[4]));
    defparam n66561_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i42997_3_lut (.I0(n66630), .I1(n65306), .I2(byte_transmit_counter_c[4]), 
            .I3(GND_net), .O(tx_data[3]));
    defparam i42997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18625_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[5] [2]), 
            .I3(\Ki[2] ), .O(n29691));   // verilog/coms.v(148[4] 304[11])
    defparam i18625_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_76_i2_4_lut (.I0(\data_out_frame[9] [4]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[20]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5440));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_76_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13692_3_lut_4_lut (.I0(n27860), .I1(reset), .I2(rx_data[5]), 
            .I3(\data_in_frame[22] [5]), .O(n29537));
    defparam i13692_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18621_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[5] [1]), 
            .I3(\Ki[1] ), .O(n29692));   // verilog/coms.v(148[4] 304[11])
    defparam i18621_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13848_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[2]_c [7]), 
            .I3(\Kp[15] ), .O(n29693));   // verilog/coms.v(148[4] 304[11])
    defparam i13848_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49505 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [3]), .I2(\data_out_frame[23] [3]), 
            .I3(byte_transmit_counter[1]), .O(n66555));
    defparam byte_transmit_counter_0__bdd_4_lut_49505.LUT_INIT = 16'he4aa;
    SB_LUT4 i13849_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[2]_c [6]), 
            .I3(\Kp[14] ), .O(n29694));   // verilog/coms.v(148[4] 304[11])
    defparam i13849_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13850_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[2]_c [5]), 
            .I3(\Kp[13] ), .O(n29695));   // verilog/coms.v(148[4] 304[11])
    defparam i13850_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13851_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[2]_c [4]), 
            .I3(\Kp[12] ), .O(n29696));   // verilog/coms.v(148[4] 304[11])
    defparam i13851_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13852_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[2]_c [3]), 
            .I3(\Kp[11] ), .O(n29697));   // verilog/coms.v(148[4] 304[11])
    defparam i13852_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13688_3_lut_4_lut (.I0(n27860), .I1(reset), .I2(rx_data[4]), 
            .I3(\data_in_frame[22] [4]), .O(n29533));
    defparam i13688_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n66555_bdd_4_lut (.I0(n66555), .I1(\data_out_frame[21] [3]), 
            .I2(\data_out_frame[20] [3]), .I3(byte_transmit_counter[1]), 
            .O(n66558));
    defparam n66555_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13853_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[2]_c [2]), 
            .I3(\Kp[10] ), .O(n29698));   // verilog/coms.v(148[4] 304[11])
    defparam i13853_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13685_3_lut_4_lut (.I0(n27860), .I1(reset), .I2(rx_data[3]), 
            .I3(\data_in_frame[22] [3]), .O(n29530));
    defparam i13685_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13854_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[2]_c [1]), 
            .I3(\Kp[9] ), .O(n29699));   // verilog/coms.v(148[4] 304[11])
    defparam i13854_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13855_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[2] [0]), 
            .I3(\Kp[8] ), .O(n29700));   // verilog/coms.v(148[4] 304[11])
    defparam i13855_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13856_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[3][7] ), 
            .I3(\Kp[7] ), .O(n29701));   // verilog/coms.v(148[4] 304[11])
    defparam i13856_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13857_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[3][6] ), 
            .I3(\Kp[6] ), .O(n29702));   // verilog/coms.v(148[4] 304[11])
    defparam i13857_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13858_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[3][5] ), 
            .I3(\Kp[5] ), .O(n29703));   // verilog/coms.v(148[4] 304[11])
    defparam i13858_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i18810_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[3] [4]), 
            .I3(\Kp[4] ), .O(n29704));   // verilog/coms.v(148[4] 304[11])
    defparam i18810_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_75_i2_4_lut (.I0(\data_out_frame[9] [3]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[19]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5439));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_75_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13860_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[3][3] ), 
            .I3(\Kp[3] ), .O(n29705));   // verilog/coms.v(148[4] 304[11])
    defparam i13860_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13861_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[3] [2]), 
            .I3(\Kp[2] ), .O(n29706));   // verilog/coms.v(148[4] 304[11])
    defparam i13861_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_49492 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [0]), .I2(\data_out_frame[23] [0]), 
            .I3(byte_transmit_counter[1]), .O(n66549));
    defparam byte_transmit_counter_0__bdd_4_lut_49492.LUT_INIT = 16'he4aa;
    SB_LUT4 i13862_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[3] [1]), 
            .I3(\Kp[1] ), .O(n29707));   // verilog/coms.v(148[4] 304[11])
    defparam i13862_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_74_i2_4_lut (.I0(\data_out_frame[9] [2]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[18]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5438));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_74_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i11_4_lut_4_lut_adj_1705 (.I0(n27860), .I1(reset), .I2(rx_data[2]), 
            .I3(\data_in_frame[22] [2]), .O(n54663));
    defparam i11_4_lut_4_lut_adj_1705.LUT_INIT = 16'hfe10;
    SB_LUT4 i13863_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[11] [7]), 
            .I3(IntegralLimit[23]), .O(n29708));   // verilog/coms.v(148[4] 304[11])
    defparam i13863_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13679_3_lut_4_lut (.I0(n27860), .I1(reset), .I2(rx_data[1]), 
            .I3(\data_in_frame[22] [1]), .O(n29524));
    defparam i13679_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n66549_bdd_4_lut (.I0(n66549), .I1(\data_out_frame[21] [0]), 
            .I2(\data_out_frame[20] [0]), .I3(byte_transmit_counter[1]), 
            .O(n66552));
    defparam n66549_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1706 (.I0(\FRAME_MATCHER.i[0] ), .I1(n38266), 
            .I2(n3484), .I3(n37097), .O(n27860));
    defparam i1_2_lut_4_lut_adj_1706.LUT_INIT = 16'hbfff;
    SB_LUT4 i13864_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[11] [6]), 
            .I3(IntegralLimit[22]), .O(n29709));   // verilog/coms.v(148[4] 304[11])
    defparam i13864_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13865_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[11] [5]), 
            .I3(IntegralLimit[21]), .O(n29710));   // verilog/coms.v(148[4] 304[11])
    defparam i13865_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_73_i2_4_lut (.I0(\data_out_frame[9] [1]), .I1(\FRAME_MATCHER.i_31__N_2509 ), 
            .I2(encoder1_position_scaled[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5437));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_73_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13866_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[11] [4]), 
            .I3(IntegralLimit[20]), .O(n29711));   // verilog/coms.v(148[4] 304[11])
    defparam i13866_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13867_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[11] [3]), 
            .I3(IntegralLimit[19]), .O(n29712));   // verilog/coms.v(148[4] 304[11])
    defparam i13867_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_49529 (.I0(byte_transmit_counter[1]), 
            .I1(n60081), .I2(n60082), .I3(byte_transmit_counter[2]), .O(n66543));
    defparam byte_transmit_counter_1__bdd_4_lut_49529.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1707 (.I0(reset), .I1(n10_c), .I2(n56368), 
            .I3(GND_net), .O(n55507));
    defparam i1_2_lut_3_lut_adj_1707.LUT_INIT = 16'hefef;
    SB_LUT4 i13868_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[11] [2]), 
            .I3(IntegralLimit[18]), .O(n29713));   // verilog/coms.v(148[4] 304[11])
    defparam i13868_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13869_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[11] [1]), 
            .I3(IntegralLimit[17]), .O(n29714));   // verilog/coms.v(148[4] 304[11])
    defparam i13869_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i11_3_lut_4_lut_adj_1708 (.I0(n27860), .I1(reset), .I2(\data_in_frame[22] [0]), 
            .I3(rx_data[0]), .O(n54577));
    defparam i11_3_lut_4_lut_adj_1708.LUT_INIT = 16'hf1e0;
    SB_LUT4 select_787_Select_159_i2_4_lut (.I0(\data_out_frame[19] [7]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[15]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5302));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_159_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13870_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[11] [0]), 
            .I3(IntegralLimit[16]), .O(n29715));   // verilog/coms.v(148[4] 304[11])
    defparam i13870_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13871_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[12] [7]), 
            .I3(IntegralLimit[15]), .O(n29716));   // verilog/coms.v(148[4] 304[11])
    defparam i13871_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_145_i2_4_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[17]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_145_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 n66543_bdd_4_lut (.I0(n66543), .I1(n60124), .I2(n60123), .I3(byte_transmit_counter[2]), 
            .O(n66546));
    defparam n66543_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13872_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[12] [6]), 
            .I3(IntegralLimit[14]), .O(n29717));   // verilog/coms.v(148[4] 304[11])
    defparam i13872_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i13873_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[12] [5]), 
            .I3(IntegralLimit[13]), .O(n29718));   // verilog/coms.v(148[4] 304[11])
    defparam i13873_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 select_787_Select_158_i2_4_lut (.I0(\data_out_frame[19] [6]), 
            .I1(\FRAME_MATCHER.i_31__N_2509 ), .I2(displacement[14]), .I3(\FRAME_MATCHER.state_31__N_2612 [3]), 
            .O(n2_adj_5301));   // verilog/coms.v(148[4] 304[11])
    defparam select_787_Select_158_i2_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i13874_3_lut_4_lut (.I0(Kp_23__N_1748), .I1(n32097), .I2(\data_in_frame[12] [4]), 
            .I3(IntegralLimit[12]), .O(n29719));   // verilog/coms.v(148[4] 304[11])
    defparam i13874_3_lut_4_lut.LUT_INIT = 16'hf780;
    uart_tx tx (.tx_data({tx_data}), .clk16MHz(clk16MHz), .r_SM_Main({Open_50, 
            \r_SM_Main[1] , Open_51}), .GND_net(GND_net), .r_Clock_Count({r_Clock_Count}), 
            .n39972(n39972), .tx_o(tx_o), .n20722(n20722), .\r_SM_Main[0] (\r_SM_Main[0] ), 
            .VCC_net(VCC_net), .n27315(n27315), .n23(n23), .\o_Rx_DV_N_3488[12] (\o_Rx_DV_N_3488[12] ), 
            .n5228(n5228), .\o_Rx_DV_N_3488[24] (\o_Rx_DV_N_3488[24] ), 
            .n27(n27), .n29(n29), .n39919(n39919), .n29589(n29589), 
            .\r_Bit_Index[0] (\r_Bit_Index[0] ), .n51433(n51433), .tx_active(tx_active), 
            .n39937(n39937), .n57036(n57036), .n31(n31), .\r_SM_Main_2__N_3545[0] (\r_SM_Main_2__N_3545[0] ), 
            .n58374(n58374), .n58502(n58502), .o_Tx_Serial_N_3598(o_Tx_Serial_N_3598), 
            .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(110[25:94])
    uart_rx rx (.baudrate({baudrate}), .GND_net(GND_net), .VCC_net(VCC_net), 
            .r_SM_Main({r_SM_Main}), .clk16MHz(clk16MHz), .r_Rx_Data(r_Rx_Data), 
            .RX_N_2(RX_N_2), .r_Clock_Count({r_Clock_Count_adj_20}), .\o_Rx_DV_N_3488[24] (\o_Rx_DV_N_3488[24] ), 
            .n27(n27), .n25108(n25108), .n29(n29), .n23(n23), .\o_Rx_DV_N_3488[12] (\o_Rx_DV_N_3488[12] ), 
            .n5225(n5225), .\o_Rx_DV_N_3488[8] (\o_Rx_DV_N_3488[8] ), .\o_Rx_DV_N_3488[7] (\o_Rx_DV_N_3488[7] ), 
            .\o_Rx_DV_N_3488[6] (\o_Rx_DV_N_3488[6] ), .\o_Rx_DV_N_3488[5] (\o_Rx_DV_N_3488[5] ), 
            .\o_Rx_DV_N_3488[4] (\o_Rx_DV_N_3488[4] ), .\o_Rx_DV_N_3488[3] (\o_Rx_DV_N_3488[3] ), 
            .\o_Rx_DV_N_3488[2] (\o_Rx_DV_N_3488[2] ), .\o_Rx_DV_N_3488[1] (\o_Rx_DV_N_3488[1] ), 
            .\o_Rx_DV_N_3488[0] (\o_Rx_DV_N_3488[0] ), .n27312(n27312), 
            .n29592(n29592), .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_17 ), 
            .n51425(n51425), .rx_data_ready(rx_data_ready), .n29596(n29596), 
            .rx_data({rx_data}), .n29582(n29582), .n29581(n29581), .n29580(n29580), 
            .n29578(n29578), .n29577(n29577), .n29576(n29576), .n29575(n29575), 
            .\r_SM_Main_2__N_3446[1] (\r_SM_Main_2__N_3446[1] ), .n56281(n56281), 
            .n6(n6_adj_18), .n55184(n55184), .n58618(n58618), .n4(n4_adj_19), 
            .n27308(n27308), .n58594(n58594), .n58896(n58896), .n58898(n58898), 
            .n58932(n58932), .n58844(n58844), .n58970(n58970), .n58934(n58934), 
            .n58880(n58880), .n58952(n58952)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(96[25:68])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (tx_data, clk16MHz, r_SM_Main, GND_net, r_Clock_Count, 
            n39972, tx_o, n20722, \r_SM_Main[0] , VCC_net, n27315, 
            n23, \o_Rx_DV_N_3488[12] , n5228, \o_Rx_DV_N_3488[24] , 
            n27, n29, n39919, n29589, \r_Bit_Index[0] , n51433, 
            tx_active, n39937, n57036, n31, \r_SM_Main_2__N_3545[0] , 
            n58374, n58502, o_Tx_Serial_N_3598, tx_enable) /* synthesis syn_module_defined=1 */ ;
    input [7:0]tx_data;
    input clk16MHz;
    output [2:0]r_SM_Main;
    input GND_net;
    output [8:0]r_Clock_Count;
    input n39972;
    output tx_o;
    input n20722;
    output \r_SM_Main[0] ;
    input VCC_net;
    output n27315;
    input n23;
    input \o_Rx_DV_N_3488[12] ;
    input n5228;
    input \o_Rx_DV_N_3488[24] ;
    input n27;
    input n29;
    output n39919;
    input n29589;
    output \r_Bit_Index[0] ;
    input n51433;
    output tx_active;
    input n39937;
    output n57036;
    output n31;
    input \r_SM_Main_2__N_3545[0] ;
    output n58374;
    output n58502;
    output o_Tx_Serial_N_3598;
    output tx_enable;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(41[6:14])
    
    wire n22335;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(35[16:25])
    
    wire n3;
    wire [2:0]r_SM_Main_c;   // verilog/uart_tx.v(32[16:25])
    wire [8:0]n41;
    
    wire n49282, n49281, n1, n49280, n49279, n49278, n49277, n49276, 
        n49275, n28647;
    wire [2:0]n460;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(34[16:27])
    
    wire n28355, n58508, n63101, n63098, n67139, n58574, n58580, 
        n56396, n59991, n59992, n59995, n59994, n14, n15, n66597;
    
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk16MHz), .E(n22335), 
            .D(tx_data[7]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3), .R(r_SM_Main_c[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk16MHz), .E(n22335), 
            .D(tx_data[6]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk16MHz), .E(n22335), 
            .D(tx_data[5]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk16MHz), .E(n22335), 
            .D(tx_data[4]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk16MHz), .E(n22335), 
            .D(tx_data[3]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk16MHz), .E(n22335), 
            .D(tx_data[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk16MHz), .E(n22335), 
            .D(tx_data[1]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 r_Clock_Count_2056_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n49282), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2056_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n49281), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_9 (.CI(n49281), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n49282));
    SB_DFFE o_Tx_Serial_51 (.Q(tx_o), .C(clk16MHz), .E(n1), .D(n39972));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 r_Clock_Count_2056_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n49280), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_8 (.CI(n49280), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n49281));
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk16MHz), .E(n22335), 
            .D(tx_data[0]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(\r_SM_Main[0] ), .C(clk16MHz), .D(n20722), 
            .R(r_SM_Main_c[2]));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 r_Clock_Count_2056_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n49279), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_7 (.CI(n49279), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n49280));
    SB_LUT4 r_Clock_Count_2056_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n49278), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_6 (.CI(n49278), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n49279));
    SB_LUT4 r_Clock_Count_2056_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n49277), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_5 (.CI(n49277), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n49278));
    SB_LUT4 r_Clock_Count_2056_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n49276), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_4 (.CI(n49276), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n49277));
    SB_LUT4 r_Clock_Count_2056_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n49275), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_3 (.CI(n49275), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n49276));
    SB_LUT4 r_Clock_Count_2056_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2056_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2056_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n49275));
    SB_DFFESR r_Clock_Count_2056__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n1), .D(n41[0]), .R(n28647));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i8 (.Q(r_Clock_Count[8]), .C(clk16MHz), 
            .E(n1), .D(n41[8]), .R(n28647));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n1), .D(n41[7]), .R(n28647));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n1), .D(n41[6]), .R(n28647));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n1), .D(n41[5]), .R(n28647));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n1), .D(n41[4]), .R(n28647));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n1), .D(n41[3]), .R(n28647));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n1), .D(n41[2]), .R(n28647));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Clock_Count_2056__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n1), .D(n41[1]), .R(n28647));   // verilog/uart_tx.v(119[34:51])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n27315), 
            .D(n460[1]), .R(n28355));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n27315), 
            .D(n460[2]), .R(n28355));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i1_4_lut (.I0(n23), .I1(\o_Rx_DV_N_3488[12] ), .I2(n5228), 
            .I3(\r_SM_Main[0] ), .O(n58508));
    defparam i1_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1086 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n27), .I2(n29), 
            .I3(n58508), .O(n39919));
    defparam i1_4_lut_adj_1086.LUT_INIT = 16'h0100;
    SB_LUT4 i46792_3_lut (.I0(\r_SM_Main[0] ), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n5228), .I3(GND_net), .O(n63101));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i46792_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i46787_4_lut (.I0(n63101), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n63098));   // verilog/uart_tx.v(44[7] 143[14])
    defparam i46787_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(n39919), .I1(n63098), 
            .I2(r_SM_Main[1]), .I3(n27), .O(n3));   // verilog/uart_tx.v(44[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'hfaca;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main_c[2]), .C(clk16MHz), .D(n67139));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .D(n29589));   // verilog/uart_tx.v(41[10] 144[8])
    SB_DFF r_Tx_Active_53 (.Q(tx_active), .C(clk16MHz), .D(n51433));   // verilog/uart_tx.v(41[10] 144[8])
    SB_LUT4 i2336_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n460[2]));   // verilog/uart_tx.v(99[36:51])
    defparam i2336_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i39279_rep_28_2_lut (.I0(n39937), .I1(r_SM_Main[1]), .I2(GND_net), 
            .I3(GND_net), .O(n57036));
    defparam i39279_rep_28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut (.I0(\o_Rx_DV_N_3488[12] ), .I1(n5228), .I2(n31), 
            .I3(GND_net), .O(n58574));
    defparam i1_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_4_lut_adj_1087 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n58574), .O(n58580));
    defparam i1_4_lut_adj_1087.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1088 (.I0(n58580), .I1(n56396), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n28355));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i1_4_lut_adj_1088.LUT_INIT = 16'h0323;
    SB_LUT4 i2329_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n460[1]));   // verilog/uart_tx.v(99[36:51])
    defparam i2329_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i42929_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n59991));
    defparam i42929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42930_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n59992));
    defparam i42930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42933_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n59995));
    defparam i42933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42932_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n59994));
    defparam i42932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1089 (.I0(\r_Bit_Index[0] ), .I1(r_Bit_Index[1]), 
            .I2(r_Bit_Index[2]), .I3(GND_net), .O(n31));   // verilog/uart_tx.v(41[10] 144[8])
    defparam i1_3_lut_adj_1089.LUT_INIT = 16'h8080;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main_c[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut (.I0(\r_SM_Main_2__N_3545[0] ), .I1(r_SM_Main_c[2]), 
            .I2(\r_SM_Main[0] ), .I3(r_SM_Main[1]), .O(n22335));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i49319_4_lut (.I0(r_SM_Main_c[2]), .I1(n39937), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main[0] ), .O(n28647));
    defparam i49319_4_lut.LUT_INIT = 16'h1115;
    SB_LUT4 i5_3_lut (.I0(\r_SM_Main[0] ), .I1(\o_Rx_DV_N_3488[24] ), .I2(n27), 
            .I3(GND_net), .O(n14));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3488[12] ), .I2(n23), .I3(n5228), 
            .O(n15));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(n1), .I2(n14), .I3(r_SM_Main[1]), 
            .O(n67139));
    defparam i8_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main_c[2]), .I2(\r_SM_Main[0] ), 
            .I3(n31), .O(n58374));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0301;
    SB_LUT4 i1_4_lut_4_lut (.I0(\r_SM_Main[0] ), .I1(r_SM_Main_c[2]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3545[0] ), .O(n58502));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h3130;
    SB_LUT4 i49230_2_lut_4_lut (.I0(n39937), .I1(r_SM_Main[1]), .I2(r_SM_Main_c[2]), 
            .I3(\r_SM_Main[0] ), .O(n27315));
    defparam i49230_2_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i39389_2_lut (.I0(r_SM_Main_c[2]), .I1(\r_SM_Main[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n56396));
    defparam i39389_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n59994), 
            .I2(n59995), .I3(r_Bit_Index[2]), .O(n66597));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n66597_bdd_4_lut (.I0(n66597), .I1(n59992), .I2(n59991), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_3598));
    defparam n66597_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(39[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (baudrate, GND_net, VCC_net, r_SM_Main, clk16MHz, r_Rx_Data, 
            RX_N_2, r_Clock_Count, \o_Rx_DV_N_3488[24] , n27, n25108, 
            n29, n23, \o_Rx_DV_N_3488[12] , n5225, \o_Rx_DV_N_3488[8] , 
            \o_Rx_DV_N_3488[7] , \o_Rx_DV_N_3488[6] , \o_Rx_DV_N_3488[5] , 
            \o_Rx_DV_N_3488[4] , \o_Rx_DV_N_3488[3] , \o_Rx_DV_N_3488[2] , 
            \o_Rx_DV_N_3488[1] , \o_Rx_DV_N_3488[0] , n27312, n29592, 
            \r_Bit_Index[0] , n51425, rx_data_ready, n29596, rx_data, 
            n29582, n29581, n29580, n29578, n29577, n29576, n29575, 
            \r_SM_Main_2__N_3446[1] , n56281, n6, n55184, n58618, 
            n4, n27308, n58594, n58896, n58898, n58932, n58844, 
            n58970, n58934, n58880, n58952) /* synthesis syn_module_defined=1 */ ;
    input [31:0]baudrate;
    input GND_net;
    input VCC_net;
    output [2:0]r_SM_Main;
    input clk16MHz;
    output r_Rx_Data;
    input RX_N_2;
    output [7:0]r_Clock_Count;
    output \o_Rx_DV_N_3488[24] ;
    output n27;
    output n25108;
    output n29;
    output n23;
    output \o_Rx_DV_N_3488[12] ;
    input n5225;
    output \o_Rx_DV_N_3488[8] ;
    output \o_Rx_DV_N_3488[7] ;
    output \o_Rx_DV_N_3488[6] ;
    output \o_Rx_DV_N_3488[5] ;
    output \o_Rx_DV_N_3488[4] ;
    output \o_Rx_DV_N_3488[3] ;
    output \o_Rx_DV_N_3488[2] ;
    output \o_Rx_DV_N_3488[1] ;
    output \o_Rx_DV_N_3488[0] ;
    output n27312;
    input n29592;
    output \r_Bit_Index[0] ;
    input n51425;
    output rx_data_ready;
    input n29596;
    output [7:0]rx_data;
    input n29582;
    input n29581;
    input n29580;
    input n29578;
    input n29577;
    input n29576;
    input n29575;
    input \r_SM_Main_2__N_3446[1] ;
    output n56281;
    output n6;
    output n55184;
    input n58618;
    output n4;
    output n27308;
    output n58594;
    input n58896;
    output n58898;
    input n58932;
    output n58844;
    output n58970;
    output n58934;
    output n58880;
    output n58952;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(41[6:14])
    
    wire n65772, n37, n65559, n2723, n27_c, n2722, n29_c, n2721, 
        n31, n2610;
    wire [23:0]n8184;
    wire [23:0]n294;
    
    wire n2727;
    wire [23:0]n8158;
    
    wire n2487, n1460, n48951, n48952, n2611, n2728, n66107, n41, 
        n63231, n66235, n2612, n2729, n2488, n1011, n48950, n17, 
        n19, n2607, n2724, n2489, n856, n48949, n2608, n2725, 
        n2609, n2726, n2366;
    wire [23:0]n8132;
    
    wire n21, n23_c, n25, n2490, n698, n48948, n2491, n858, 
        n48947, n2718, n37_adj_5013, n58480, n538, n56585, n2353, 
        n2638, n48946, n2354, n2519, n48945, n63963, n64949, n65383, 
        n65375, n35, n33, n63970, n2730, n14, n65595, n39, n65596, 
        n2100, n66236, n22, n45, n40, n43, n41_adj_5014, n63952, 
        n20, n63950, n65575, n64475, n2099, n66187, n2098, n48, 
        n18, n26, n16, n63997, n65981, n59304, n65982, n65854, 
        n65717, n2355, n2397, n48944, n2356, n2272, n48943, n66051, 
        n64473, n66053, n59254, n59302, n58984, n59312, n59308, 
        n59310, n25187, n2357, n2144, n48942, n2358, n2013, n48941, 
        n2476, n2596, n21311, n9620, n44, n2477, n2597, n2481, 
        n2601, n2359, n1879, n48940, n37_adj_5015, n2478, n2598, 
        n2360, n1742, n48939, n43_adj_5016, n2480, n2600, n39_adj_5017, 
        n2479, n2599, n2361, n1602, n48938, n59226, n59228, n41_adj_5018, 
        n2482, n2602, n2362, n1459, n48937, n59824, n2484, n2604, 
        n2483, n2603, n59174, n59954, n58804, n31_adj_5019, n33_adj_5020, 
        n35_adj_5021, n2485, n2605, n2486, n2606, n59890, n27_adj_5022, 
        n2363, n48936, n29_adj_5023, n56344, n59392, n58832, n2364, 
        n48935, n19_adj_5024, n21_adj_5025, n2365, n48934, n59886, 
        n59888, n59810, n59964, n63384, n66281, n23_adj_5026, n25_adj_5027, 
        n17_adj_5028, n64091, n64078, n65731, n16_adj_5029, n65605, 
        n65606, n64087, n64967, n22_adj_5030, n65573, n64465, n48_adj_5031, 
        n25229, n20_adj_5032, n28, n59238, n38422, n59096, n18_adj_5033, 
        n64068, n65979, n57124, n57547, n62993, n65980, n48933, 
        n59240, n59170, n62994, n65856, n64971, n65603, n59692, 
        n56317, n64463, n66138, n2367, n48932, n56321, n66139, 
        n25205, n56573, n804, n21309, n39_adj_5034, n45_adj_5035, 
        n43_adj_5036, n41_adj_5037, n33_adj_5038, n35_adj_5039, n37_adj_5040, 
        n29_adj_5041, n31_adj_5042, n21_adj_5043, n23_adj_5044, n25_adj_5045, 
        n27_adj_5046, n58478, n56589, n19_adj_5047, n64137, n64133, 
        n65739, n18_adj_5048, n65609;
    wire [23:0]n8106;
    
    wire n2227, n48931, n65610, n64135, n65005, n24, n26_adj_5049, 
        n64459, n2228, n48930, n22_adj_5050, n30, n20_adj_5051, 
        n64125, n65977, n65978, n65858, n44_adj_5052, n803, n65007, 
        n65570, n64457, n65572, n46, n56323;
    wire [23:0]n7976;
    
    wire n1552, n48662, n960, n9784, n21323, n21325, n2229, n48929, 
        n1553, n48661, n2230, n48928, n2231, n48927, n1554, n48660, 
        n2232, n48926, n1555, n48659, n2233, n48925, n2234, n48924, 
        n959, n3, r_Rx_Data_R, n2235, n48923, n9791, n46_adj_5053, 
        n2236, n48922, n1111, n1556, n48658, n2237, n48921, n2238, 
        n48920, n1557, n48657, n1558, n48656, n59946, n56569, 
        n2239, n48919, n1559, n48655, n2240, n48918, n1560, n48654, 
        n58476, n56593;
    wire [23:0]n7898;
    
    wire n1261;
    wire [23:0]n7924;
    
    wire n1408;
    wire [23:0]n7950;
    
    wire n1693;
    wire [23:0]n8002;
    
    wire n1831;
    wire [23:0]n8028;
    
    wire n1966;
    wire [7:0]n1;
    
    wire n49243, n49242;
    wire [23:0]n8054;
    
    wire n49241, n49240, n49239, n49238, n49237;
    wire [23:0]n8080;
    
    wire n59252, n59296, n48406, n48405, n58448, n59294, n59202, 
        n59004, n59974, n48404, n58524, n25202, n59012, n59008, 
        n59010, n59030, n59020, n59016, n59018, n59014, n59032, 
        n48403;
    wire [24:0]o_Rx_DV_N_3488;
    
    wire n3_adj_5063, n63088, n48402, n58522, n55210, n63094, n63085, 
        n63091, n48401, n58520, n48400, n48399, n58518, n63390, 
        n42_adj_5064, n48398, n58516, n48626, n48397, n58446, n1409, 
        n48625, n1410, n48624, n48396, n58514, n48395, n1411, 
        n48623, n48895, n48394, n42_adj_5065, n1113, n48894, n1412, 
        n48622, n1413, n48621, n48393, n48893, n48392, n1414, 
        n48620, n48391, n2101, n48892, n1415, n48619, n58472, 
        n56611, n48390, n48389, n59874, n2102, n48891, n48618, 
        n1262, n48617, n48388, n48387, n1263, n48616, n2103, n48890, 
        n48386, n59872, n59248, n1264, n48615, n48385, n59812, 
        n59926, n59968, n2104, n48889, n1265, n48614, n1695, n1833, 
        n1968, n43_adj_5066, n23_adj_5067, n29_adj_5068, n27_adj_5069, 
        n25_adj_5070, n63217, n35_adj_5071, n33_adj_5072, n31_adj_5073, 
        n63211, n22_adj_5074, n28_adj_5075, n30_adj_5076, n26_adj_5077, 
        n37_adj_5078, n34, n24_adj_5079, n63207, n66109, n2713, 
        n58484, n2845, n1266, n48613, n48384, n39_adj_5080, n66110, 
        n41_adj_5081, n65988, n65437, n63213, n65761, n2105, n48888, 
        n2106, n48887, n1267, n48612, n48383, n2107, n48886, n2108, 
        n48885, n58470, n56615, n2109, n48884, n57452, n42_adj_5082, 
        n2110, n27426, n28645, n66013, n66014, n48_adj_5083, n48602, 
        n1112, n48601;
    wire [23:0]n8314;
    
    wire n3151, n3186, n49090, n3152, n3082, n49089, n3153, n3188, 
        n49088, n3154, n3084, n49087, n3155, n2977, n49086, n3156, 
        n2867, n49085, n3157, n2754, n49084, n48600, n1114, n48599, 
        n3158, n49083, n3159, n49082, n3160, n49081, n3161, n49080, 
        n3162, n49079, n3163, n49078, n3164, n49077, n3165, n49076, 
        n3166, n49075, n3167, n49074, n3168, n49073, n3169, n49072, 
        n3170, n49071, n3171, n49070, n3172, n49069, n1115, n48598, 
        n1116, n48597, n58492, n49068, n56561;
    wire [23:0]n8288;
    
    wire n3046, n49067, n3047, n49066, n3048, n49065, n3049, n49064, 
        n3050, n49063, n3051, n49062, n3052, n49061, n58468, n56619, 
        n3053, n49060, n3054, n49059, n3055, n49058, n3056, n49057, 
        n25199, n3057, n49056, n3058, n49055, n3059, n49054, n3060, 
        n49053, n21_adj_5084, n27_adj_5085, n25_adj_5086, n23_adj_5087, 
        n63184, n3061, n49052, n3062, n49051, n3063, n49050, n33_adj_5088, 
        n31_adj_5089, n29_adj_5090, n64179, n3064, n49049, n3065, 
        n49048, n3066, n49047, n58490, n56565;
    wire [23:0]n8262;
    
    wire n2938, n49046, n2939, n49045, n2940, n49044, n2941, n49043, 
        n2942, n49042, n2943, n49041, n2944, n49040, n2945, n49039, 
        n2946, n49038, n2947, n49037, n2948, n49036, n2949, n49035, 
        n2950, n49034, n2951, n49033, n2952, n49032, n2953, n49031, 
        n2954, n49030, n2955, n49029, n2956, n49028, n2957, n49027, 
        n58488, n26_adj_5091, n28_adj_5092;
    wire [23:0]n8236;
    
    wire n2827, n49026, n2828, n49025, n2829, n49024, n24_adj_5093, 
        n35_adj_5094, n32, n2830, n49023, n2831, n49022, n2832, 
        n49021, n22_adj_5095, n64171, n65973, n37_adj_5096, n65974, 
        n39_adj_5097, n65864, n2833, n49020, n2834, n49019, n2835, 
        n49018, n2836, n49017, n2837, n49016, n65743, n20_adj_5098, 
        n63182, n65975, n2838, n49015, n2839, n49014, n2840, n49013, 
        n2841, n49012, n2842, n49011, n2843, n49010, n2844, n49009, 
        n49008, n58486;
    wire [23:0]n8210;
    
    wire n49007, n2714, n49006, n41_adj_5099, n64447, n2715, n49005, 
        n2716, n49004, n2717, n49003, n1699, n1700, n63316, n34_adj_5100, 
        n66136, n66137, n49002, n2719, n49001, n2720, n49000, 
        n48999, n48998, n1835, n39_adj_5101, n1836, n37_adj_5102, 
        n48997, n48996, n48995, n43_adj_5103, n66059, n1839, n31_adj_5104, 
        n63329, n48994, n1838, n33_adj_5105, n34_adj_5106, n1837, 
        n35_adj_5107, n48_adj_5108, n1834, n41_adj_5109, n63341, n1840, 
        n29_adj_5110, n63274, n48993, n36;
    wire [2:0]n479;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(34[17:28])
    
    wire n28373, n40_adj_5111, n48992, n48991, n48990, n32_adj_5112, 
        n40_adj_5113, n1841, n28_adj_5114, n65785, n56577, n48989, 
        n48988, n48987, n65786, n63270, n30_adj_5115, n63266, n65783, 
        n48986, n63357, n65551, n66094, n48985, n1832, n66095, 
        n48984, n1977, n58424, n58422, n59298, n1969, n1698, n1971, 
        n48814, n1967, n48813, n48812, n1697, n48811, n1970, n48810, 
        n48809, n1972, n48983, n25211, n48808, n1973, n48807, 
        n1974, n48806, n48982, n1975, n48805, n1976, n48804, n48803, 
        n48981, n41_adj_5116, n48980, n38_adj_5117, n48979, n48784, 
        n48783, n48978, n48782, n48977, n48781, n67140, n48780, 
        n48779, n48778, n48777, n48776, n43_adj_5118, n42_adj_5119, 
        n48775, n48774, n58474, n56602, n65797, n65798, n48976, 
        n48975, n48974, n48973, n58482, n56581, n65996, n36_adj_5120, 
        n48717, n1694, n48716, n48715, n1696, n48714, n48962, 
        n48713, n48961, n48712, n48711, n48710, n1701, n48709, 
        n1702, n48960, n38_adj_5121, n40_adj_5122, n48959, n48958, 
        n48957, n48956, n48955, n48954, n48953, n63348, n66103, 
        n66104, n59934, n45_adj_5123, n962, n31_adj_5124, n29_adj_5125, 
        n33_adj_5126, n35_adj_5127, n39_adj_5128, n37_adj_5129, n39_adj_5130, 
        n41_adj_5131, n37_adj_5132, n43_adj_5133, n31_adj_5134, n29_adj_5135, 
        n33_adj_5136, n35_adj_5137, n39_adj_5138, n58400, n38424, 
        n58748, n58766, n59896, n59966, n39_adj_5139, n41_adj_5140, 
        n961, n59936, n43_adj_5141, n34_adj_5142, n65795, n65796, 
        n64290, n38_adj_5143, n44_adj_5144, n65141, n48_adj_5145, 
        n59876, n59908, n59394, n59396, n28_adj_5146, n63229, n30_adj_5147, 
        n58586, n59212, n56622, n59190, n3_adj_5148, n59194, n58592, 
        n42_adj_5149, n5, n59198, n8, n65799, n65800, n63003, 
        n48_adj_5150, n63000, n62997, n58548, n58554, n59282, n25163, 
        n59854, n59960, n2, n10007, n44_adj_5151, n805, n39_adj_5152, 
        n41_adj_5153, n33_adj_5154, n43_adj_5155, n35_adj_5156, n37_adj_5157, 
        n29_adj_5158, n39_adj_5159, n31_adj_5160, n59270, n23_adj_5161, 
        n41_adj_5162, n25_adj_5163, n37_adj_5164, n7, n45_adj_5165, 
        n43_adj_5166, n9, n17_adj_5167, n19_adj_5168, n21_adj_5169, 
        n11, n13, n15, n27_adj_5170, n63681, n63701, n16_adj_5171, 
        n63653, n8_adj_5172, n24_adj_5173, n3274, n63722, n64688, 
        n32_adj_5174, n65793, n64680, n65794, n65895, n64282, n65229, 
        n14_adj_5175, n66066, n63927, n16_adj_5176, n12, n48_adj_5177, 
        n4_c, n65498, n18_adj_5178, n65499, n65143, n63888, n20_adj_5179, 
        n65541, n65791, n65792, n63671, n14_adj_5180, n15_adj_5181, 
        n55436, n10, n48_adj_5182, n28_adj_5183, n30_adj_5184, n63675, 
        n63246, n66005, n30_adj_5185, n64527, n66196, n66197, n6_adj_5186, 
        n65500, n65501, n63655, n65587, n64525, n66118, n63657, 
        n66054, n64533, n12_adj_5187, n63866, n14_adj_5188, n58436, 
        n3253, n66056, n59250, n58444, n16_adj_5190, n63834, n18_adj_5191, 
        n33_adj_5192, n31_adj_5193, n37_adj_5194, n35_adj_5195, n21_adj_5196, 
        n23_adj_5197, n9_adj_5198, n11_adj_5199, n19_adj_5200, n25_adj_5201, 
        n27_adj_5202, n10_adj_5203, n14_adj_5204, n13_adj_5205, n15_adj_5206, 
        n17_adj_5207, n63061, n63779, n16_adj_5208, n29_adj_5209, 
        n59398, n25214, n12_adj_5210, n63812, n63747, n64736, n65271, 
        n65267, n63749, n6_adj_5211, n65510, n14_adj_5212, n32_adj_5213, 
        n65511, n63741, n12_adj_5214, n63735, n66003, n64513, n8_adj_5215, 
        n65512, n65513, n63759, n64722, n62954, n62951, n10_adj_5216, 
        n65585, n64511, n65679, n66194, n65817, n66249, n66250, 
        n66240, n66043, n66044, n35_adj_5217, n39_adj_5218, n33_adj_5219, 
        n37_adj_5220, n27_adj_5221, n29_adj_5222, n23_adj_5223, n25_adj_5224, 
        n11_adj_5225, n59232, n13_adj_5226, n21_adj_5227, n15_adj_5228, 
        n17_adj_5229, n19_adj_5230, n31_adj_5231, n63795, n59230, 
        n64786, n65293, n65291, n59148, n63797, n8_adj_5232, n65518, 
        n65519, n46_adj_5233, n48_adj_5234, n59182, n34_adj_5235, 
        n25152, n63781, n65999, n64501, n65520, n65521, n64768, 
        n20_adj_5236, n64499, n65689, n66192, n65581, n66251, n66252, 
        n66242, n65758, n42_adj_5237, n65801, n65802, n48_adj_5238, 
        n66238, n40_adj_5239, n66246, n35_adj_5240, n37_adj_5241, 
        n41_adj_5242, n39_adj_5243, n29_adj_5244, n31_adj_5245, n23_adj_5246, 
        n25_adj_5247, n27_adj_5248, n13_adj_5249, n15_adj_5250, n17_adj_5251, 
        n19_adj_5252, n21_adj_5253, n33_adj_5254, n63845, n64827, 
        n65315, n65313, n63847, n10_adj_5255, n65548, n65549, n36_adj_5256, 
        n63837, n65997, n64489, n22_adj_5257, n65991, n65992, n65840, 
        n65697, n66190, n64487, n66247, n66248, n41_adj_5258, n39_adj_5259, 
        n37_adj_5260, n43_adj_5261, n41_adj_5262, n27_adj_5263, n63255, 
        n31_adj_5264, n33_adj_5265, n25_adj_5266, n27_adj_5267, n29_adj_5268, 
        n15_adj_5269, n17_adj_5270, n19_adj_5271, n21_adj_5272, n23_adj_5273, 
        n35_adj_5274, n63908, n64881, n65345, n65343, n63910, n12_adj_5275, 
        n65589, n38_adj_5276, n26_adj_5277, n65781, n65782, n38_adj_5278, 
        n65590, n63898, n63249, n65985, n66105, n65555, n66233, 
        n66234, n64481, n66189, n48_adj_5279, n24_adj_5280, n65983, 
        n65984, n65850, n65709, n66184, n59300, n64479, n66237, 
        n56605, n32_adj_5281, n65789, n65790, n64272, n65145, n65545, 
        n65787, n65788, n48_adj_5282, n59280, n25178, n27_adj_5283, 
        n63235, n38_adj_5284, n56596, n26_adj_5285, n65771;
    
    SB_LUT4 i48497_3_lut (.I0(n65772), .I1(baudrate[8]), .I2(n37), .I3(GND_net), 
            .O(n65559));   // verilog/uart_rx.v(119[33:55])
    defparam i48497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i27_2_lut (.I0(n2723), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n27_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i29_2_lut (.I0(n2722), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i31_2_lut (.I0(n2721), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1836_3_lut (.I0(n2610), .I1(n8184[9]), .I2(n294[6]), 
            .I3(GND_net), .O(n2727));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2752_7_lut (.I0(GND_net), .I1(n2487), .I2(n1460), .I3(n48951), 
            .O(n8158[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_7 (.CI(n48951), .I0(n2487), .I1(n1460), .CO(n48952));
    SB_LUT4 div_37_i1837_3_lut (.I0(n2611), .I1(n8184[8]), .I2(n294[6]), 
            .I3(GND_net), .O(n2728));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49173_4_lut (.I0(n65559), .I1(n66107), .I2(n41), .I3(n63231), 
            .O(n66235));   // verilog/uart_rx.v(119[33:55])
    defparam i49173_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_37_i1838_3_lut (.I0(n2612), .I1(n8184[7]), .I2(n294[6]), 
            .I3(GND_net), .O(n2729));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2752_6_lut (.I0(GND_net), .I1(n2488), .I2(n1011), .I3(n48950), 
            .O(n8158[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1845_i17_2_lut (.I0(n2728), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i19_2_lut (.I0(n2727), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1833_3_lut (.I0(n2607), .I1(n8184[12]), .I2(n294[6]), 
            .I3(GND_net), .O(n2724));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1833_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2752_6 (.CI(n48950), .I0(n2488), .I1(n1011), .CO(n48951));
    SB_LUT4 add_2752_5_lut (.I0(GND_net), .I1(n2489), .I2(n856), .I3(n48949), 
            .O(n8158[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1834_3_lut (.I0(n2608), .I1(n8184[11]), .I2(n294[6]), 
            .I3(GND_net), .O(n2725));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1834_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2752_5 (.CI(n48949), .I0(n2489), .I1(n856), .CO(n48950));
    SB_LUT4 div_37_i1835_3_lut (.I0(n2609), .I1(n8184[10]), .I2(n294[6]), 
            .I3(GND_net), .O(n2726));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1675_3_lut (.I0(n2366), .I1(n8132[10]), .I2(n294[8]), 
            .I3(GND_net), .O(n2489));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i21_2_lut (.I0(n2726), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i23_2_lut (.I0(n2725), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n23_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i25_2_lut (.I0(n2724), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2752_4_lut (.I0(GND_net), .I1(n2490), .I2(n698), .I3(n48948), 
            .O(n8158[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_4 (.CI(n48948), .I0(n2490), .I1(n698), .CO(n48949));
    SB_LUT4 add_2752_3_lut (.I0(GND_net), .I1(n2491), .I2(n858), .I3(n48947), 
            .O(n8158[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_3 (.CI(n48947), .I0(n2491), .I1(n858), .CO(n48948));
    SB_LUT4 div_37_LessThan_1845_i37_2_lut (.I0(n2718), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2752_2_lut (.I0(n56585), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n58480)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2752_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n48947));
    SB_LUT4 add_2751_17_lut (.I0(GND_net), .I1(n2353), .I2(n2638), .I3(n48946), 
            .O(n8132[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2751_16_lut (.I0(GND_net), .I1(n2354), .I2(n2519), .I3(n48945), 
            .O(n8132[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46901_4_lut (.I0(n37_adj_5013), .I1(n25), .I2(n23_c), .I3(n21), 
            .O(n63963));
    defparam i46901_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47887_4_lut (.I0(n19), .I1(n17), .I2(n2729), .I3(baudrate[2]), 
            .O(n64949));
    defparam i47887_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i48321_4_lut (.I0(n25), .I1(n23_c), .I2(n21), .I3(n64949), 
            .O(n65383));
    defparam i48321_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48313_4_lut (.I0(n31), .I1(n29_c), .I2(n27_c), .I3(n65383), 
            .O(n65375));
    defparam i48313_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY add_2751_16 (.CI(n48945), .I0(n2354), .I1(n2519), .CO(n48946));
    SB_LUT4 i46908_4_lut (.I0(n37_adj_5013), .I1(n35), .I2(n33), .I3(n65375), 
            .O(n63970));
    defparam i46908_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1845_i14_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2730), .I3(GND_net), .O(n14));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i14_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48533_3_lut (.I0(n14), .I1(baudrate[13]), .I2(n37_adj_5013), 
            .I3(GND_net), .O(n65595));   // verilog/uart_rx.v(119[33:55])
    defparam i48533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48534_3_lut (.I0(n65595), .I1(baudrate[14]), .I2(n39), .I3(GND_net), 
            .O(n65596));   // verilog/uart_rx.v(119[33:55])
    defparam i48534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49174_3_lut (.I0(n66235), .I1(baudrate[11]), .I2(n2100), 
            .I3(GND_net), .O(n66236));   // verilog/uart_rx.v(119[33:55])
    defparam i49174_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i40_3_lut (.I0(n22), .I1(baudrate[17]), 
            .I2(n45), .I3(GND_net), .O(n40));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46890_4_lut (.I0(n43), .I1(n41_adj_5014), .I2(n39), .I3(n63963), 
            .O(n63952));
    defparam i46890_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48513_4_lut (.I0(n40), .I1(n20), .I2(n45), .I3(n63950), 
            .O(n65575));   // verilog/uart_rx.v(119[33:55])
    defparam i48513_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47413_3_lut (.I0(n65596), .I1(baudrate[15]), .I2(n41_adj_5014), 
            .I3(GND_net), .O(n64475));   // verilog/uart_rx.v(119[33:55])
    defparam i47413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49125_3_lut (.I0(n66236), .I1(baudrate[12]), .I2(n2099), 
            .I3(GND_net), .O(n66187));   // verilog/uart_rx.v(119[33:55])
    defparam i49125_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49070_3_lut (.I0(n66187), .I1(baudrate[13]), .I2(n2098), 
            .I3(GND_net), .O(n48));   // verilog/uart_rx.v(119[33:55])
    defparam i49070_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i26_3_lut (.I0(n18), .I1(baudrate[9]), 
            .I2(n29_c), .I3(GND_net), .O(n26));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48919_4_lut (.I0(n26), .I1(n16), .I2(n29_c), .I3(n63997), 
            .O(n65981));   // verilog/uart_rx.v(119[33:55])
    defparam i48919_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut (.I0(baudrate[27]), .I1(baudrate[24]), .I2(baudrate[29]), 
            .I3(baudrate[30]), .O(n59304));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48920_3_lut (.I0(n65981), .I1(baudrate[10]), .I2(n31), .I3(GND_net), 
            .O(n65982));   // verilog/uart_rx.v(119[33:55])
    defparam i48920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48792_3_lut (.I0(n65982), .I1(baudrate[11]), .I2(n33), .I3(GND_net), 
            .O(n65854));   // verilog/uart_rx.v(119[33:55])
    defparam i48792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48655_4_lut (.I0(n43), .I1(n41_adj_5014), .I2(n39), .I3(n63970), 
            .O(n65717));
    defparam i48655_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2751_15_lut (.I0(GND_net), .I1(n2355), .I2(n2397), .I3(n48944), 
            .O(n8132[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_15 (.CI(n48944), .I0(n2355), .I1(n2397), .CO(n48945));
    SB_LUT4 add_2751_14_lut (.I0(GND_net), .I1(n2356), .I2(n2272), .I3(n48943), 
            .O(n8132[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_14 (.CI(n48943), .I0(n2356), .I1(n2272), .CO(n48944));
    SB_LUT4 i48989_4_lut (.I0(n64475), .I1(n65575), .I2(n45), .I3(n63952), 
            .O(n66051));   // verilog/uart_rx.v(119[33:55])
    defparam i48989_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47411_3_lut (.I0(n65854), .I1(baudrate[12]), .I2(n35), .I3(GND_net), 
            .O(n64473));   // verilog/uart_rx.v(119[33:55])
    defparam i47411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48991_4_lut (.I0(n64473), .I1(n66051), .I2(n45), .I3(n65717), 
            .O(n66053));   // verilog/uart_rx.v(119[33:55])
    defparam i48991_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_3_lut (.I0(n59254), .I1(n59302), .I2(n58984), .I3(GND_net), 
            .O(n59312));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_990 (.I0(n59312), .I1(n59308), .I2(n59310), .I3(n59304), 
            .O(n25187));
    defparam i1_4_lut_adj_990.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2751_13_lut (.I0(GND_net), .I1(n2357), .I2(n2144), .I3(n48942), 
            .O(n8132[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_13 (.CI(n48942), .I0(n2357), .I1(n2144), .CO(n48943));
    SB_LUT4 add_2751_12_lut (.I0(GND_net), .I1(n2358), .I2(n2013), .I3(n48941), 
            .O(n8132[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1743_3_lut (.I0(n2476), .I1(n8158[23]), .I2(n294[7]), 
            .I3(GND_net), .O(n2596));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4038_2_lut (.I0(n21311), .I1(n9620), .I2(GND_net), .I3(GND_net), 
            .O(n44));   // verilog/uart_rx.v(119[33:55])
    defparam i4038_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1754_3_lut (.I0(n2487), .I1(n8158[12]), .I2(n294[7]), 
            .I3(GND_net), .O(n2607));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(baudrate[14]), .I1(baudrate[15]), .I2(GND_net), 
            .I3(GND_net), .O(n59302));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1744_3_lut (.I0(n2477), .I1(n8158[22]), .I2(n294[7]), 
            .I3(GND_net), .O(n2597));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1748_3_lut (.I0(n2481), .I1(n8158[18]), .I2(n294[7]), 
            .I3(GND_net), .O(n2601));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2751_12 (.CI(n48941), .I0(n2358), .I1(n2013), .CO(n48942));
    SB_LUT4 add_2751_11_lut (.I0(GND_net), .I1(n2359), .I2(n1879), .I3(n48940), 
            .O(n8132[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_11 (.CI(n48940), .I0(n2359), .I1(n1879), .CO(n48941));
    SB_LUT4 div_37_LessThan_1766_i37_2_lut (.I0(n2601), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5015));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1745_3_lut (.I0(n2478), .I1(n8158[21]), .I2(n294[7]), 
            .I3(GND_net), .O(n2598));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2751_10_lut (.I0(GND_net), .I1(n2360), .I2(n1742), .I3(n48939), 
            .O(n8132[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_10 (.CI(n48939), .I0(n2360), .I1(n1742), .CO(n48940));
    SB_LUT4 div_37_LessThan_1766_i43_2_lut (.I0(n2598), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5016));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1747_3_lut (.I0(n2480), .I1(n8158[19]), .I2(n294[7]), 
            .I3(GND_net), .O(n2600));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i39_2_lut (.I0(n2600), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5017));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1746_3_lut (.I0(n2479), .I1(n8158[20]), .I2(n294[7]), 
            .I3(GND_net), .O(n2599));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2751_9_lut (.I0(GND_net), .I1(n2361), .I2(n1602), .I3(n48938), 
            .O(n8132[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_991 (.I0(baudrate[12]), .I1(baudrate[13]), .I2(GND_net), 
            .I3(GND_net), .O(n59226));
    defparam i1_2_lut_adj_991.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_992 (.I0(baudrate[10]), .I1(baudrate[11]), .I2(GND_net), 
            .I3(GND_net), .O(n59228));
    defparam i1_2_lut_adj_992.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_1766_i41_2_lut (.I0(n2599), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5018));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2751_9 (.CI(n48938), .I0(n2361), .I1(n1602), .CO(n48939));
    SB_LUT4 div_37_i1749_3_lut (.I0(n2482), .I1(n8158[17]), .I2(n294[7]), 
            .I3(GND_net), .O(n2602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2751_8_lut (.I0(GND_net), .I1(n2362), .I2(n1459), .I3(n48937), 
            .O(n8132[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i42772_2_lut (.I0(baudrate[21]), .I1(baudrate[22]), .I2(GND_net), 
            .I3(GND_net), .O(n59824));
    defparam i42772_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1751_3_lut (.I0(n2484), .I1(n8158[15]), .I2(n294[7]), 
            .I3(GND_net), .O(n2604));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1750_3_lut (.I0(n2483), .I1(n8158[16]), .I2(n294[7]), 
            .I3(GND_net), .O(n2603));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42901_4_lut (.I0(n59824), .I1(n59174), .I2(n59228), .I3(baudrate[9]), 
            .O(n59954));
    defparam i42901_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_993 (.I0(baudrate[23]), .I1(baudrate[28]), .I2(baudrate[27]), 
            .I3(baudrate[0]), .O(n58804));
    defparam i1_4_lut_adj_993.LUT_INIT = 16'h0100;
    SB_LUT4 div_37_LessThan_1766_i31_2_lut (.I0(n2604), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5019));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i33_2_lut (.I0(n2603), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5020));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i35_2_lut (.I0(n2602), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5021));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2751_8 (.CI(n48937), .I0(n2362), .I1(n1459), .CO(n48938));
    SB_LUT4 div_37_i1752_3_lut (.I0(n2485), .I1(n8158[14]), .I2(n294[7]), 
            .I3(GND_net), .O(n2605));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1753_3_lut (.I0(n2486), .I1(n8158[13]), .I2(n294[7]), 
            .I3(GND_net), .O(n2606));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42837_4_lut (.I0(baudrate[25]), .I1(baudrate[31]), .I2(baudrate[24]), 
            .I3(baudrate[29]), .O(n59890));
    defparam i42837_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i27_2_lut (.I0(n2606), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5022));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2751_7_lut (.I0(GND_net), .I1(n2363), .I2(n1460), .I3(n48936), 
            .O(n8132[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_7 (.CI(n48936), .I0(n2363), .I1(n1460), .CO(n48937));
    SB_LUT4 div_37_LessThan_1766_i29_2_lut (.I0(n2605), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5023));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1757_3_lut (.I0(n2490), .I1(n8158[9]), .I2(n294[7]), 
            .I3(GND_net), .O(n2610));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_994 (.I0(n56344), .I1(n58804), .I2(n59392), .I3(baudrate[16]), 
            .O(n58832));
    defparam i1_4_lut_adj_994.LUT_INIT = 16'h0004;
    SB_LUT4 div_37_i1756_3_lut (.I0(n2489), .I1(n8158[10]), .I2(n294[7]), 
            .I3(GND_net), .O(n2609));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2751_6_lut (.I0(GND_net), .I1(n2364), .I2(n1011), .I3(n48935), 
            .O(n8132[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1766_i19_2_lut (.I0(n2610), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5024));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i19_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2751_6 (.CI(n48935), .I0(n2364), .I1(n1011), .CO(n48936));
    SB_LUT4 div_37_LessThan_1766_i21_2_lut (.I0(n2609), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5025));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2751_5_lut (.I0(GND_net), .I1(n2365), .I2(n856), .I3(n48934), 
            .O(n8132[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2751_5 (.CI(n48934), .I0(n2365), .I1(n856), .CO(n48935));
    SB_LUT4 i42911_4_lut (.I0(n59890), .I1(n59886), .I2(n59888), .I3(n59810), 
            .O(n59964));
    defparam i42911_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1758_3_lut (.I0(n2491), .I1(n8158[8]), .I2(n294[7]), 
            .I3(GND_net), .O(n2611));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49219_4_lut (.I0(n59954), .I1(n63384), .I2(n59964), .I3(n58832), 
            .O(n66281));
    defparam i49219_4_lut.LUT_INIT = 16'hc9cc;
    SB_LUT4 div_37_i1755_3_lut (.I0(n2488), .I1(n8158[11]), .I2(n294[7]), 
            .I3(GND_net), .O(n2608));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1766_i23_2_lut (.I0(n2608), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5026));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i25_2_lut (.I0(n2607), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5027));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1766_i17_2_lut (.I0(n2611), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5028));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47029_4_lut (.I0(n23_adj_5026), .I1(n21_adj_5025), .I2(n19_adj_5024), 
            .I3(n17_adj_5028), .O(n64091));
    defparam i47029_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47016_4_lut (.I0(n29_adj_5023), .I1(n27_adj_5022), .I2(n25_adj_5027), 
            .I3(n64091), .O(n64078));
    defparam i47016_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48669_4_lut (.I0(n35_adj_5021), .I1(n33_adj_5020), .I2(n31_adj_5019), 
            .I3(n64078), .O(n65731));
    defparam i48669_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1766_i16_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2612), .I3(GND_net), .O(n16_adj_5029));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48543_3_lut (.I0(n16_adj_5029), .I1(baudrate[13]), .I2(n39_adj_5017), 
            .I3(GND_net), .O(n65605));   // verilog/uart_rx.v(119[33:55])
    defparam i48543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48544_3_lut (.I0(n65605), .I1(baudrate[14]), .I2(n41_adj_5018), 
            .I3(GND_net), .O(n65606));   // verilog/uart_rx.v(119[33:55])
    defparam i48544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47905_4_lut (.I0(n41_adj_5018), .I1(n39_adj_5017), .I2(n27_adj_5022), 
            .I3(n64087), .O(n64967));
    defparam i47905_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i48511_3_lut (.I0(n22_adj_5030), .I1(baudrate[7]), .I2(n27_adj_5022), 
            .I3(GND_net), .O(n65573));   // verilog/uart_rx.v(119[33:55])
    defparam i48511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47403_3_lut (.I0(n65606), .I1(baudrate[15]), .I2(n43_adj_5016), 
            .I3(GND_net), .O(n64465));   // verilog/uart_rx.v(119[33:55])
    defparam i47403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49227_2_lut (.I0(n48_adj_5031), .I1(n25229), .I2(GND_net), 
            .I3(GND_net), .O(n294[21]));
    defparam i49227_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_37_LessThan_1766_i28_3_lut (.I0(n20_adj_5032), .I1(baudrate[9]), 
            .I2(n31_adj_5019), .I3(GND_net), .O(n28));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_995 (.I0(n59238), .I1(n59302), .I2(baudrate[16]), 
            .I3(n38422), .O(n59096));
    defparam i1_4_lut_adj_995.LUT_INIT = 16'h0100;
    SB_LUT4 i48917_4_lut (.I0(n28), .I1(n18_adj_5033), .I2(n31_adj_5019), 
            .I3(n64068), .O(n65979));   // verilog/uart_rx.v(119[33:55])
    defparam i48917_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47112_3_lut (.I0(n57124), .I1(n57547), .I2(baudrate[2]), 
            .I3(GND_net), .O(n62993));   // verilog/uart_rx.v(119[33:55])
    defparam i47112_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i48918_3_lut (.I0(n65979), .I1(baudrate[10]), .I2(n33_adj_5020), 
            .I3(GND_net), .O(n65980));   // verilog/uart_rx.v(119[33:55])
    defparam i48918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2751_4_lut (.I0(GND_net), .I1(n2366), .I2(n698), .I3(n48933), 
            .O(n8132[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46930_4_lut (.I0(n56344), .I1(n59096), .I2(n59240), .I3(n59170), 
            .O(n62994));   // verilog/uart_rx.v(119[33:55])
    defparam i46930_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i48794_3_lut (.I0(n65980), .I1(baudrate[11]), .I2(n35_adj_5021), 
            .I3(GND_net), .O(n65856));   // verilog/uart_rx.v(119[33:55])
    defparam i48794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47909_4_lut (.I0(n41_adj_5018), .I1(n39_adj_5017), .I2(n37_adj_5015), 
            .I3(n65731), .O(n64971));
    defparam i47909_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i48541_4_lut (.I0(n64465), .I1(n65573), .I2(n43_adj_5016), 
            .I3(n64967), .O(n65603));   // verilog/uart_rx.v(119[33:55])
    defparam i48541_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i427_4_lut (.I0(n62994), .I1(n62993), .I2(n294[21]), 
            .I3(n59692), .O(n56317));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i427_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i47401_3_lut (.I0(n65856), .I1(baudrate[12]), .I2(n37_adj_5015), 
            .I3(GND_net), .O(n64463));   // verilog/uart_rx.v(119[33:55])
    defparam i47401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49076_4_lut (.I0(n64463), .I1(n65603), .I2(n43_adj_5016), 
            .I3(n64971), .O(n66138));   // verilog/uart_rx.v(119[33:55])
    defparam i49076_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_2751_4 (.CI(n48933), .I0(n2366), .I1(n698), .CO(n48934));
    SB_LUT4 add_2751_3_lut (.I0(GND_net), .I1(n2367), .I2(n858), .I3(n48932), 
            .O(n8132[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i534_3_lut (.I0(n56317), .I1(n294[20]), .I2(baudrate[3]), 
            .I3(GND_net), .O(n56321));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i534_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i49077_3_lut (.I0(n66138), .I1(baudrate[16]), .I2(n2597), 
            .I3(GND_net), .O(n66139));   // verilog/uart_rx.v(119[33:55])
    defparam i49077_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1662_3_lut (.I0(n2353), .I1(n8132[23]), .I2(n294[8]), 
            .I3(GND_net), .O(n2476));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39559_1_lut (.I0(n25205), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56573));
    defparam i39559_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1672_3_lut (.I0(n2363), .I1(n8132[13]), .I2(n294[8]), 
            .I3(GND_net), .O(n2486));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5808_4_lut (.I0(n804), .I1(n38422), .I2(n21309), .I3(baudrate[2]), 
            .O(n21311));   // verilog/uart_rx.v(119[33:55])
    defparam i5808_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 div_37_i1666_3_lut (.I0(n2357), .I1(n8132[19]), .I2(n294[8]), 
            .I3(GND_net), .O(n2480));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i39_2_lut (.I0(n2480), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5034));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1663_3_lut (.I0(n2354), .I1(n8132[22]), .I2(n294[8]), 
            .I3(GND_net), .O(n2477));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i45_2_lut (.I0(n2477), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5035));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1664_3_lut (.I0(n2355), .I1(n8132[21]), .I2(n294[8]), 
            .I3(GND_net), .O(n2478));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i43_2_lut (.I0(n2478), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5036));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1665_3_lut (.I0(n2356), .I1(n8132[20]), .I2(n294[8]), 
            .I3(GND_net), .O(n2479));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i41_2_lut (.I0(n2479), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5037));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1667_3_lut (.I0(n2358), .I1(n8132[18]), .I2(n294[8]), 
            .I3(GND_net), .O(n2481));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1669_3_lut (.I0(n2360), .I1(n8132[16]), .I2(n294[8]), 
            .I3(GND_net), .O(n2483));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1668_3_lut (.I0(n2359), .I1(n8132[17]), .I2(n294[8]), 
            .I3(GND_net), .O(n2482));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i33_2_lut (.I0(n2483), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5038));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i35_2_lut (.I0(n2482), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5039));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i37_2_lut (.I0(n2481), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5040));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1670_3_lut (.I0(n2361), .I1(n8132[15]), .I2(n294[8]), 
            .I3(GND_net), .O(n2484));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1671_3_lut (.I0(n2362), .I1(n8132[14]), .I2(n294[8]), 
            .I3(GND_net), .O(n2485));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1685_i29_2_lut (.I0(n2485), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5041));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i31_2_lut (.I0(n2484), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5042));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i21_2_lut (.I0(n2489), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5043));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i23_2_lut (.I0(n2488), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5044));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i25_2_lut (.I0(n2487), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5045));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1685_i27_2_lut (.I0(n2486), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i27_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2751_3 (.CI(n48932), .I0(n2367), .I1(n858), .CO(n48933));
    SB_LUT4 add_2751_2_lut (.I0(n56589), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n58478)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2751_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_37_LessThan_1685_i19_2_lut (.I0(n2490), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47075_4_lut (.I0(n25_adj_5045), .I1(n23_adj_5044), .I2(n21_adj_5043), 
            .I3(n19_adj_5047), .O(n64137));
    defparam i47075_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47071_4_lut (.I0(n31_adj_5042), .I1(n29_adj_5041), .I2(n27_adj_5046), 
            .I3(n64137), .O(n64133));
    defparam i47071_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48677_4_lut (.I0(n37_adj_5040), .I1(n35_adj_5039), .I2(n33_adj_5038), 
            .I3(n64133), .O(n65739));
    defparam i48677_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_2751_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n48932));
    SB_LUT4 i48547_3_lut (.I0(n18_adj_5048), .I1(baudrate[13]), .I2(n41_adj_5037), 
            .I3(GND_net), .O(n65609));   // verilog/uart_rx.v(119[33:55])
    defparam i48547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2750_16_lut (.I0(GND_net), .I1(n2227), .I2(n2519), .I3(n48931), 
            .O(n8106[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48548_3_lut (.I0(n65609), .I1(baudrate[14]), .I2(n43_adj_5036), 
            .I3(GND_net), .O(n65610));   // verilog/uart_rx.v(119[33:55])
    defparam i48548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47943_4_lut (.I0(n43_adj_5036), .I1(n41_adj_5037), .I2(n29_adj_5041), 
            .I3(n64135), .O(n65005));
    defparam i47943_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_LessThan_1685_i26_3_lut (.I0(n24), .I1(baudrate[7]), 
            .I2(n29_adj_5041), .I3(GND_net), .O(n26_adj_5049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47397_3_lut (.I0(n65610), .I1(baudrate[15]), .I2(n45_adj_5035), 
            .I3(GND_net), .O(n64459));   // verilog/uart_rx.v(119[33:55])
    defparam i47397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2750_15_lut (.I0(GND_net), .I1(n2228), .I2(n2397), .I3(n48930), 
            .O(n8106[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1685_i30_3_lut (.I0(n22_adj_5050), .I1(baudrate[9]), 
            .I2(n33_adj_5038), .I3(GND_net), .O(n30));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48915_4_lut (.I0(n30), .I1(n20_adj_5051), .I2(n33_adj_5038), 
            .I3(n64125), .O(n65977));   // verilog/uart_rx.v(119[33:55])
    defparam i48915_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48916_3_lut (.I0(n65977), .I1(baudrate[10]), .I2(n35_adj_5039), 
            .I3(GND_net), .O(n65978));   // verilog/uart_rx.v(119[33:55])
    defparam i48916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48796_3_lut (.I0(n65978), .I1(baudrate[11]), .I2(n37_adj_5040), 
            .I3(GND_net), .O(n65858));   // verilog/uart_rx.v(119[33:55])
    defparam i48796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i535_4_lut (.I0(n66281), .I1(n44_adj_5052), .I2(n294[20]), 
            .I3(baudrate[2]), .O(n803));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i535_4_lut.LUT_INIT = 16'h9565;
    SB_LUT4 i47945_4_lut (.I0(n43_adj_5036), .I1(n41_adj_5037), .I2(n39_adj_5034), 
            .I3(n65739), .O(n65007));
    defparam i47945_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i48508_4_lut (.I0(n64459), .I1(n26_adj_5049), .I2(n45_adj_5035), 
            .I3(n65005), .O(n65570));   // verilog/uart_rx.v(119[33:55])
    defparam i48508_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47395_3_lut (.I0(n65858), .I1(baudrate[12]), .I2(n39_adj_5034), 
            .I3(GND_net), .O(n64457));   // verilog/uart_rx.v(119[33:55])
    defparam i47395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48510_4_lut (.I0(n64457), .I1(n65570), .I2(n45_adj_5035), 
            .I3(n65007), .O(n65572));   // verilog/uart_rx.v(119[33:55])
    defparam i48510_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i4045_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n9620), .I3(n21311), 
            .O(n46));   // verilog/uart_rx.v(119[33:55])
    defparam i4045_4_lut.LUT_INIT = 16'hbbb2;
    SB_LUT4 div_37_i639_4_lut (.I0(n56321), .I1(n294[19]), .I2(n46), .I3(baudrate[4]), 
            .O(n56323));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i639_4_lut.LUT_INIT = 16'h6aa6;
    SB_CARRY add_2750_15 (.CI(n48930), .I0(n2228), .I1(n2397), .CO(n48931));
    SB_LUT4 add_2745_11_lut (.I0(GND_net), .I1(n1552), .I2(n1879), .I3(n48662), 
            .O(n7976[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5819_4_lut (.I0(n960), .I1(n9784), .I2(n21323), .I3(baudrate[3]), 
            .O(n21325));   // verilog/uart_rx.v(119[33:55])
    defparam i5819_4_lut.LUT_INIT = 16'ha8aa;
    SB_LUT4 add_2750_14_lut (.I0(GND_net), .I1(n2229), .I2(n2272), .I3(n48929), 
            .O(n8106[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_14 (.CI(n48929), .I0(n2229), .I1(n2272), .CO(n48930));
    SB_LUT4 add_2745_10_lut (.I0(GND_net), .I1(n1553), .I2(n1742), .I3(n48661), 
            .O(n7976[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2750_13_lut (.I0(GND_net), .I1(n2230), .I2(n2144), .I3(n48928), 
            .O(n8106[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_13 (.CI(n48928), .I0(n2230), .I1(n2144), .CO(n48929));
    SB_CARRY add_2745_10 (.CI(n48661), .I0(n1553), .I1(n1742), .CO(n48662));
    SB_LUT4 add_2750_12_lut (.I0(GND_net), .I1(n2231), .I2(n2013), .I3(n48927), 
            .O(n8106[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_12 (.CI(n48927), .I0(n2231), .I1(n2013), .CO(n48928));
    SB_LUT4 add_2745_9_lut (.I0(GND_net), .I1(n1554), .I2(n1602), .I3(n48660), 
            .O(n7976[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2745_9 (.CI(n48660), .I0(n1554), .I1(n1602), .CO(n48661));
    SB_LUT4 add_2750_11_lut (.I0(GND_net), .I1(n2232), .I2(n1879), .I3(n48926), 
            .O(n8106[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2745_8_lut (.I0(GND_net), .I1(n1555), .I2(n1459), .I3(n48659), 
            .O(n7976[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_11 (.CI(n48926), .I0(n2232), .I1(n1879), .CO(n48927));
    SB_LUT4 add_2750_10_lut (.I0(GND_net), .I1(n2233), .I2(n1742), .I3(n48925), 
            .O(n8106[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_10 (.CI(n48925), .I0(n2233), .I1(n1742), .CO(n48926));
    SB_LUT4 add_2750_9_lut (.I0(GND_net), .I1(n2234), .I2(n1602), .I3(n48924), 
            .O(n8106[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i640_4_lut (.I0(n803), .I1(baudrate[3]), .I2(n294[19]), 
            .I3(n44), .O(n959));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i640_4_lut.LUT_INIT = 16'h6a9a;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk16MHz), .D(n3), .R(r_SM_Main[2]));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Data_56 (.Q(r_Rx_Data), .C(clk16MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(42[10] 46[8])
    SB_CARRY add_2750_9 (.CI(n48924), .I0(n2234), .I1(n1602), .CO(n48925));
    SB_LUT4 add_2750_8_lut (.I0(GND_net), .I1(n2235), .I2(n1459), .I3(n48923), 
            .O(n8106[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Data_R_55 (.Q(r_Rx_Data_R), .C(clk16MHz), .D(RX_N_2));   // verilog/uart_rx.v(42[10] 46[8])
    SB_CARRY add_2745_8 (.CI(n48659), .I0(n1555), .I1(n1459), .CO(n48660));
    SB_CARRY add_2750_8 (.CI(n48923), .I0(n2235), .I1(n1459), .CO(n48924));
    SB_LUT4 i4216_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n9791), .I3(n21325), 
            .O(n46_adj_5053));   // verilog/uart_rx.v(119[33:55])
    defparam i4216_4_lut.LUT_INIT = 16'hbbb2;
    SB_LUT4 add_2750_7_lut (.I0(GND_net), .I1(n2236), .I2(n1460), .I3(n48922), 
            .O(n8106[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i742_4_lut (.I0(n56323), .I1(n294[18]), .I2(n46_adj_5053), 
            .I3(baudrate[5]), .O(n1111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i742_4_lut.LUT_INIT = 16'h9559;
    SB_LUT4 add_2745_7_lut (.I0(GND_net), .I1(n1556), .I2(n1460), .I3(n48658), 
            .O(n7976[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_7 (.CI(n48922), .I0(n2236), .I1(n1460), .CO(n48923));
    SB_LUT4 add_2750_6_lut (.I0(GND_net), .I1(n2237), .I2(n1011), .I3(n48921), 
            .O(n8106[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2750_6 (.CI(n48921), .I0(n2237), .I1(n1011), .CO(n48922));
    SB_CARRY add_2745_7 (.CI(n48658), .I0(n1556), .I1(n1460), .CO(n48659));
    SB_LUT4 add_2750_5_lut (.I0(GND_net), .I1(n2238), .I2(n856), .I3(n48920), 
            .O(n8106[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2745_6_lut (.I0(GND_net), .I1(n1557), .I2(n1011), .I3(n48657), 
            .O(n7976[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2745_6 (.CI(n48657), .I0(n1557), .I1(n1011), .CO(n48658));
    SB_CARRY add_2750_5 (.CI(n48920), .I0(n2238), .I1(n856), .CO(n48921));
    SB_LUT4 add_2745_5_lut (.I0(GND_net), .I1(n1558), .I2(n856), .I3(n48656), 
            .O(n7976[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2745_5 (.CI(n48656), .I0(n1558), .I1(n856), .CO(n48657));
    SB_LUT4 i42894_1_lut (.I0(n59946), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56569));
    defparam i42894_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2750_4_lut (.I0(GND_net), .I1(n2239), .I2(n698), .I3(n48919), 
            .O(n8106[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2745_4_lut (.I0(GND_net), .I1(n1559), .I2(n698), .I3(n48655), 
            .O(n7976[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2745_4 (.CI(n48655), .I0(n1559), .I1(n698), .CO(n48656));
    SB_CARRY add_2750_4 (.CI(n48919), .I0(n2239), .I1(n698), .CO(n48920));
    SB_LUT4 add_2750_3_lut (.I0(GND_net), .I1(n2240), .I2(n858), .I3(n48918), 
            .O(n8106[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2745_3_lut (.I0(GND_net), .I1(n1560), .I2(n858), .I3(n48654), 
            .O(n7976[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2745_3 (.CI(n48654), .I0(n1560), .I1(n858), .CO(n48655));
    SB_LUT4 add_2745_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n7976[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2745_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2745_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n48654));
    SB_CARRY add_2750_3 (.CI(n48918), .I0(n2240), .I1(n858), .CO(n48919));
    SB_LUT4 add_2750_2_lut (.I0(n56593), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n58476)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2750_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2750_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n48918));
    SB_LUT4 div_37_i843_3_lut (.I0(n1111), .I1(n7898[23]), .I2(n294[17]), 
            .I3(GND_net), .O(n1261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i942_3_lut (.I0(n1261), .I1(n7924[23]), .I2(n294[16]), 
            .I3(GND_net), .O(n1408));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1039_3_lut (.I0(n1408), .I1(n7950[23]), .I2(n294[15]), 
            .I3(GND_net), .O(n1552));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1134_3_lut (.I0(n1552), .I1(n7976[23]), .I2(n294[14]), 
            .I3(GND_net), .O(n1693));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1227_3_lut (.I0(n1693), .I1(n8002[23]), .I2(n294[13]), 
            .I3(GND_net), .O(n1831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1318_3_lut (.I0(n1831), .I1(n8028[23]), .I2(n294[12]), 
            .I3(GND_net), .O(n1966));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_Clock_Count_2053_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n49243), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2053_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n49242), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1407_3_lut (.I0(n1966), .I1(n8054[23]), .I2(n294[11]), 
            .I3(GND_net), .O(n2098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1407_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY r_Clock_Count_2053_add_4_8 (.CI(n49242), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n49243));
    SB_LUT4 r_Clock_Count_2053_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n49241), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_7 (.CI(n49241), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n49242));
    SB_LUT4 r_Clock_Count_2053_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n49240), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_6 (.CI(n49240), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n49241));
    SB_LUT4 r_Clock_Count_2053_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n49239), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_5 (.CI(n49239), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n49240));
    SB_LUT4 r_Clock_Count_2053_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n49238), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_4 (.CI(n49238), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n49239));
    SB_LUT4 r_Clock_Count_2053_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n49237), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_3 (.CI(n49237), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n49238));
    SB_LUT4 r_Clock_Count_2053_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2053_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2053_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n49237));
    SB_LUT4 div_37_i1494_3_lut (.I0(n2098), .I1(n8080[23]), .I2(n294[10]), 
            .I3(GND_net), .O(n2227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_996 (.I0(baudrate[29]), .I1(baudrate[24]), .I2(GND_net), 
            .I3(GND_net), .O(n59252));
    defparam i1_2_lut_adj_996.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_997 (.I0(baudrate[20]), .I1(baudrate[21]), .I2(GND_net), 
            .I3(GND_net), .O(n59296));
    defparam i1_2_lut_adj_997.LUT_INIT = 16'heeee;
    SB_LUT4 sub_38_add_2_26_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n48406), .O(\o_Rx_DV_N_3488[24] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_25_lut (.I0(n58448), .I1(n25108), .I2(VCC_net), 
            .I3(n48405), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_25 (.CI(n48405), .I0(n25108), .I1(VCC_net), 
            .CO(n48406));
    SB_LUT4 i1_2_lut_adj_998 (.I0(baudrate[31]), .I1(baudrate[26]), .I2(GND_net), 
            .I3(GND_net), .O(n59254));
    defparam i1_2_lut_adj_998.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_999 (.I0(n59294), .I1(n59202), .I2(n58984), .I3(baudrate[19]), 
            .O(n59004));
    defparam i1_4_lut_adj_999.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_38_add_2_24_lut (.I0(n58524), .I1(n59974), .I2(VCC_net), 
            .I3(n48404), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i1_4_lut_adj_1000 (.I0(n59004), .I1(n59254), .I2(n59296), 
            .I3(n59252), .O(n25202));
    defparam i1_4_lut_adj_1000.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_341_i48_3_lut (.I0(n57124), .I1(baudrate[2]), 
            .I2(n57547), .I3(GND_net), .O(n48_adj_5031));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_341_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_4_lut_adj_1001 (.I0(n59012), .I1(n59008), .I2(n59010), 
            .I3(n59810), .O(n59030));
    defparam i1_4_lut_adj_1001.LUT_INIT = 16'hfffe;
    SB_CARRY sub_38_add_2_24 (.CI(n48404), .I0(n59974), .I1(VCC_net), 
            .CO(n48405));
    SB_LUT4 i1_4_lut_adj_1002 (.I0(n59020), .I1(n59016), .I2(n59018), 
            .I3(n59014), .O(n59032));
    defparam i1_4_lut_adj_1002.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_38_add_2_23_lut (.I0(o_Rx_DV_N_3488[18]), .I1(n294[21]), 
            .I2(VCC_net), .I3(n48403), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_23 (.CI(n48403), .I0(n294[21]), .I1(VCC_net), 
            .CO(n48404));
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk16MHz), .D(n3_adj_5063), 
            .R(r_SM_Main[2]));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 i1_3_lut_adj_1003 (.I0(n59032), .I1(n25202), .I2(n59030), 
            .I3(GND_net), .O(n25229));
    defparam i1_3_lut_adj_1003.LUT_INIT = 16'hfefe;
    SB_LUT4 i46800_4_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n5225), .I3(\o_Rx_DV_N_3488[8] ), .O(n63088));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i46800_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 sub_38_add_2_22_lut (.I0(n58522), .I1(n294[20]), .I2(VCC_net), 
            .I3(n48402), .O(n58524)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_22 (.CI(n48402), .I0(n294[20]), .I1(VCC_net), 
            .CO(n48403));
    SB_LUT4 i46934_4_lut (.I0(r_Rx_Data), .I1(\o_Rx_DV_N_3488[12] ), .I2(n55210), 
            .I3(r_SM_Main[0]), .O(n63094));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i46934_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i46797_4_lut (.I0(n63088), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n63085));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i46797_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i46803_4_lut (.I0(n63094), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n63091));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i46803_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_1_i3_4_lut (.I0(n63091), .I1(n63085), 
            .I2(r_SM_Main[1]), .I3(n27), .O(n3_adj_5063));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_1_i3_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 sub_38_add_2_21_lut (.I0(n58520), .I1(n294[19]), .I2(VCC_net), 
            .I3(n48401), .O(n58522)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_21 (.CI(n48401), .I0(n294[19]), .I1(VCC_net), 
            .CO(n48402));
    SB_LUT4 sub_38_add_2_20_lut (.I0(GND_net), .I1(n294[18]), .I2(VCC_net), 
            .I3(n48400), .O(o_Rx_DV_N_3488[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_20 (.CI(n48400), .I0(n294[18]), .I1(VCC_net), 
            .CO(n48401));
    SB_LUT4 sub_38_add_2_19_lut (.I0(n58518), .I1(n294[17]), .I2(VCC_net), 
            .I3(n48399), .O(n58520)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_19 (.CI(n48399), .I0(n294[17]), .I1(VCC_net), 
            .CO(n48400));
    SB_LUT4 i46328_2_lut (.I0(baudrate[1]), .I1(n294[20]), .I2(GND_net), 
            .I3(GND_net), .O(n63390));   // verilog/uart_rx.v(119[33:55])
    defparam i46328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47012_4_lut (.I0(n25229), .I1(n63390), .I2(n48_adj_5031), 
            .I3(baudrate[0]), .O(n804));
    defparam i47012_4_lut.LUT_INIT = 16'h3633;
    SB_LUT4 div_37_i641_4_lut (.I0(n804), .I1(n42_adj_5064), .I2(n294[19]), 
            .I3(baudrate[2]), .O(n960));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i641_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 sub_38_add_2_18_lut (.I0(n58516), .I1(n294[16]), .I2(VCC_net), 
            .I3(n48398), .O(n58518)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_18 (.CI(n48398), .I0(n294[16]), .I1(VCC_net), 
            .CO(n48399));
    SB_LUT4 add_2744_10_lut (.I0(GND_net), .I1(n1408), .I2(n1742), .I3(n48626), 
            .O(n7950[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_17_lut (.I0(n58446), .I1(n294[15]), .I2(VCC_net), 
            .I3(n48397), .O(n58448)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_17 (.CI(n48397), .I0(n294[15]), .I1(VCC_net), 
            .CO(n48398));
    SB_LUT4 add_2744_9_lut (.I0(GND_net), .I1(n1409), .I2(n1602), .I3(n48625), 
            .O(n7950[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2744_9 (.CI(n48625), .I0(n1409), .I1(n1602), .CO(n48626));
    SB_LUT4 add_2744_8_lut (.I0(GND_net), .I1(n1410), .I2(n1459), .I3(n48624), 
            .O(n7950[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_16_lut (.I0(n58514), .I1(n294[14]), .I2(VCC_net), 
            .I3(n48396), .O(n58516)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_16 (.CI(n48396), .I0(n294[14]), .I1(VCC_net), 
            .CO(n48397));
    SB_LUT4 sub_38_add_2_15_lut (.I0(o_Rx_DV_N_3488[10]), .I1(n294[13]), 
            .I2(VCC_net), .I3(n48395), .O(n58514)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_2744_8 (.CI(n48624), .I0(n1410), .I1(n1459), .CO(n48625));
    SB_LUT4 add_2744_7_lut (.I0(GND_net), .I1(n1411), .I2(n1460), .I3(n48623), 
            .O(n7950[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_15 (.CI(n48395), .I0(n294[13]), .I1(VCC_net), 
            .CO(n48396));
    SB_LUT4 add_2749_14_lut (.I0(GND_net), .I1(n2098), .I2(n2397), .I3(n48895), 
            .O(n8080[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2744_7 (.CI(n48623), .I0(n1411), .I1(n1460), .CO(n48624));
    SB_LUT4 sub_38_add_2_14_lut (.I0(GND_net), .I1(n294[12]), .I2(VCC_net), 
            .I3(n48394), .O(\o_Rx_DV_N_3488[12] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i744_4_lut (.I0(n960), .I1(baudrate[3]), .I2(n294[18]), 
            .I3(n42_adj_5065), .O(n1113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i744_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 add_2749_13_lut (.I0(GND_net), .I1(n2099), .I2(n2272), .I3(n48894), 
            .O(n8080[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2744_6_lut (.I0(GND_net), .I1(n1412), .I2(n1011), .I3(n48622), 
            .O(n7950[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_13 (.CI(n48894), .I0(n2099), .I1(n2272), .CO(n48895));
    SB_CARRY add_2744_6 (.CI(n48622), .I0(n1412), .I1(n1011), .CO(n48623));
    SB_CARRY sub_38_add_2_14 (.CI(n48394), .I0(n294[12]), .I1(VCC_net), 
            .CO(n48395));
    SB_LUT4 add_2744_5_lut (.I0(GND_net), .I1(n1413), .I2(n856), .I3(n48621), 
            .O(n7950[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_13_lut (.I0(o_Rx_DV_N_3488[9]), .I1(n294[11]), 
            .I2(VCC_net), .I3(n48393), .O(n58446)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_13_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_38_add_2_13 (.CI(n48393), .I0(n294[11]), .I1(VCC_net), 
            .CO(n48394));
    SB_LUT4 i1_2_lut_adj_1004 (.I0(baudrate[15]), .I1(baudrate[16]), .I2(GND_net), 
            .I3(GND_net), .O(n59008));
    defparam i1_2_lut_adj_1004.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1005 (.I0(baudrate[11]), .I1(baudrate[12]), .I2(GND_net), 
            .I3(GND_net), .O(n59012));
    defparam i1_2_lut_adj_1005.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1006 (.I0(baudrate[9]), .I1(baudrate[10]), .I2(GND_net), 
            .I3(GND_net), .O(n59014));
    defparam i1_2_lut_adj_1006.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1007 (.I0(baudrate[7]), .I1(baudrate[8]), .I2(GND_net), 
            .I3(GND_net), .O(n59016));
    defparam i1_2_lut_adj_1007.LUT_INIT = 16'heeee;
    SB_LUT4 add_2749_12_lut (.I0(GND_net), .I1(n2100), .I2(n2144), .I3(n48893), 
            .O(n8080[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_12_lut (.I0(GND_net), .I1(n294[10]), .I2(VCC_net), 
            .I3(n48392), .O(o_Rx_DV_N_3488[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2744_5 (.CI(n48621), .I0(n1413), .I1(n856), .CO(n48622));
    SB_CARRY add_2749_12 (.CI(n48893), .I0(n2100), .I1(n2144), .CO(n48894));
    SB_LUT4 add_2744_4_lut (.I0(GND_net), .I1(n1414), .I2(n698), .I3(n48620), 
            .O(n7950[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2744_4 (.CI(n48620), .I0(n1414), .I1(n698), .CO(n48621));
    SB_LUT4 i39337_2_lut (.I0(baudrate[2]), .I1(baudrate[3]), .I2(GND_net), 
            .I3(GND_net), .O(n56344));
    defparam i39337_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY sub_38_add_2_12 (.CI(n48392), .I0(n294[10]), .I1(VCC_net), 
            .CO(n48393));
    SB_LUT4 sub_38_add_2_11_lut (.I0(GND_net), .I1(n294[9]), .I2(VCC_net), 
            .I3(n48391), .O(o_Rx_DV_N_3488[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2749_11_lut (.I0(GND_net), .I1(n2101), .I2(n2013), .I3(n48892), 
            .O(n8080[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2744_3_lut (.I0(GND_net), .I1(n1415), .I2(n858), .I3(n48619), 
            .O(n7950[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_11 (.CI(n48391), .I0(n294[9]), .I1(VCC_net), 
            .CO(n48392));
    SB_CARRY add_2744_3 (.CI(n48619), .I0(n1415), .I1(n858), .CO(n48620));
    SB_LUT4 add_2744_2_lut (.I0(n56611), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n58472)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2744_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_38_add_2_10_lut (.I0(GND_net), .I1(n294[8]), .I2(VCC_net), 
            .I3(n48390), .O(\o_Rx_DV_N_3488[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_10 (.CI(n48390), .I0(n294[8]), .I1(VCC_net), 
            .CO(n48391));
    SB_LUT4 sub_38_add_2_9_lut (.I0(GND_net), .I1(n294[7]), .I2(VCC_net), 
            .I3(n48389), .O(\o_Rx_DV_N_3488[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2744_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n48619));
    SB_CARRY add_2749_11 (.CI(n48892), .I0(n2101), .I1(n2013), .CO(n48893));
    SB_LUT4 i42821_3_lut (.I0(baudrate[31]), .I1(baudrate[21]), .I2(baudrate[27]), 
            .I3(GND_net), .O(n59874));
    defparam i42821_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 add_2749_10_lut (.I0(GND_net), .I1(n2102), .I2(n1879), .I3(n48891), 
            .O(n8080[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2743_9_lut (.I0(GND_net), .I1(n1261), .I2(n1602), .I3(n48618), 
            .O(n7924[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2743_8_lut (.I0(GND_net), .I1(n1262), .I2(n1459), .I3(n48617), 
            .O(n7924[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_9 (.CI(n48389), .I0(n294[7]), .I1(VCC_net), 
            .CO(n48390));
    SB_LUT4 sub_38_add_2_8_lut (.I0(GND_net), .I1(n294[6]), .I2(VCC_net), 
            .I3(n48388), .O(\o_Rx_DV_N_3488[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_8 (.CI(n48388), .I0(n294[6]), .I1(VCC_net), 
            .CO(n48389));
    SB_CARRY add_2743_8 (.CI(n48617), .I0(n1262), .I1(n1459), .CO(n48618));
    SB_CARRY add_2749_10 (.CI(n48891), .I0(n2102), .I1(n1879), .CO(n48892));
    SB_LUT4 sub_38_add_2_7_lut (.I0(GND_net), .I1(n294[5]), .I2(VCC_net), 
            .I3(n48387), .O(\o_Rx_DV_N_3488[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2743_7_lut (.I0(GND_net), .I1(n1263), .I2(n1460), .I3(n48616), 
            .O(n7924[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2749_9_lut (.I0(GND_net), .I1(n2103), .I2(n1742), .I3(n48890), 
            .O(n8080[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2743_7 (.CI(n48616), .I0(n1263), .I1(n1460), .CO(n48617));
    SB_CARRY sub_38_add_2_7 (.CI(n48387), .I0(n294[5]), .I1(VCC_net), 
            .CO(n48388));
    SB_LUT4 sub_38_add_2_6_lut (.I0(GND_net), .I1(n294[4]), .I2(VCC_net), 
            .I3(n48386), .O(\o_Rx_DV_N_3488[4] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_9 (.CI(n48890), .I0(n2103), .I1(n1742), .CO(n48891));
    SB_LUT4 div_37_i845_3_lut (.I0(n1113), .I1(n7898[21]), .I2(n294[17]), 
            .I3(GND_net), .O(n1263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42893_4_lut (.I0(n59874), .I1(n59294), .I2(n59872), .I3(n59248), 
            .O(n59946));
    defparam i42893_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2743_6_lut (.I0(GND_net), .I1(n1264), .I2(n1011), .I3(n48615), 
            .O(n7924[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2743_6 (.CI(n48615), .I0(n1264), .I1(n1011), .CO(n48616));
    SB_CARRY sub_38_add_2_6 (.CI(n48386), .I0(n294[4]), .I1(VCC_net), 
            .CO(n48387));
    SB_LUT4 sub_38_add_2_5_lut (.I0(GND_net), .I1(n294[3]), .I2(VCC_net), 
            .I3(n48385), .O(\o_Rx_DV_N_3488[3] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i42760_2_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(GND_net), 
            .I3(GND_net), .O(n59812));
    defparam i42760_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i944_3_lut (.I0(n1263), .I1(n7924[21]), .I2(n294[16]), 
            .I3(GND_net), .O(n1410));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1008 (.I0(baudrate[17]), .I1(baudrate[18]), .I2(GND_net), 
            .I3(GND_net), .O(n59810));
    defparam i1_2_lut_adj_1008.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i1041_3_lut (.I0(n1410), .I1(n7950[21]), .I2(n294[15]), 
            .I3(GND_net), .O(n1554));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i42873_4_lut (.I0(n59014), .I1(n59010), .I2(n59012), .I3(n59008), 
            .O(n59926));
    defparam i42873_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i42915_4_lut (.I0(n59946), .I1(n59886), .I2(n56344), .I3(baudrate[4]), 
            .O(n59968));
    defparam i42915_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i49473_4_lut (.I0(n59926), .I1(n59810), .I2(n59968), .I3(n59812), 
            .O(n59974));
    defparam i49473_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 add_2749_8_lut (.I0(GND_net), .I1(n2104), .I2(n1602), .I3(n48889), 
            .O(n8080[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2743_5_lut (.I0(GND_net), .I1(n1265), .I2(n856), .I3(n48614), 
            .O(n7924[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1136_3_lut (.I0(n1554), .I1(n7976[21]), .I2(n294[14]), 
            .I3(GND_net), .O(n1695));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1229_3_lut (.I0(n1695), .I1(n8002[21]), .I2(n294[13]), 
            .I3(GND_net), .O(n1833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1320_3_lut (.I0(n1833), .I1(n8028[21]), .I2(n294[12]), 
            .I3(GND_net), .O(n1968));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1409_3_lut (.I0(n1968), .I1(n8054[21]), .I2(n294[11]), 
            .I3(GND_net), .O(n2100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1496_3_lut (.I0(n2100), .I1(n8080[21]), .I2(n294[10]), 
            .I3(GND_net), .O(n2229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i43_2_lut (.I0(n2229), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5066));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i23_2_lut (.I0(n2239), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5067));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46155_4_lut (.I0(n29_adj_5068), .I1(n27_adj_5069), .I2(n25_adj_5070), 
            .I3(n23_adj_5067), .O(n63217));
    defparam i46155_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46149_4_lut (.I0(n35_adj_5071), .I1(n33_adj_5072), .I2(n31_adj_5073), 
            .I3(n63217), .O(n63211));
    defparam i46149_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1517_i22_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2240), .I3(GND_net), .O(n22_adj_5074));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i22_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1517_i30_3_lut (.I0(n28_adj_5075), .I1(baudrate[7]), 
            .I2(n33_adj_5072), .I3(GND_net), .O(n30_adj_5076));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i34_3_lut (.I0(n26_adj_5077), .I1(baudrate[9]), 
            .I2(n37_adj_5078), .I3(GND_net), .O(n34));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49047_4_lut (.I0(n34), .I1(n24_adj_5079), .I2(n37_adj_5078), 
            .I3(n63207), .O(n66109));   // verilog/uart_rx.v(119[33:55])
    defparam i49047_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2743_5 (.CI(n48614), .I0(n1265), .I1(n856), .CO(n48615));
    SB_LUT4 i1_2_lut_4_lut (.I0(n66053), .I1(baudrate[18]), .I2(n2713), 
            .I3(n58484), .O(n2845));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h7100;
    SB_CARRY sub_38_add_2_5 (.CI(n48385), .I0(n294[3]), .I1(VCC_net), 
            .CO(n48386));
    SB_CARRY add_2749_8 (.CI(n48889), .I0(n2104), .I1(n1602), .CO(n48890));
    SB_LUT4 add_2743_4_lut (.I0(GND_net), .I1(n1266), .I2(n698), .I3(n48613), 
            .O(n7924[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_4_lut (.I0(GND_net), .I1(n294[2]), .I2(VCC_net), 
            .I3(n48384), .O(\o_Rx_DV_N_3488[2] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49048_3_lut (.I0(n66109), .I1(baudrate[10]), .I2(n39_adj_5080), 
            .I3(GND_net), .O(n66110));   // verilog/uart_rx.v(119[33:55])
    defparam i49048_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_38_add_2_4 (.CI(n48384), .I0(n294[2]), .I1(VCC_net), 
            .CO(n48385));
    SB_LUT4 i48926_3_lut (.I0(n66110), .I1(baudrate[11]), .I2(n41_adj_5081), 
            .I3(GND_net), .O(n65988));   // verilog/uart_rx.v(119[33:55])
    defparam i48926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48375_4_lut (.I0(n41_adj_5081), .I1(n39_adj_5080), .I2(n37_adj_5078), 
            .I3(n63211), .O(n65437));
    defparam i48375_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48699_4_lut (.I0(n30_adj_5076), .I1(n22_adj_5074), .I2(n33_adj_5072), 
            .I3(n63213), .O(n65761));   // verilog/uart_rx.v(119[33:55])
    defparam i48699_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2749_7_lut (.I0(GND_net), .I1(n2105), .I2(n1459), .I3(n48888), 
            .O(n8080[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_7 (.CI(n48888), .I0(n2105), .I1(n1459), .CO(n48889));
    SB_LUT4 add_2749_6_lut (.I0(GND_net), .I1(n2106), .I2(n1460), .I3(n48887), 
            .O(n8080[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2743_4 (.CI(n48613), .I0(n1266), .I1(n698), .CO(n48614));
    SB_LUT4 add_2743_3_lut (.I0(GND_net), .I1(n1267), .I2(n858), .I3(n48612), 
            .O(n7924[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_38_add_2_3_lut (.I0(GND_net), .I1(n294[1]), .I2(VCC_net), 
            .I3(n48383), .O(\o_Rx_DV_N_3488[1] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2743_3 (.CI(n48612), .I0(n1267), .I1(n858), .CO(n48613));
    SB_CARRY add_2749_6 (.CI(n48887), .I0(n2106), .I1(n1460), .CO(n48888));
    SB_LUT4 add_2749_5_lut (.I0(GND_net), .I1(n2107), .I2(n1011), .I3(n48886), 
            .O(n8080[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_5 (.CI(n48886), .I0(n2107), .I1(n1011), .CO(n48887));
    SB_LUT4 add_2749_4_lut (.I0(GND_net), .I1(n2108), .I2(n856), .I3(n48885), 
            .O(n8080[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_4 (.CI(n48885), .I0(n2108), .I1(n856), .CO(n48886));
    SB_LUT4 add_2743_2_lut (.I0(n56615), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n58470)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2743_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2749_3_lut (.I0(GND_net), .I1(n2109), .I2(n698), .I3(n48884), 
            .O(n8080[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2743_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n48612));
    SB_CARRY sub_38_add_2_3 (.CI(n48383), .I0(n294[1]), .I1(VCC_net), 
            .CO(n48384));
    SB_CARRY add_2749_3 (.CI(n48884), .I0(n2109), .I1(n698), .CO(n48885));
    SB_LUT4 sub_38_add_2_2_lut (.I0(GND_net), .I1(n57452), .I2(GND_net), 
            .I3(VCC_net), .O(\o_Rx_DV_N_3488[0] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_38_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_38_add_2_2 (.CI(VCC_net), .I0(n57452), .I1(GND_net), 
            .CO(n48383));
    SB_LUT4 i48782_3_lut (.I0(n65988), .I1(baudrate[12]), .I2(n43_adj_5066), 
            .I3(GND_net), .O(n42_adj_5082));   // verilog/uart_rx.v(119[33:55])
    defparam i48782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2749_2_lut (.I0(GND_net), .I1(n2110), .I2(n858), .I3(VCC_net), 
            .O(n8080[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2749_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2749_2 (.CI(VCC_net), .I0(n2110), .I1(n858), .CO(n48884));
    SB_DFFESR r_Clock_Count_2053__i0 (.Q(r_Clock_Count[0]), .C(clk16MHz), 
            .E(n27426), .D(n1[0]), .R(n28645));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 i48951_4_lut (.I0(n42_adj_5082), .I1(n65761), .I2(n43_adj_5066), 
            .I3(n65437), .O(n66013));   // verilog/uart_rx.v(119[33:55])
    defparam i48951_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48952_3_lut (.I0(n66013), .I1(baudrate[13]), .I2(n2228), 
            .I3(GND_net), .O(n66014));   // verilog/uart_rx.v(119[33:55])
    defparam i48952_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49449_2_lut_4_lut (.I0(n66053), .I1(baudrate[18]), .I2(n2713), 
            .I3(n25202), .O(n294[5]));   // verilog/uart_rx.v(119[33:55])
    defparam i49449_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i48507_3_lut (.I0(n66014), .I1(baudrate[14]), .I2(n2227), 
            .I3(GND_net), .O(n48_adj_5083));   // verilog/uart_rx.v(119[33:55])
    defparam i48507_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2742_8_lut (.I0(GND_net), .I1(n1111), .I2(n1459), .I3(n48602), 
            .O(n7898[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2742_7_lut (.I0(GND_net), .I1(n1112), .I2(n1460), .I3(n48601), 
            .O(n7898[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1009 (.I0(n25187), .I1(n48), .I2(baudrate[0]), 
            .I3(GND_net), .O(n2240));
    defparam i1_3_lut_adj_1009.LUT_INIT = 16'hefef;
    SB_LUT4 add_2758_25_lut (.I0(GND_net), .I1(n3151), .I2(n3186), .I3(n49090), 
            .O(n8314[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2758_24_lut (.I0(GND_net), .I1(n3152), .I2(n3082), .I3(n49089), 
            .O(n8314[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_24 (.CI(n49089), .I0(n3152), .I1(n3082), .CO(n49090));
    SB_LUT4 add_2758_23_lut (.I0(GND_net), .I1(n3153), .I2(n3188), .I3(n49088), 
            .O(n8314[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_23 (.CI(n49088), .I0(n3153), .I1(n3188), .CO(n49089));
    SB_LUT4 add_2758_22_lut (.I0(GND_net), .I1(n3154), .I2(n3084), .I3(n49087), 
            .O(n8314[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_22 (.CI(n49087), .I0(n3154), .I1(n3084), .CO(n49088));
    SB_LUT4 add_2758_21_lut (.I0(GND_net), .I1(n3155), .I2(n2977), .I3(n49086), 
            .O(n8314[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_21 (.CI(n49086), .I0(n3155), .I1(n2977), .CO(n49087));
    SB_LUT4 add_2758_20_lut (.I0(GND_net), .I1(n3156), .I2(n2867), .I3(n49085), 
            .O(n8314[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_20 (.CI(n49085), .I0(n3156), .I1(n2867), .CO(n49086));
    SB_LUT4 add_2758_19_lut (.I0(GND_net), .I1(n3157), .I2(n2754), .I3(n49084), 
            .O(n8314[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_19 (.CI(n49084), .I0(n3157), .I1(n2754), .CO(n49085));
    SB_CARRY add_2742_7 (.CI(n48601), .I0(n1112), .I1(n1460), .CO(n48602));
    SB_LUT4 add_2742_6_lut (.I0(GND_net), .I1(n1113), .I2(n1011), .I3(n48600), 
            .O(n7898[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2742_6 (.CI(n48600), .I0(n1113), .I1(n1011), .CO(n48601));
    SB_LUT4 add_2742_5_lut (.I0(GND_net), .I1(n1114), .I2(n856), .I3(n48599), 
            .O(n7898[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2742_5 (.CI(n48599), .I0(n1114), .I1(n856), .CO(n48600));
    SB_LUT4 add_2758_18_lut (.I0(GND_net), .I1(n3158), .I2(n2638), .I3(n49083), 
            .O(n8314[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_18 (.CI(n49083), .I0(n3158), .I1(n2638), .CO(n49084));
    SB_LUT4 add_2758_17_lut (.I0(GND_net), .I1(n3159), .I2(n2519), .I3(n49082), 
            .O(n8314[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_17 (.CI(n49082), .I0(n3159), .I1(n2519), .CO(n49083));
    SB_LUT4 add_2758_16_lut (.I0(GND_net), .I1(n3160), .I2(n2397), .I3(n49081), 
            .O(n8314[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_16 (.CI(n49081), .I0(n3160), .I1(n2397), .CO(n49082));
    SB_LUT4 add_2758_15_lut (.I0(GND_net), .I1(n3161), .I2(n2272), .I3(n49080), 
            .O(n8314[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_15 (.CI(n49080), .I0(n3161), .I1(n2272), .CO(n49081));
    SB_LUT4 add_2758_14_lut (.I0(GND_net), .I1(n3162), .I2(n2144), .I3(n49079), 
            .O(n8314[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_14 (.CI(n49079), .I0(n3162), .I1(n2144), .CO(n49080));
    SB_LUT4 add_2758_13_lut (.I0(GND_net), .I1(n3163), .I2(n2013), .I3(n49078), 
            .O(n8314[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_13 (.CI(n49078), .I0(n3163), .I1(n2013), .CO(n49079));
    SB_LUT4 add_2758_12_lut (.I0(GND_net), .I1(n3164), .I2(n1879), .I3(n49077), 
            .O(n8314[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_12 (.CI(n49077), .I0(n3164), .I1(n1879), .CO(n49078));
    SB_LUT4 add_2758_11_lut (.I0(GND_net), .I1(n3165), .I2(n1742), .I3(n49076), 
            .O(n8314[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_11 (.CI(n49076), .I0(n3165), .I1(n1742), .CO(n49077));
    SB_LUT4 add_2758_10_lut (.I0(GND_net), .I1(n3166), .I2(n1602), .I3(n49075), 
            .O(n8314[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_10 (.CI(n49075), .I0(n3166), .I1(n1602), .CO(n49076));
    SB_LUT4 add_2758_9_lut (.I0(GND_net), .I1(n3167), .I2(n1459), .I3(n49074), 
            .O(n8314[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_9 (.CI(n49074), .I0(n3167), .I1(n1459), .CO(n49075));
    SB_LUT4 add_2758_8_lut (.I0(GND_net), .I1(n3168), .I2(n1460), .I3(n49073), 
            .O(n8314[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_8 (.CI(n49073), .I0(n3168), .I1(n1460), .CO(n49074));
    SB_LUT4 div_37_i1592_3_lut (.I0(n2240), .I1(n8106[10]), .I2(n294[9]), 
            .I3(GND_net), .O(n2366));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2758_7_lut (.I0(GND_net), .I1(n3169), .I2(n1011), .I3(n49072), 
            .O(n8314[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_7 (.CI(n49072), .I0(n3169), .I1(n1011), .CO(n49073));
    SB_LUT4 add_2758_6_lut (.I0(GND_net), .I1(n3170), .I2(n856), .I3(n49071), 
            .O(n8314[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_6 (.CI(n49071), .I0(n3170), .I1(n856), .CO(n49072));
    SB_LUT4 add_2758_5_lut (.I0(GND_net), .I1(n3171), .I2(n698), .I3(n49070), 
            .O(n8314[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_5 (.CI(n49070), .I0(n3171), .I1(n698), .CO(n49071));
    SB_LUT4 add_2758_4_lut (.I0(GND_net), .I1(n3172), .I2(n858), .I3(n49069), 
            .O(n8314[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2742_4_lut (.I0(GND_net), .I1(n1115), .I2(n698), .I3(n48598), 
            .O(n7898[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2742_4 (.CI(n48598), .I0(n1115), .I1(n698), .CO(n48599));
    SB_LUT4 add_2742_3_lut (.I0(GND_net), .I1(n1116), .I2(n858), .I3(n48597), 
            .O(n7898[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2758_4 (.CI(n49069), .I0(n3172), .I1(n858), .CO(n49070));
    SB_LUT4 add_2758_3_lut (.I0(n56561), .I1(GND_net), .I2(n538), .I3(n49068), 
            .O(n58492)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2758_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2758_3 (.CI(n49068), .I0(GND_net), .I1(n538), .CO(n49069));
    SB_CARRY add_2758_2 (.CI(VCC_net), .I0(GND_net), .I1(VCC_net), .CO(n49068));
    SB_LUT4 add_2757_23_lut (.I0(GND_net), .I1(n3046), .I2(n3082), .I3(n49067), 
            .O(n8288[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2757_22_lut (.I0(GND_net), .I1(n3047), .I2(n3188), .I3(n49066), 
            .O(n8288[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_22 (.CI(n49066), .I0(n3047), .I1(n3188), .CO(n49067));
    SB_LUT4 add_2757_21_lut (.I0(GND_net), .I1(n3048), .I2(n3084), .I3(n49065), 
            .O(n8288[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_21 (.CI(n49065), .I0(n3048), .I1(n3084), .CO(n49066));
    SB_LUT4 add_2757_20_lut (.I0(GND_net), .I1(n3049), .I2(n2977), .I3(n49064), 
            .O(n8288[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_20 (.CI(n49064), .I0(n3049), .I1(n2977), .CO(n49065));
    SB_LUT4 add_2757_19_lut (.I0(GND_net), .I1(n3050), .I2(n2867), .I3(n49063), 
            .O(n8288[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_19 (.CI(n49063), .I0(n3050), .I1(n2867), .CO(n49064));
    SB_LUT4 add_2757_18_lut (.I0(GND_net), .I1(n3051), .I2(n2754), .I3(n49062), 
            .O(n8288[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_18 (.CI(n49062), .I0(n3051), .I1(n2754), .CO(n49063));
    SB_LUT4 add_2757_17_lut (.I0(GND_net), .I1(n3052), .I2(n2638), .I3(n49061), 
            .O(n8288[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2742_3 (.CI(n48597), .I0(n1116), .I1(n858), .CO(n48598));
    SB_CARRY add_2757_17 (.CI(n49061), .I0(n3052), .I1(n2638), .CO(n49062));
    SB_LUT4 add_2742_2_lut (.I0(n56619), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n58468)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2742_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2742_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n48597));
    SB_LUT4 add_2757_16_lut (.I0(GND_net), .I1(n3053), .I2(n2519), .I3(n49060), 
            .O(n8288[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_16 (.CI(n49060), .I0(n3053), .I1(n2519), .CO(n49061));
    SB_LUT4 add_2757_15_lut (.I0(GND_net), .I1(n3054), .I2(n2397), .I3(n49059), 
            .O(n8288[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_15 (.CI(n49059), .I0(n3054), .I1(n2397), .CO(n49060));
    SB_LUT4 add_2757_14_lut (.I0(GND_net), .I1(n3055), .I2(n2272), .I3(n49058), 
            .O(n8288[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_14 (.CI(n49058), .I0(n3055), .I1(n2272), .CO(n49059));
    SB_LUT4 add_2757_13_lut (.I0(GND_net), .I1(n3056), .I2(n2144), .I3(n49057), 
            .O(n8288[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i42649_2_lut (.I0(baudrate[17]), .I1(n25199), .I2(GND_net), 
            .I3(GND_net), .O(n59692));
    defparam i42649_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_2757_13 (.CI(n49057), .I0(n3056), .I1(n2144), .CO(n49058));
    SB_LUT4 add_2757_12_lut (.I0(GND_net), .I1(n3057), .I2(n2013), .I3(n49056), 
            .O(n8288[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_12 (.CI(n49056), .I0(n3057), .I1(n2013), .CO(n49057));
    SB_LUT4 add_2757_11_lut (.I0(GND_net), .I1(n3058), .I2(n1879), .I3(n49055), 
            .O(n8288[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_11 (.CI(n49055), .I0(n3058), .I1(n1879), .CO(n49056));
    SB_LUT4 add_2757_10_lut (.I0(GND_net), .I1(n3059), .I2(n1742), .I3(n49054), 
            .O(n8288[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_10 (.CI(n49054), .I0(n3059), .I1(n1742), .CO(n49055));
    SB_LUT4 add_2757_9_lut (.I0(GND_net), .I1(n3060), .I2(n1602), .I3(n49053), 
            .O(n8288[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1602_i21_2_lut (.I0(n2366), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46122_4_lut (.I0(n27_adj_5085), .I1(n25_adj_5086), .I2(n23_adj_5087), 
            .I3(n21_adj_5084), .O(n63184));
    defparam i46122_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2757_9 (.CI(n49053), .I0(n3060), .I1(n1602), .CO(n49054));
    SB_LUT4 add_2757_8_lut (.I0(GND_net), .I1(n3061), .I2(n1459), .I3(n49052), 
            .O(n8288[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_8 (.CI(n49052), .I0(n3061), .I1(n1459), .CO(n49053));
    SB_LUT4 add_2757_7_lut (.I0(GND_net), .I1(n3062), .I2(n1460), .I3(n49051), 
            .O(n8288[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_7 (.CI(n49051), .I0(n3062), .I1(n1460), .CO(n49052));
    SB_LUT4 add_2757_6_lut (.I0(GND_net), .I1(n3063), .I2(n1011), .I3(n49050), 
            .O(n8288[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47117_4_lut (.I0(n33_adj_5088), .I1(n31_adj_5089), .I2(n29_adj_5090), 
            .I3(n63184), .O(n64179));
    defparam i47117_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2757_6 (.CI(n49050), .I0(n3063), .I1(n1011), .CO(n49051));
    SB_LUT4 add_2757_5_lut (.I0(GND_net), .I1(n3064), .I2(n856), .I3(n49049), 
            .O(n8288[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_5 (.CI(n49049), .I0(n3064), .I1(n856), .CO(n49050));
    SB_LUT4 add_2757_4_lut (.I0(GND_net), .I1(n3065), .I2(n698), .I3(n49048), 
            .O(n8288[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_4 (.CI(n49048), .I0(n3065), .I1(n698), .CO(n49049));
    SB_LUT4 add_2757_3_lut (.I0(GND_net), .I1(n3066), .I2(n858), .I3(n49047), 
            .O(n8288[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2757_3 (.CI(n49047), .I0(n3066), .I1(n858), .CO(n49048));
    SB_LUT4 add_2757_2_lut (.I0(n56565), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n58490)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2757_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2757_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n49047));
    SB_LUT4 add_2756_22_lut (.I0(GND_net), .I1(n2938), .I2(n3188), .I3(n49046), 
            .O(n8262[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2756_21_lut (.I0(GND_net), .I1(n2939), .I2(n3084), .I3(n49045), 
            .O(n8262[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_21 (.CI(n49045), .I0(n2939), .I1(n3084), .CO(n49046));
    SB_LUT4 add_2756_20_lut (.I0(GND_net), .I1(n2940), .I2(n2977), .I3(n49044), 
            .O(n8262[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_20 (.CI(n49044), .I0(n2940), .I1(n2977), .CO(n49045));
    SB_LUT4 add_2756_19_lut (.I0(GND_net), .I1(n2941), .I2(n2867), .I3(n49043), 
            .O(n8262[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_19 (.CI(n49043), .I0(n2941), .I1(n2867), .CO(n49044));
    SB_LUT4 add_2756_18_lut (.I0(GND_net), .I1(n2942), .I2(n2754), .I3(n49042), 
            .O(n8262[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_18 (.CI(n49042), .I0(n2942), .I1(n2754), .CO(n49043));
    SB_LUT4 add_2756_17_lut (.I0(GND_net), .I1(n2943), .I2(n2638), .I3(n49041), 
            .O(n8262[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_17 (.CI(n49041), .I0(n2943), .I1(n2638), .CO(n49042));
    SB_LUT4 add_2756_16_lut (.I0(GND_net), .I1(n2944), .I2(n2519), .I3(n49040), 
            .O(n8262[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_16 (.CI(n49040), .I0(n2944), .I1(n2519), .CO(n49041));
    SB_LUT4 add_2756_15_lut (.I0(GND_net), .I1(n2945), .I2(n2397), .I3(n49039), 
            .O(n8262[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_15 (.CI(n49039), .I0(n2945), .I1(n2397), .CO(n49040));
    SB_LUT4 add_2756_14_lut (.I0(GND_net), .I1(n2946), .I2(n2272), .I3(n49038), 
            .O(n8262[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_14 (.CI(n49038), .I0(n2946), .I1(n2272), .CO(n49039));
    SB_LUT4 add_2756_13_lut (.I0(GND_net), .I1(n2947), .I2(n2144), .I3(n49037), 
            .O(n8262[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_13 (.CI(n49037), .I0(n2947), .I1(n2144), .CO(n49038));
    SB_LUT4 add_2756_12_lut (.I0(GND_net), .I1(n2948), .I2(n2013), .I3(n49036), 
            .O(n8262[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_12 (.CI(n49036), .I0(n2948), .I1(n2013), .CO(n49037));
    SB_LUT4 add_2756_11_lut (.I0(GND_net), .I1(n2949), .I2(n1879), .I3(n49035), 
            .O(n8262[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49316_3_lut (.I0(n25229), .I1(baudrate[1]), .I2(baudrate[2]), 
            .I3(GND_net), .O(n25108));   // verilog/uart_rx.v(119[33:55])
    defparam i49316_3_lut.LUT_INIT = 16'h0101;
    SB_CARRY add_2756_11 (.CI(n49035), .I0(n2949), .I1(n1879), .CO(n49036));
    SB_LUT4 add_2756_10_lut (.I0(GND_net), .I1(n2950), .I2(n1742), .I3(n49034), 
            .O(n8262[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_10 (.CI(n49034), .I0(n2950), .I1(n1742), .CO(n49035));
    SB_LUT4 add_2756_9_lut (.I0(GND_net), .I1(n2951), .I2(n1602), .I3(n49033), 
            .O(n8262[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_9 (.CI(n49033), .I0(n2951), .I1(n1602), .CO(n49034));
    SB_LUT4 add_2756_8_lut (.I0(GND_net), .I1(n2952), .I2(n1459), .I3(n49032), 
            .O(n8262[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_8 (.CI(n49032), .I0(n2952), .I1(n1459), .CO(n49033));
    SB_LUT4 add_2756_7_lut (.I0(GND_net), .I1(n2953), .I2(n1460), .I3(n49031), 
            .O(n8262[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_7 (.CI(n49031), .I0(n2953), .I1(n1460), .CO(n49032));
    SB_LUT4 add_2756_6_lut (.I0(GND_net), .I1(n2954), .I2(n1011), .I3(n49030), 
            .O(n8262[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_6 (.CI(n49030), .I0(n2954), .I1(n1011), .CO(n49031));
    SB_LUT4 add_2756_5_lut (.I0(GND_net), .I1(n2955), .I2(n856), .I3(n49029), 
            .O(n8262[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_5 (.CI(n49029), .I0(n2955), .I1(n856), .CO(n49030));
    SB_LUT4 add_2756_4_lut (.I0(GND_net), .I1(n2956), .I2(n698), .I3(n49028), 
            .O(n8262[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_4 (.CI(n49028), .I0(n2956), .I1(n698), .CO(n49029));
    SB_LUT4 add_2756_3_lut (.I0(GND_net), .I1(n2957), .I2(n858), .I3(n49027), 
            .O(n8262[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2756_3 (.CI(n49027), .I0(n2957), .I1(n858), .CO(n49028));
    SB_LUT4 add_2756_2_lut (.I0(n56569), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n58488)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2756_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2756_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n49027));
    SB_LUT4 div_37_LessThan_1602_i28_3_lut (.I0(n26_adj_5091), .I1(baudrate[7]), 
            .I2(n31_adj_5089), .I3(GND_net), .O(n28_adj_5092));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2755_21_lut (.I0(GND_net), .I1(n2827), .I2(n3084), .I3(n49026), 
            .O(n8236[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2755_20_lut (.I0(GND_net), .I1(n2828), .I2(n2977), .I3(n49025), 
            .O(n8236[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_20 (.CI(n49025), .I0(n2828), .I1(n2977), .CO(n49026));
    SB_LUT4 add_2755_19_lut (.I0(GND_net), .I1(n2829), .I2(n2867), .I3(n49024), 
            .O(n8236[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_19 (.CI(n49024), .I0(n2829), .I1(n2867), .CO(n49025));
    SB_LUT4 div_37_LessThan_1602_i32_3_lut (.I0(n24_adj_5093), .I1(baudrate[9]), 
            .I2(n35_adj_5094), .I3(GND_net), .O(n32));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2755_18_lut (.I0(GND_net), .I1(n2830), .I2(n2754), .I3(n49023), 
            .O(n8236[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_18 (.CI(n49023), .I0(n2830), .I1(n2754), .CO(n49024));
    SB_LUT4 add_2755_17_lut (.I0(GND_net), .I1(n2831), .I2(n2638), .I3(n49022), 
            .O(n8236[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_17 (.CI(n49022), .I0(n2831), .I1(n2638), .CO(n49023));
    SB_LUT4 add_2755_16_lut (.I0(GND_net), .I1(n2832), .I2(n2519), .I3(n49021), 
            .O(n8236[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_16 (.CI(n49021), .I0(n2832), .I1(n2519), .CO(n49022));
    SB_LUT4 i48911_4_lut (.I0(n32), .I1(n22_adj_5095), .I2(n35_adj_5094), 
            .I3(n64171), .O(n65973));   // verilog/uart_rx.v(119[33:55])
    defparam i48911_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48912_3_lut (.I0(n65973), .I1(baudrate[10]), .I2(n37_adj_5096), 
            .I3(GND_net), .O(n65974));   // verilog/uart_rx.v(119[33:55])
    defparam i48912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48802_3_lut (.I0(n65974), .I1(baudrate[11]), .I2(n39_adj_5097), 
            .I3(GND_net), .O(n65864));   // verilog/uart_rx.v(119[33:55])
    defparam i48802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2171_1_lut (.I0(baudrate[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1011));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2171_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2755_15_lut (.I0(GND_net), .I1(n2833), .I2(n2397), .I3(n49020), 
            .O(n8236[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_15 (.CI(n49020), .I0(n2833), .I1(n2397), .CO(n49021));
    SB_LUT4 add_2755_14_lut (.I0(GND_net), .I1(n2834), .I2(n2272), .I3(n49019), 
            .O(n8236[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_14 (.CI(n49019), .I0(n2834), .I1(n2272), .CO(n49020));
    SB_LUT4 add_2755_13_lut (.I0(GND_net), .I1(n2835), .I2(n2144), .I3(n49018), 
            .O(n8236[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1674_3_lut (.I0(n2365), .I1(n8132[11]), .I2(n294[8]), 
            .I3(GND_net), .O(n2488));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2755_13 (.CI(n49018), .I0(n2835), .I1(n2144), .CO(n49019));
    SB_LUT4 add_2755_12_lut (.I0(GND_net), .I1(n2836), .I2(n2013), .I3(n49017), 
            .O(n8236[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_12 (.CI(n49017), .I0(n2836), .I1(n2013), .CO(n49018));
    SB_LUT4 add_2755_11_lut (.I0(GND_net), .I1(n2837), .I2(n1879), .I3(n49016), 
            .O(n8236[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48681_4_lut (.I0(n39_adj_5097), .I1(n37_adj_5096), .I2(n35_adj_5094), 
            .I3(n64179), .O(n65743));
    defparam i48681_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48913_4_lut (.I0(n28_adj_5092), .I1(n20_adj_5098), .I2(n31_adj_5089), 
            .I3(n63182), .O(n65975));   // verilog/uart_rx.v(119[33:55])
    defparam i48913_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2755_11 (.CI(n49016), .I0(n2837), .I1(n1879), .CO(n49017));
    SB_LUT4 add_2755_10_lut (.I0(GND_net), .I1(n2838), .I2(n1742), .I3(n49015), 
            .O(n8236[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_10 (.CI(n49015), .I0(n2838), .I1(n1742), .CO(n49016));
    SB_LUT4 add_2755_9_lut (.I0(GND_net), .I1(n2839), .I2(n1602), .I3(n49014), 
            .O(n8236[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_9 (.CI(n49014), .I0(n2839), .I1(n1602), .CO(n49015));
    SB_LUT4 add_2755_8_lut (.I0(GND_net), .I1(n2840), .I2(n1459), .I3(n49013), 
            .O(n8236[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_8 (.CI(n49013), .I0(n2840), .I1(n1459), .CO(n49014));
    SB_LUT4 add_2755_7_lut (.I0(GND_net), .I1(n2841), .I2(n1460), .I3(n49012), 
            .O(n8236[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_7 (.CI(n49012), .I0(n2841), .I1(n1460), .CO(n49013));
    SB_LUT4 add_2755_6_lut (.I0(GND_net), .I1(n2842), .I2(n1011), .I3(n49011), 
            .O(n8236[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_6 (.CI(n49011), .I0(n2842), .I1(n1011), .CO(n49012));
    SB_LUT4 add_2755_5_lut (.I0(GND_net), .I1(n2843), .I2(n856), .I3(n49010), 
            .O(n8236[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_5 (.CI(n49010), .I0(n2843), .I1(n856), .CO(n49011));
    SB_LUT4 add_2755_4_lut (.I0(GND_net), .I1(n2844), .I2(n698), .I3(n49009), 
            .O(n8236[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_4 (.CI(n49009), .I0(n2844), .I1(n698), .CO(n49010));
    SB_LUT4 add_2755_3_lut (.I0(GND_net), .I1(n2845), .I2(n858), .I3(n49008), 
            .O(n8236[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2755_3 (.CI(n49008), .I0(n2845), .I1(n858), .CO(n49009));
    SB_LUT4 add_2755_2_lut (.I0(n56573), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n58486)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2755_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2755_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n49008));
    SB_LUT4 add_2754_20_lut (.I0(GND_net), .I1(n2713), .I2(n2977), .I3(n49007), 
            .O(n8210[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_20_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR r_Clock_Count_2053__i7 (.Q(r_Clock_Count[7]), .C(clk16MHz), 
            .E(n27426), .D(n1[7]), .R(n28645));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i6 (.Q(r_Clock_Count[6]), .C(clk16MHz), 
            .E(n27426), .D(n1[6]), .R(n28645));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i5 (.Q(r_Clock_Count[5]), .C(clk16MHz), 
            .E(n27426), .D(n1[5]), .R(n28645));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i4 (.Q(r_Clock_Count[4]), .C(clk16MHz), 
            .E(n27426), .D(n1[4]), .R(n28645));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i3 (.Q(r_Clock_Count[3]), .C(clk16MHz), 
            .E(n27426), .D(n1[3]), .R(n28645));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i2 (.Q(r_Clock_Count[2]), .C(clk16MHz), 
            .E(n27426), .D(n1[2]), .R(n28645));   // verilog/uart_rx.v(121[34:51])
    SB_DFFESR r_Clock_Count_2053__i1 (.Q(r_Clock_Count[1]), .C(clk16MHz), 
            .E(n27426), .D(n1[1]), .R(n28645));   // verilog/uart_rx.v(121[34:51])
    SB_LUT4 add_2754_19_lut (.I0(GND_net), .I1(n2714), .I2(n2867), .I3(n49006), 
            .O(n8210[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_19 (.CI(n49006), .I0(n2714), .I1(n2867), .CO(n49007));
    SB_LUT4 i47385_3_lut (.I0(n65864), .I1(baudrate[12]), .I2(n41_adj_5099), 
            .I3(GND_net), .O(n64447));   // verilog/uart_rx.v(119[33:55])
    defparam i47385_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2754_18_lut (.I0(GND_net), .I1(n2715), .I2(n2754), .I3(n49005), 
            .O(n8210[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_18 (.CI(n49005), .I0(n2715), .I1(n2754), .CO(n49006));
    SB_LUT4 add_2754_17_lut (.I0(GND_net), .I1(n2716), .I2(n2638), .I3(n49004), 
            .O(n8210[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_17 (.CI(n49004), .I0(n2716), .I1(n2638), .CO(n49005));
    SB_LUT4 add_2754_16_lut (.I0(GND_net), .I1(n2717), .I2(n2519), .I3(n49003), 
            .O(n8210[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46254_3_lut_4_lut (.I0(n1699), .I1(baudrate[4]), .I2(baudrate[3]), 
            .I3(n1700), .O(n63316));   // verilog/uart_rx.v(119[33:55])
    defparam i46254_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1157_i34_3_lut_3_lut (.I0(n1699), .I1(baudrate[4]), 
            .I2(baudrate[3]), .I3(GND_net), .O(n34_adj_5100));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i49074_4_lut (.I0(n64447), .I1(n65975), .I2(n41_adj_5099), 
            .I3(n65743), .O(n66136));   // verilog/uart_rx.v(119[33:55])
    defparam i49074_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49075_3_lut (.I0(n66136), .I1(baudrate[13]), .I2(n2355), 
            .I3(GND_net), .O(n66137));   // verilog/uart_rx.v(119[33:55])
    defparam i49075_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2754_16 (.CI(n49003), .I0(n2717), .I1(n2519), .CO(n49004));
    SB_LUT4 add_2754_15_lut (.I0(GND_net), .I1(n2718), .I2(n2397), .I3(n49002), 
            .O(n8210[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_15 (.CI(n49002), .I0(n2718), .I1(n2397), .CO(n49003));
    SB_LUT4 add_2754_14_lut (.I0(GND_net), .I1(n2719), .I2(n2272), .I3(n49001), 
            .O(n8210[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_14 (.CI(n49001), .I0(n2719), .I1(n2272), .CO(n49002));
    SB_LUT4 add_2754_13_lut (.I0(GND_net), .I1(n2720), .I2(n2144), .I3(n49000), 
            .O(n8210[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_13 (.CI(n49000), .I0(n2720), .I1(n2144), .CO(n49001));
    SB_LUT4 add_2754_12_lut (.I0(GND_net), .I1(n2721), .I2(n2013), .I3(n48999), 
            .O(n8210[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_12 (.CI(n48999), .I0(n2721), .I1(n2013), .CO(n49000));
    SB_LUT4 add_2754_11_lut (.I0(GND_net), .I1(n2722), .I2(n1879), .I3(n48998), 
            .O(n8210[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_11 (.CI(n48998), .I0(n2722), .I1(n1879), .CO(n48999));
    SB_LUT4 div_37_LessThan_1250_i39_2_lut (.I0(n1835), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1250_i37_2_lut (.I0(n1836), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2754_10_lut (.I0(GND_net), .I1(n2723), .I2(n1742), .I3(n48997), 
            .O(n8210[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_10 (.CI(n48997), .I0(n2723), .I1(n1742), .CO(n48998));
    SB_LUT4 add_2754_9_lut (.I0(GND_net), .I1(n2724), .I2(n1602), .I3(n48996), 
            .O(n8210[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_9 (.CI(n48996), .I0(n2724), .I1(n1602), .CO(n48997));
    SB_LUT4 add_2754_8_lut (.I0(GND_net), .I1(n2725), .I2(n1459), .I3(n48995), 
            .O(n8210[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1250_i43_2_lut (.I0(n1833), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i43_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_2754_8 (.CI(n48995), .I0(n2725), .I1(n1459), .CO(n48996));
    SB_LUT4 i48997_3_lut (.I0(n66137), .I1(baudrate[14]), .I2(n2354), 
            .I3(GND_net), .O(n66059));   // verilog/uart_rx.v(119[33:55])
    defparam i48997_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1250_i31_2_lut (.I0(n1839), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46267_3_lut_4_lut (.I0(n1558), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1559), .O(n63329));   // verilog/uart_rx.v(119[33:55])
    defparam i46267_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_2754_7_lut (.I0(GND_net), .I1(n2726), .I2(n1460), .I3(n48994), 
            .O(n8210[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1250_i33_2_lut (.I0(n1838), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1062_i34_3_lut_3_lut (.I0(n1558), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n34_adj_5106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i34_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_LessThan_1250_i35_2_lut (.I0(n1837), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47391_3_lut (.I0(n66059), .I1(baudrate[15]), .I2(n2353), 
            .I3(GND_net), .O(n48_adj_5108));   // verilog/uart_rx.v(119[33:55])
    defparam i47391_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1250_i41_2_lut (.I0(n1834), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46279_3_lut_4_lut (.I0(n1413), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1414), .O(n63341));   // verilog/uart_rx.v(119[33:55])
    defparam i46279_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1250_i29_2_lut (.I0(n1840), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5110));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46212_4_lut (.I0(n35_adj_5107), .I1(n33_adj_5105), .I2(n31_adj_5104), 
            .I3(n29_adj_5110), .O(n63274));
    defparam i46212_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2754_7 (.CI(n48994), .I0(n2726), .I1(n1460), .CO(n48995));
    SB_LUT4 add_2754_6_lut (.I0(GND_net), .I1(n2727), .I2(n1011), .I3(n48993), 
            .O(n8210[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_965_i36_3_lut_3_lut (.I0(n1413), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n36));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i36_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk16MHz), .E(n27312), 
            .D(n479[1]), .R(n28373));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 div_37_LessThan_765_i40_3_lut_3_lut (.I0(n1114), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n40_adj_5111));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i40_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_i1590_3_lut (.I0(n2238), .I1(n8106[12]), .I2(n294[9]), 
            .I3(GND_net), .O(n2364));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2170_1_lut (.I0(baudrate[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1460));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2170_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk16MHz), .E(n27312), 
            .D(n479[2]), .R(n28373));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2754_6 (.CI(n48993), .I0(n2727), .I1(n1011), .CO(n48994));
    SB_LUT4 add_2754_5_lut (.I0(GND_net), .I1(n2728), .I2(n856), .I3(n48992), 
            .O(n8210[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_5 (.CI(n48992), .I0(n2728), .I1(n856), .CO(n48993));
    SB_LUT4 div_37_i1673_3_lut (.I0(n2364), .I1(n8132[12]), .I2(n294[8]), 
            .I3(GND_net), .O(n2487));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2754_4_lut (.I0(GND_net), .I1(n2729), .I2(n698), .I3(n48991), 
            .O(n8210[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2754_4 (.CI(n48991), .I0(n2729), .I1(n698), .CO(n48992));
    SB_LUT4 add_2754_3_lut (.I0(GND_net), .I1(n2730), .I2(n858), .I3(n48990), 
            .O(n8210[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_1250_i40_3_lut (.I0(n32_adj_5112), .I1(baudrate[9]), 
            .I2(n43_adj_5103), .I3(GND_net), .O(n40_adj_5113));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1250_i28_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1841), .I3(GND_net), .O(n28_adj_5114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i28_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48723_3_lut (.I0(n28_adj_5114), .I1(baudrate[5]), .I2(n35_adj_5107), 
            .I3(GND_net), .O(n65785));   // verilog/uart_rx.v(119[33:55])
    defparam i48723_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2754_3 (.CI(n48990), .I0(n2730), .I1(n858), .CO(n48991));
    SB_LUT4 add_2754_2_lut (.I0(n56577), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n58484)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2754_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2754_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n48990));
    SB_LUT4 add_2753_19_lut (.I0(GND_net), .I1(n2596), .I2(n2867), .I3(n48989), 
            .O(n8184[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2753_18_lut (.I0(GND_net), .I1(n2597), .I2(n2754), .I3(n48988), 
            .O(n8184[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_18 (.CI(n48988), .I0(n2597), .I1(n2754), .CO(n48989));
    SB_LUT4 add_2753_17_lut (.I0(GND_net), .I1(n2598), .I2(n2638), .I3(n48987), 
            .O(n8184[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48724_3_lut (.I0(n65785), .I1(baudrate[6]), .I2(n37_adj_5102), 
            .I3(GND_net), .O(n65786));   // verilog/uart_rx.v(119[33:55])
    defparam i48724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46208_4_lut (.I0(n41_adj_5109), .I1(n39_adj_5101), .I2(n37_adj_5102), 
            .I3(n63274), .O(n63270));
    defparam i46208_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48721_4_lut (.I0(n40_adj_5113), .I1(n30_adj_5115), .I2(n43_adj_5103), 
            .I3(n63266), .O(n65783));   // verilog/uart_rx.v(119[33:55])
    defparam i48721_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2753_17 (.CI(n48987), .I0(n2598), .I1(n2638), .CO(n48988));
    SB_LUT4 add_2753_16_lut (.I0(GND_net), .I1(n2599), .I2(n2519), .I3(n48986), 
            .O(n8184[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_16 (.CI(n48986), .I0(n2599), .I1(n2519), .CO(n48987));
    SB_LUT4 i46295_3_lut_4_lut (.I0(n1114), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1115), .O(n63357));   // verilog/uart_rx.v(119[33:55])
    defparam i46295_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i48489_3_lut (.I0(n65786), .I1(baudrate[7]), .I2(n39_adj_5101), 
            .I3(GND_net), .O(n65551));   // verilog/uart_rx.v(119[33:55])
    defparam i48489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49032_4_lut (.I0(n65551), .I1(n65783), .I2(n43_adj_5103), 
            .I3(n63270), .O(n66094));   // verilog/uart_rx.v(119[33:55])
    defparam i49032_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2753_15_lut (.I0(GND_net), .I1(n2600), .I2(n2397), .I3(n48985), 
            .O(n8184[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49033_3_lut (.I0(n66094), .I1(baudrate[10]), .I2(n1832), 
            .I3(GND_net), .O(n66095));   // verilog/uart_rx.v(119[33:55])
    defparam i49033_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2753_15 (.CI(n48985), .I0(n2600), .I1(n2397), .CO(n48986));
    SB_LUT4 add_2753_14_lut (.I0(GND_net), .I1(n2601), .I2(n2272), .I3(n48984), 
            .O(n8184[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1418_3_lut (.I0(n1977), .I1(n8054[12]), .I2(n294[11]), 
            .I3(GND_net), .O(n2109));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1505_3_lut (.I0(n2109), .I1(n8080[12]), .I2(n294[10]), 
            .I3(GND_net), .O(n2238));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1579_3_lut (.I0(n2227), .I1(n8106[23]), .I2(n294[9]), 
            .I3(GND_net), .O(n2353));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1010 (.I0(n59308), .I1(n58424), .I2(n58422), 
            .I3(n59298), .O(n25199));
    defparam i1_4_lut_adj_1010.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1580_3_lut (.I0(n2228), .I1(n8106[22]), .I2(n294[9]), 
            .I3(GND_net), .O(n2354));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1580_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2753_14 (.CI(n48984), .I0(n2601), .I1(n2272), .CO(n48985));
    SB_LUT4 div_37_i1581_3_lut (.I0(n2229), .I1(n8106[21]), .I2(n294[9]), 
            .I3(GND_net), .O(n2355));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1410_3_lut (.I0(n1969), .I1(n8054[20]), .I2(n294[11]), 
            .I3(GND_net), .O(n2101));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1497_3_lut (.I0(n2101), .I1(n8080[20]), .I2(n294[10]), 
            .I3(GND_net), .O(n2230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1582_3_lut (.I0(n2230), .I1(n8106[20]), .I2(n294[9]), 
            .I3(GND_net), .O(n2356));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i41_2_lut (.I0(n2356), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1139_3_lut (.I0(n1557), .I1(n7976[18]), .I2(n294[14]), 
            .I3(GND_net), .O(n1698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1232_3_lut (.I0(n1698), .I1(n8002[18]), .I2(n294[13]), 
            .I3(GND_net), .O(n1836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1323_3_lut (.I0(n1836), .I1(n8028[18]), .I2(n294[12]), 
            .I3(GND_net), .O(n1971));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2748_14_lut (.I0(GND_net), .I1(n1966), .I2(n2272), .I3(n48814), 
            .O(n8054[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2748_13_lut (.I0(GND_net), .I1(n1967), .I2(n2144), .I3(n48813), 
            .O(n8054[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1412_3_lut (.I0(n1971), .I1(n8054[18]), .I2(n294[11]), 
            .I3(GND_net), .O(n2103));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1499_3_lut (.I0(n2103), .I1(n8080[18]), .I2(n294[10]), 
            .I3(GND_net), .O(n2232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1584_3_lut (.I0(n2232), .I1(n8106[18]), .I2(n294[9]), 
            .I3(GND_net), .O(n2358));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1584_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2748_13 (.CI(n48813), .I0(n1967), .I1(n2144), .CO(n48814));
    SB_LUT4 add_2748_12_lut (.I0(GND_net), .I1(n1968), .I2(n2013), .I3(n48812), 
            .O(n8054[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_12 (.CI(n48812), .I0(n1968), .I1(n2013), .CO(n48813));
    SB_LUT4 div_37_LessThan_1602_i37_2_lut (.I0(n2358), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5096));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1043_3_lut (.I0(n1412), .I1(n7950[19]), .I2(n294[15]), 
            .I3(GND_net), .O(n1556));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1138_3_lut (.I0(n1556), .I1(n7976[19]), .I2(n294[14]), 
            .I3(GND_net), .O(n1697));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2748_11_lut (.I0(GND_net), .I1(n1969), .I2(n1879), .I3(n48811), 
            .O(n8054[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_11 (.CI(n48811), .I0(n1969), .I1(n1879), .CO(n48812));
    SB_LUT4 div_37_i1231_3_lut (.I0(n1697), .I1(n8002[19]), .I2(n294[13]), 
            .I3(GND_net), .O(n1835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1322_3_lut (.I0(n1835), .I1(n8028[19]), .I2(n294[12]), 
            .I3(GND_net), .O(n1970));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1411_3_lut (.I0(n1970), .I1(n8054[19]), .I2(n294[11]), 
            .I3(GND_net), .O(n2102));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1498_3_lut (.I0(n2102), .I1(n8080[19]), .I2(n294[10]), 
            .I3(GND_net), .O(n2231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2748_10_lut (.I0(GND_net), .I1(n1970), .I2(n1742), .I3(n48810), 
            .O(n8054[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_10 (.CI(n48810), .I0(n1970), .I1(n1742), .CO(n48811));
    SB_LUT4 div_37_i1583_3_lut (.I0(n2231), .I1(n8106[19]), .I2(n294[9]), 
            .I3(GND_net), .O(n2357));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i39_2_lut (.I0(n2357), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5097));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i948_3_lut (.I0(n1267), .I1(n7924[17]), .I2(n294[16]), 
            .I3(GND_net), .O(n1414));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1045_3_lut (.I0(n1414), .I1(n7950[17]), .I2(n294[15]), 
            .I3(GND_net), .O(n1558));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1140_3_lut (.I0(n1558), .I1(n7976[17]), .I2(n294[14]), 
            .I3(GND_net), .O(n1699));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2748_9_lut (.I0(GND_net), .I1(n1971), .I2(n1602), .I3(n48809), 
            .O(n8054[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_i1233_3_lut (.I0(n1699), .I1(n8002[17]), .I2(n294[13]), 
            .I3(GND_net), .O(n1837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1324_3_lut (.I0(n1837), .I1(n8028[17]), .I2(n294[12]), 
            .I3(GND_net), .O(n1972));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1413_3_lut (.I0(n1972), .I1(n8054[17]), .I2(n294[11]), 
            .I3(GND_net), .O(n2104));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1500_3_lut (.I0(n2104), .I1(n8080[17]), .I2(n294[10]), 
            .I3(GND_net), .O(n2233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2753_13_lut (.I0(GND_net), .I1(n2602), .I2(n2144), .I3(n48983), 
            .O(n8184[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i39551_1_lut (.I0(n25211), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56565));
    defparam i39551_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2748_9 (.CI(n48809), .I0(n1971), .I1(n1602), .CO(n48810));
    SB_CARRY add_2753_13 (.CI(n48983), .I0(n2602), .I1(n2144), .CO(n48984));
    SB_LUT4 div_37_i1585_3_lut (.I0(n2233), .I1(n8106[17]), .I2(n294[9]), 
            .I3(GND_net), .O(n2359));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2748_8_lut (.I0(GND_net), .I1(n1972), .I2(n1459), .I3(n48808), 
            .O(n8054[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_8 (.CI(n48808), .I0(n1972), .I1(n1459), .CO(n48809));
    SB_LUT4 add_2748_7_lut (.I0(GND_net), .I1(n1973), .I2(n1460), .I3(n48807), 
            .O(n8054[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_7 (.CI(n48807), .I0(n1973), .I1(n1460), .CO(n48808));
    SB_LUT4 div_37_LessThan_1602_i35_2_lut (.I0(n2359), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5094));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2748_6_lut (.I0(GND_net), .I1(n1974), .I2(n1011), .I3(n48806), 
            .O(n8054[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2753_12_lut (.I0(GND_net), .I1(n2603), .I2(n2013), .I3(n48982), 
            .O(n8184[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_6 (.CI(n48806), .I0(n1974), .I1(n1011), .CO(n48807));
    SB_CARRY add_2753_12 (.CI(n48982), .I0(n2603), .I1(n2013), .CO(n48983));
    SB_LUT4 add_2748_5_lut (.I0(GND_net), .I1(n1975), .I2(n856), .I3(n48805), 
            .O(n8054[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_5 (.CI(n48805), .I0(n1975), .I1(n856), .CO(n48806));
    SB_LUT4 add_2748_4_lut (.I0(GND_net), .I1(n1976), .I2(n698), .I3(n48804), 
            .O(n8054[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_4 (.CI(n48804), .I0(n1976), .I1(n698), .CO(n48805));
    SB_LUT4 i1_2_lut_adj_1011 (.I0(n58476), .I1(n48_adj_5083), .I2(GND_net), 
            .I3(GND_net), .O(n2367));
    defparam i1_2_lut_adj_1011.LUT_INIT = 16'h2222;
    SB_LUT4 add_2748_3_lut (.I0(GND_net), .I1(n1977), .I2(n858), .I3(n48803), 
            .O(n8054[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_3 (.CI(n48803), .I0(n1977), .I1(n858), .CO(n48804));
    SB_LUT4 add_2748_2_lut (.I0(GND_net), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n8054[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2748_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2753_11_lut (.I0(GND_net), .I1(n2604), .I2(n1879), .I3(n48981), 
            .O(n8184[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2748_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n48803));
    SB_CARRY add_2753_11 (.CI(n48981), .I0(n2604), .I1(n1879), .CO(n48982));
    SB_LUT4 div_37_LessThan_866_i41_2_lut (.I0(n1264), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5116));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_2753_10_lut (.I0(GND_net), .I1(n2605), .I2(n1742), .I3(n48980), 
            .O(n8184[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_10 (.CI(n48980), .I0(n2605), .I1(n1742), .CO(n48981));
    SB_LUT4 div_37_LessThan_765_i38_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1116), .I3(GND_net), .O(n38_adj_5117));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i38_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk16MHz), .D(n29592));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_DV_58 (.Q(rx_data_ready), .C(clk16MHz), .D(n51425));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2753_9_lut (.I0(GND_net), .I1(n2606), .I2(n1602), .I3(n48979), 
            .O(n8184[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_9 (.CI(n48979), .I0(n2606), .I1(n1602), .CO(n48980));
    SB_LUT4 add_2747_13_lut (.I0(GND_net), .I1(n1831), .I2(n2144), .I3(n48784), 
            .O(n8028[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk16MHz), .D(n29596));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2747_12_lut (.I0(GND_net), .I1(n1832), .I2(n2013), .I3(n48783), 
            .O(n8028[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2753_8_lut (.I0(GND_net), .I1(n2607), .I2(n1459), .I3(n48978), 
            .O(n8184[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk16MHz), .D(n29582));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2747_12 (.CI(n48783), .I0(n1832), .I1(n2013), .CO(n48784));
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk16MHz), .D(n29581));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk16MHz), .D(n29580));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk16MHz), .D(n29578));   // verilog/uart_rx.v(50[10] 145[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk16MHz), .D(n29577));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2747_11_lut (.I0(GND_net), .I1(n1833), .I2(n1879), .I3(n48782), 
            .O(n8028[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_11 (.CI(n48782), .I0(n1833), .I1(n1879), .CO(n48783));
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk16MHz), .D(n29576));   // verilog/uart_rx.v(50[10] 145[8])
    SB_CARRY add_2753_8 (.CI(n48978), .I0(n2607), .I1(n1459), .CO(n48979));
    SB_LUT4 add_2753_7_lut (.I0(GND_net), .I1(n2608), .I2(n1460), .I3(n48977), 
            .O(n8184[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk16MHz), .D(n29575));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2747_10_lut (.I0(GND_net), .I1(n1834), .I2(n1742), .I3(n48781), 
            .O(n8028[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_10 (.CI(n48781), .I0(n1834), .I1(n1742), .CO(n48782));
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk16MHz), .D(n67140));   // verilog/uart_rx.v(50[10] 145[8])
    SB_LUT4 add_2747_9_lut (.I0(GND_net), .I1(n1835), .I2(n1602), .I3(n48780), 
            .O(n8028[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_9 (.CI(n48780), .I0(n1835), .I1(n1602), .CO(n48781));
    SB_LUT4 add_2747_8_lut (.I0(GND_net), .I1(n1836), .I2(n1459), .I3(n48779), 
            .O(n8028[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_8 (.CI(n48779), .I0(n1836), .I1(n1459), .CO(n48780));
    SB_LUT4 add_2747_7_lut (.I0(GND_net), .I1(n1837), .I2(n1460), .I3(n48778), 
            .O(n8028[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_7 (.CI(n48778), .I0(n1837), .I1(n1460), .CO(n48779));
    SB_LUT4 add_2747_6_lut (.I0(GND_net), .I1(n1838), .I2(n1011), .I3(n48777), 
            .O(n8028[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_6 (.CI(n48777), .I0(n1838), .I1(n1011), .CO(n48778));
    SB_LUT4 add_2747_5_lut (.I0(GND_net), .I1(n1839), .I2(n856), .I3(n48776), 
            .O(n8028[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_37_LessThan_765_i42_3_lut (.I0(n40_adj_5111), .I1(baudrate[4]), 
            .I2(n43_adj_5118), .I3(GND_net), .O(n42_adj_5119));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i42_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2747_5 (.CI(n48776), .I0(n1839), .I1(n856), .CO(n48777));
    SB_LUT4 add_2747_4_lut (.I0(GND_net), .I1(n1840), .I2(n698), .I3(n48775), 
            .O(n8028[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_4 (.CI(n48775), .I0(n1840), .I1(n698), .CO(n48776));
    SB_LUT4 add_2747_3_lut (.I0(GND_net), .I1(n1841), .I2(n858), .I3(n48774), 
            .O(n8028[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2747_3 (.CI(n48774), .I0(n1841), .I1(n858), .CO(n48775));
    SB_LUT4 add_2747_2_lut (.I0(n56602), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n58474)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2747_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2747_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n48774));
    SB_LUT4 i48735_4_lut (.I0(n42_adj_5119), .I1(n38_adj_5117), .I2(n43_adj_5118), 
            .I3(n63357), .O(n65797));   // verilog/uart_rx.v(119[33:55])
    defparam i48735_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48736_3_lut (.I0(n65797), .I1(baudrate[5]), .I2(n1112), .I3(GND_net), 
            .O(n65798));   // verilog/uart_rx.v(119[33:55])
    defparam i48736_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_2753_7 (.CI(n48977), .I0(n2608), .I1(n1460), .CO(n48978));
    SB_LUT4 add_2753_6_lut (.I0(GND_net), .I1(n2609), .I2(n1011), .I3(n48976), 
            .O(n8184[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_6 (.CI(n48976), .I0(n2609), .I1(n1011), .CO(n48977));
    SB_LUT4 add_2753_5_lut (.I0(GND_net), .I1(n2610), .I2(n856), .I3(n48975), 
            .O(n8184[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_5 (.CI(n48975), .I0(n2610), .I1(n856), .CO(n48976));
    SB_LUT4 add_2753_4_lut (.I0(GND_net), .I1(n2611), .I2(n698), .I3(n48974), 
            .O(n8184[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_4 (.CI(n48974), .I0(n2611), .I1(n698), .CO(n48975));
    SB_LUT4 add_2753_3_lut (.I0(GND_net), .I1(n2612), .I2(n858), .I3(n48973), 
            .O(n8184[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2753_3 (.CI(n48973), .I0(n2612), .I1(n858), .CO(n48974));
    SB_LUT4 add_2753_2_lut (.I0(n56581), .I1(GND_net), .I2(n538), .I3(VCC_net), 
            .O(n58482)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2753_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2753_2 (.CI(VCC_net), .I0(GND_net), .I1(n538), .CO(n48973));
    SB_LUT4 i1_2_lut_4_lut_adj_1012 (.I0(n65996), .I1(baudrate[7]), .I2(n1261), 
            .I3(n58470), .O(n1415));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1012.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_LessThan_866_i36_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1267), .I3(GND_net), .O(n36_adj_5120));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i36_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2746_11_lut (.I0(GND_net), .I1(n1693), .I2(n2013), .I3(n48717), 
            .O(n8002[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2746_10_lut (.I0(GND_net), .I1(n1694), .I2(n1879), .I3(n48716), 
            .O(n8002[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_10 (.CI(n48716), .I0(n1694), .I1(n1879), .CO(n48717));
    SB_LUT4 add_2746_9_lut (.I0(GND_net), .I1(n1695), .I2(n1742), .I3(n48715), 
            .O(n8002[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_9 (.CI(n48715), .I0(n1695), .I1(n1742), .CO(n48716));
    SB_LUT4 add_2746_8_lut (.I0(GND_net), .I1(n1696), .I2(n1602), .I3(n48714), 
            .O(n8002[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_8 (.CI(n48714), .I0(n1696), .I1(n1602), .CO(n48715));
    SB_LUT4 add_2752_18_lut (.I0(GND_net), .I1(n2476), .I2(n2754), .I3(n48962), 
            .O(n8158[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2746_7_lut (.I0(GND_net), .I1(n1697), .I2(n1459), .I3(n48713), 
            .O(n8002[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_7 (.CI(n48713), .I0(n1697), .I1(n1459), .CO(n48714));
    SB_LUT4 add_2752_17_lut (.I0(GND_net), .I1(n2477), .I2(n2638), .I3(n48961), 
            .O(n8158[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2746_6_lut (.I0(GND_net), .I1(n1698), .I2(n1460), .I3(n48712), 
            .O(n8002[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_6 (.CI(n48712), .I0(n1698), .I1(n1460), .CO(n48713));
    SB_LUT4 add_2746_5_lut (.I0(GND_net), .I1(n1699), .I2(n1011), .I3(n48711), 
            .O(n8002[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_5 (.CI(n48711), .I0(n1699), .I1(n1011), .CO(n48712));
    SB_LUT4 add_2746_4_lut (.I0(GND_net), .I1(n1700), .I2(n856), .I3(n48710), 
            .O(n8002[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_4 (.CI(n48710), .I0(n1700), .I1(n856), .CO(n48711));
    SB_LUT4 add_2746_3_lut (.I0(GND_net), .I1(n1701), .I2(n698), .I3(n48709), 
            .O(n8002[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_17 (.CI(n48961), .I0(n2477), .I1(n2638), .CO(n48962));
    SB_CARRY add_2746_3 (.CI(n48709), .I0(n1701), .I1(n698), .CO(n48710));
    SB_LUT4 add_2746_2_lut (.I0(GND_net), .I1(n1702), .I2(n858), .I3(VCC_net), 
            .O(n8002[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2746_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2746_2 (.CI(VCC_net), .I0(n1702), .I1(n858), .CO(n48709));
    SB_LUT4 add_2752_16_lut (.I0(GND_net), .I1(n2478), .I2(n2519), .I3(n48960), 
            .O(n8158[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_16 (.CI(n48960), .I0(n2478), .I1(n2519), .CO(n48961));
    SB_LUT4 div_37_LessThan_866_i40_3_lut (.I0(n38_adj_5121), .I1(baudrate[4]), 
            .I2(n41_adj_5116), .I3(GND_net), .O(n40_adj_5122));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2752_15_lut (.I0(GND_net), .I1(n2479), .I2(n2397), .I3(n48959), 
            .O(n8158[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_15 (.CI(n48959), .I0(n2479), .I1(n2397), .CO(n48960));
    SB_LUT4 add_2752_14_lut (.I0(GND_net), .I1(n2480), .I2(n2272), .I3(n48958), 
            .O(n8158[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_14 (.CI(n48958), .I0(n2480), .I1(n2272), .CO(n48959));
    SB_LUT4 add_2752_13_lut (.I0(GND_net), .I1(n2481), .I2(n2144), .I3(n48957), 
            .O(n8158[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_13 (.CI(n48957), .I0(n2481), .I1(n2144), .CO(n48958));
    SB_LUT4 add_2752_12_lut (.I0(GND_net), .I1(n2482), .I2(n2013), .I3(n48956), 
            .O(n8158[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_12 (.CI(n48956), .I0(n2482), .I1(n2013), .CO(n48957));
    SB_LUT4 add_2752_11_lut (.I0(GND_net), .I1(n2483), .I2(n1879), .I3(n48955), 
            .O(n8158[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_11 (.CI(n48955), .I0(n2483), .I1(n1879), .CO(n48956));
    SB_LUT4 add_2752_10_lut (.I0(GND_net), .I1(n2484), .I2(n1742), .I3(n48954), 
            .O(n8158[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_10 (.CI(n48954), .I0(n2484), .I1(n1742), .CO(n48955));
    SB_LUT4 add_2752_9_lut (.I0(GND_net), .I1(n2485), .I2(n1602), .I3(n48953), 
            .O(n8158[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49041_4_lut (.I0(n40_adj_5122), .I1(n36_adj_5120), .I2(n41_adj_5116), 
            .I3(n63348), .O(n66103));   // verilog/uart_rx.v(119[33:55])
    defparam i49041_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2752_9 (.CI(n48953), .I0(n2485), .I1(n1602), .CO(n48954));
    SB_LUT4 i49042_3_lut (.I0(n66103), .I1(baudrate[5]), .I2(n1263), .I3(GND_net), 
            .O(n66104));   // verilog/uart_rx.v(119[33:55])
    defparam i49042_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_2752_8_lut (.I0(GND_net), .I1(n2486), .I2(n1459), .I3(n48952), 
            .O(n8158[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2752_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2752_8 (.CI(n48952), .I0(n2486), .I1(n1459), .CO(n48953));
    SB_LUT4 i48934_3_lut (.I0(n66104), .I1(baudrate[6]), .I2(n1262), .I3(GND_net), 
            .O(n65996));   // verilog/uart_rx.v(119[33:55])
    defparam i48934_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49328_2_lut_4_lut (.I0(n65996), .I1(baudrate[7]), .I2(n1261), 
            .I3(n59934), .O(n294[16]));   // verilog/uart_rx.v(119[33:55])
    defparam i49328_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1046_3_lut (.I0(n1415), .I1(n7950[16]), .I2(n294[15]), 
            .I3(GND_net), .O(n1559));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1141_3_lut (.I0(n1559), .I1(n7976[16]), .I2(n294[14]), 
            .I3(GND_net), .O(n1700));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1234_3_lut (.I0(n1700), .I1(n8002[16]), .I2(n294[13]), 
            .I3(GND_net), .O(n1838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_866_i38_3_lut_3_lut (.I0(n1265), .I1(baudrate[3]), 
            .I2(baudrate[2]), .I3(GND_net), .O(n38_adj_5121));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_866_i38_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 div_37_i1325_3_lut (.I0(n1838), .I1(n8028[16]), .I2(n294[12]), 
            .I3(GND_net), .O(n1973));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1414_3_lut (.I0(n1973), .I1(n8054[16]), .I2(n294[11]), 
            .I3(GND_net), .O(n2105));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1501_3_lut (.I0(n2105), .I1(n8080[16]), .I2(n294[10]), 
            .I3(GND_net), .O(n2234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46286_3_lut_4_lut (.I0(n1265), .I1(baudrate[3]), .I2(baudrate[2]), 
            .I3(n1266), .O(n63348));   // verilog/uart_rx.v(119[33:55])
    defparam i46286_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_4_lut_adj_1013 (.I0(n65798), .I1(baudrate[6]), .I2(n1111), 
            .I3(n58468), .O(n1267));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1013.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_LessThan_965_i45_2_lut (.I0(n1409), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_5123));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i39563_1_lut (.I0(n25202), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56577));
    defparam i39563_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i47008_3_lut (.I0(n962), .I1(baudrate[1]), .I2(n294[18]), 
            .I3(GND_net), .O(n1115));
    defparam i47008_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 div_37_i847_3_lut (.I0(n1115), .I1(n7898[19]), .I2(n294[17]), 
            .I3(GND_net), .O(n1265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_765_i43_2_lut (.I0(n1113), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5118));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_765_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i31_2_lut (.I0(n1974), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5124));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i29_2_lut (.I0(n1975), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5125));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i33_2_lut (.I0(n1973), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5126));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i35_2_lut (.I0(n1972), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5127));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i39_2_lut (.I0(n1970), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5128));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i37_2_lut (.I0(n1971), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5129));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i39_2_lut (.I0(n1697), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5130));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i41_2_lut (.I0(n1696), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5131));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i37_2_lut (.I0(n1698), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5132));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1157_i43_2_lut (.I0(n1695), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5133));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i31_2_lut (.I0(n2106), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5134));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i29_2_lut (.I0(n2107), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5135));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i33_2_lut (.I0(n2105), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5136));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i35_2_lut (.I0(n2104), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5137));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i39_2_lut (.I0(n2102), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5138));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1430_i37_2_lut (.I0(n2103), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i946_3_lut (.I0(n1265), .I1(n7924[19]), .I2(n294[16]), 
            .I3(GND_net), .O(n1412));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1430_i41_2_lut (.I0(n2101), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1014 (.I0(n2867), .I1(n59020), .I2(n698), .I3(n38422), 
            .O(n58400));
    defparam i1_4_lut_adj_1014.LUT_INIT = 16'h2000;
    SB_LUT4 i1_4_lut_adj_1015 (.I0(n59926), .I1(n58400), .I2(n25199), 
            .I3(n59886), .O(n57547));
    defparam i1_4_lut_adj_1015.LUT_INIT = 16'h0004;
    SB_LUT4 i1_4_lut_adj_1016 (.I0(baudrate[23]), .I1(baudrate[27]), .I2(baudrate[25]), 
            .I3(n38424), .O(n58748));
    defparam i1_4_lut_adj_1016.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1017 (.I0(n58748), .I1(baudrate[29]), .I2(baudrate[16]), 
            .I3(baudrate[28]), .O(n58766));
    defparam i1_4_lut_adj_1017.LUT_INIT = 16'h0002;
    SB_LUT4 i42913_4_lut (.I0(n59896), .I1(n59886), .I2(n59888), .I3(n59810), 
            .O(n59966));
    defparam i42913_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_965_i39_2_lut (.I0(n1412), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5139));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1018 (.I0(n59954), .I1(n59966), .I2(n56344), 
            .I3(n58766), .O(n57124));
    defparam i1_4_lut_adj_1018.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_adj_1019 (.I0(baudrate[3]), .I1(baudrate[4]), .I2(GND_net), 
            .I3(GND_net), .O(n59020));
    defparam i1_2_lut_adj_1019.LUT_INIT = 16'heeee;
    SB_LUT4 i22683_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n38424));
    defparam i22683_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22681_2_lut (.I0(baudrate[1]), .I1(baudrate[0]), .I2(GND_net), 
            .I3(GND_net), .O(n38422));
    defparam i22681_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_965_i41_2_lut (.I0(n1411), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5140));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5818_4_lut (.I0(n961), .I1(baudrate[2]), .I2(n962), .I3(baudrate[1]), 
            .O(n21323));   // verilog/uart_rx.v(119[33:55])
    defparam i5818_4_lut.LUT_INIT = 16'ha2aa;
    SB_LUT4 div_37_LessThan_1517_i29_2_lut (.I0(n2236), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5068));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i31_2_lut (.I0(n2235), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5073));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i27_2_lut (.I0(n2237), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5069));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i35_2_lut (.I0(n2233), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5071));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i25_2_lut (.I0(n2238), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5070));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i37_2_lut (.I0(n2232), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5078));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i39_2_lut (.I0(n2231), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5080));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i41_2_lut (.I0(n2230), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5081));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1517_i33_2_lut (.I0(n2234), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5072));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49267_2_lut_4_lut (.I0(n65798), .I1(baudrate[6]), .I2(n1111), 
            .I3(n59936), .O(n294[17]));   // verilog/uart_rx.v(119[33:55])
    defparam i49267_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_965_i43_2_lut (.I0(n1410), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5141));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_965_i34_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1415), .I3(GND_net), .O(n34_adj_5142));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i34_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2159_1_lut (.I0(baudrate[16]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2754));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2159_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i48733_3_lut (.I0(n34_adj_5142), .I1(baudrate[5]), .I2(n41_adj_5140), 
            .I3(GND_net), .O(n65795));   // verilog/uart_rx.v(119[33:55])
    defparam i48733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2158_1_lut (.I0(baudrate[17]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2867));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2158_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i48734_3_lut (.I0(n65795), .I1(baudrate[6]), .I2(n43_adj_5141), 
            .I3(GND_net), .O(n65796));   // verilog/uart_rx.v(119[33:55])
    defparam i48734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2157_1_lut (.I0(baudrate[18]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2977));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2157_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2156_1_lut (.I0(baudrate[19]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3084));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2156_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i47228_4_lut (.I0(n43_adj_5141), .I1(n41_adj_5140), .I2(n39_adj_5139), 
            .I3(n63341), .O(n64290));
    defparam i47228_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_37_i2155_1_lut (.I0(baudrate[20]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2155_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_965_i38_3_lut (.I0(n36), .I1(baudrate[4]), .I2(n39_adj_5139), 
            .I3(GND_net), .O(n38_adj_5143));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_965_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2083_1_lut (.I0(baudrate[21]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3082));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2083_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2153_1_lut (.I0(baudrate[22]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2153_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i48477_3_lut (.I0(n65796), .I1(baudrate[7]), .I2(n45_adj_5123), 
            .I3(GND_net), .O(n44_adj_5144));   // verilog/uart_rx.v(119[33:55])
    defparam i48477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48079_4_lut (.I0(n44_adj_5144), .I1(n38_adj_5143), .I2(n45_adj_5123), 
            .I3(n64290), .O(n65141));   // verilog/uart_rx.v(119[33:55])
    defparam i48079_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48080_3_lut (.I0(n65141), .I1(baudrate[8]), .I2(n1408), .I3(GND_net), 
            .O(n48_adj_5145));   // verilog/uart_rx.v(119[33:55])
    defparam i48080_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1020 (.I0(n58472), .I1(n48_adj_5145), .I2(GND_net), 
            .I3(GND_net), .O(n1560));
    defparam i1_2_lut_adj_1020.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i1142_3_lut (.I0(n1560), .I1(n7976[15]), .I2(n294[14]), 
            .I3(GND_net), .O(n1701));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1235_3_lut (.I0(n1701), .I1(n8002[15]), .I2(n294[13]), 
            .I3(GND_net), .O(n1839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1326_3_lut (.I0(n1839), .I1(n8028[15]), .I2(n294[12]), 
            .I3(GND_net), .O(n1974));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1415_3_lut (.I0(n1974), .I1(n8054[15]), .I2(n294[11]), 
            .I3(GND_net), .O(n2106));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1502_3_lut (.I0(n2106), .I1(n8080[15]), .I2(n294[10]), 
            .I3(GND_net), .O(n2235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1587_3_lut (.I0(n2235), .I1(n8106[15]), .I2(n294[9]), 
            .I3(GND_net), .O(n2361));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1586_3_lut (.I0(n2234), .I1(n8106[16]), .I2(n294[9]), 
            .I3(GND_net), .O(n2360));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i31_2_lut (.I0(n2361), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5089));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i33_2_lut (.I0(n2360), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5088));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i42855_2_lut (.I0(baudrate[12]), .I1(n59876), .I2(GND_net), 
            .I3(GND_net), .O(n59908));
    defparam i42855_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1021 (.I0(baudrate[27]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n59202));
    defparam i1_2_lut_adj_1021.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1022 (.I0(baudrate[25]), .I1(baudrate[29]), .I2(GND_net), 
            .I3(GND_net), .O(n59394));
    defparam i1_2_lut_adj_1022.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1023 (.I0(baudrate[24]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n59396));
    defparam i1_2_lut_adj_1023.LUT_INIT = 16'heeee;
    SB_LUT4 i2314_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n479[2]));   // verilog/uart_rx.v(103[36:51])
    defparam i2314_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 div_37_LessThan_1430_i28_3_lut_3_lut (.I0(baudrate[3]), .I1(baudrate[4]), 
            .I2(n2107), .I3(GND_net), .O(n28_adj_5146));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46167_2_lut_4_lut (.I0(n2102), .I1(baudrate[9]), .I2(n2106), 
            .I3(baudrate[5]), .O(n63229));
    defparam i46167_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1430_i30_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[9]), 
            .I2(n2102), .I3(GND_net), .O(n30_adj_5147));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_4_lut_adj_1024 (.I0(baudrate[20]), .I1(baudrate[21]), 
            .I2(baudrate[22]), .I3(baudrate[23]), .O(n59308));
    defparam i1_2_lut_4_lut_adj_1024.LUT_INIT = 16'hfffe;
    SB_LUT4 i39281_2_lut (.I0(\r_SM_Main_2__N_3446[1] ), .I1(r_SM_Main[1]), 
            .I2(GND_net), .I3(GND_net), .O(n56281));
    defparam i39281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1025 (.I0(\o_Rx_DV_N_3488[12] ), .I1(n5225), .I2(\o_Rx_DV_N_3488[8] ), 
            .I3(n55184), .O(n58586));
    defparam i1_4_lut_adj_1025.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1026 (.I0(n59394), .I1(n59212), .I2(n59294), 
            .I3(n59202), .O(n25211));
    defparam i1_4_lut_adj_1026.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1027 (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(baudrate[18]), .I3(baudrate[19]), .O(n59310));
    defparam i1_2_lut_4_lut_adj_1027.LUT_INIT = 16'hfffe;
    SB_LUT4 i22689_rep_10_2_lut (.I0(baudrate[0]), .I1(n294[19]), .I2(GND_net), 
            .I3(GND_net), .O(n56622));   // verilog/uart_rx.v(119[33:55])
    defparam i22689_rep_10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1028 (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), 
            .I2(\o_Rx_DV_N_3488[2] ), .I3(\o_Rx_DV_N_3488[1] ), .O(n59190));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1028.LUT_INIT = 16'h7bde;
    SB_LUT4 equal_271_i3_2_lut (.I0(r_Clock_Count[2]), .I1(\o_Rx_DV_N_3488[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_5148));   // verilog/uart_rx.v(69[17:62])
    defparam equal_271_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1029 (.I0(r_Clock_Count[3]), .I1(n3_adj_5148), 
            .I2(\o_Rx_DV_N_3488[4] ), .I3(n59190), .O(n59194));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1029.LUT_INIT = 16'hffde;
    SB_LUT4 i1_4_lut_adj_1030 (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n58586), .O(n58592));
    defparam i1_4_lut_adj_1030.LUT_INIT = 16'h0100;
    SB_LUT4 div_37_LessThan_662_i42_4_lut (.I0(n56622), .I1(baudrate[2]), 
            .I2(n961), .I3(baudrate[1]), .O(n42_adj_5149));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_662_i42_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 equal_271_i5_2_lut (.I0(r_Clock_Count[4]), .I1(\o_Rx_DV_N_3488[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/uart_rx.v(69[17:62])
    defparam equal_271_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1031 (.I0(r_Clock_Count[5]), .I1(n5), .I2(\o_Rx_DV_N_3488[6] ), 
            .I3(n59194), .O(n59198));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1031.LUT_INIT = 16'hffde;
    SB_LUT4 equal_271_i8_2_lut (.I0(r_Clock_Count[7]), .I1(\o_Rx_DV_N_3488[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/uart_rx.v(69[17:62])
    defparam equal_271_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1032 (.I0(r_Clock_Count[6]), .I1(n8), .I2(n59198), 
            .I3(\o_Rx_DV_N_3488[7] ), .O(n55210));   // verilog/uart_rx.v(69[17:62])
    defparam i1_4_lut_adj_1032.LUT_INIT = 16'hfdfe;
    SB_LUT4 i1_4_lut_adj_1033 (.I0(n58592), .I1(n6), .I2(r_SM_Main[1]), 
            .I3(n27), .O(n28373));   // verilog/uart_rx.v(50[10] 145[8])
    defparam i1_4_lut_adj_1033.LUT_INIT = 16'h0323;
    SB_LUT4 i48737_3_lut (.I0(n42_adj_5149), .I1(baudrate[3]), .I2(n960), 
            .I3(GND_net), .O(n65799));   // verilog/uart_rx.v(119[33:55])
    defparam i48737_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48738_3_lut (.I0(n65799), .I1(baudrate[4]), .I2(n959), .I3(GND_net), 
            .O(n65800));   // verilog/uart_rx.v(119[33:55])
    defparam i48738_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47039_2_lut (.I0(n55210), .I1(r_Rx_Data), .I2(GND_net), .I3(GND_net), 
            .O(n63003));
    defparam i47039_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i48467_3_lut (.I0(n65800), .I1(baudrate[5]), .I2(n56323), 
            .I3(GND_net), .O(n48_adj_5150));   // verilog/uart_rx.v(119[33:55])
    defparam i48467_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n55184));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i47034_4_lut (.I0(n63003), .I1(n29), .I2(n23), .I3(\o_Rx_DV_N_3488[12] ), 
            .O(n63000));
    defparam i47034_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i46186_4_lut (.I0(n63000), .I1(r_SM_Main[0]), .I2(n27), .I3(\o_Rx_DV_N_3488[24] ), 
            .O(n62997));
    defparam i46186_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i49325_4_lut (.I0(r_SM_Main[2]), .I1(n62997), .I2(\r_SM_Main_2__N_3446[1] ), 
            .I3(r_SM_Main[1]), .O(n28645));
    defparam i49325_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i1_4_lut_adj_1034 (.I0(n55210), .I1(r_SM_Main[1]), .I2(r_Rx_Data), 
            .I3(r_SM_Main[0]), .O(n58548));
    defparam i1_4_lut_adj_1034.LUT_INIT = 16'h1000;
    SB_LUT4 i1_4_lut_adj_1035 (.I0(n29), .I1(n23), .I2(\o_Rx_DV_N_3488[12] ), 
            .I3(n58548), .O(n58554));
    defparam i1_4_lut_adj_1035.LUT_INIT = 16'h0100;
    SB_LUT4 i42650_1_lut_2_lut (.I0(baudrate[17]), .I1(n25199), .I2(GND_net), 
            .I3(GND_net), .O(n56585));
    defparam i42650_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_4_lut_adj_1036 (.I0(n59240), .I1(n25211), .I2(n59282), 
            .I3(n59238), .O(n25163));
    defparam i1_4_lut_adj_1036.LUT_INIT = 16'hfffe;
    SB_LUT4 i49245_4_lut (.I0(r_SM_Main[2]), .I1(\o_Rx_DV_N_3488[24] ), 
            .I2(n27), .I3(n58554), .O(n27426));   // verilog/uart_rx.v(53[7] 144[14])
    defparam i49245_4_lut.LUT_INIT = 16'h5455;
    SB_LUT4 i1_3_lut_adj_1037 (.I0(n25163), .I1(n48_adj_5150), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1116));
    defparam i1_3_lut_adj_1037.LUT_INIT = 16'hefef;
    SB_LUT4 i42801_2_lut (.I0(\o_Rx_DV_N_3488[12] ), .I1(n55210), .I2(GND_net), 
            .I3(GND_net), .O(n59854));
    defparam i42801_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i42907_4_lut (.I0(\o_Rx_DV_N_3488[24] ), .I1(n29), .I2(n23), 
            .I3(n59854), .O(n59960));
    defparam i42907_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i2_4_lut (.I0(n58618), .I1(\r_SM_Main_2__N_3446[1] ), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n2));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i2_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i1_4_lut (.I0(r_Rx_Data), .I1(n59960), 
            .I2(r_SM_Main[0]), .I3(n27), .O(n10007));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 r_SM_Main_2__I_0_62_Mux_0_i3_3_lut (.I0(n10007), .I1(n2), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(53[7] 144[14])
    defparam r_SM_Main_2__I_0_62_Mux_0_i3_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i4209_2_lut_4_lut (.I0(n960), .I1(n9784), .I2(n21323), .I3(baudrate[3]), 
            .O(n44_adj_5151));   // verilog/uart_rx.v(119[33:55])
    defparam i4209_2_lut_4_lut.LUT_INIT = 16'ha8fe;
    SB_LUT4 div_37_i848_3_lut (.I0(n1116), .I1(n7898[18]), .I2(n294[17]), 
            .I3(GND_net), .O(n1266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2307_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n479[1]));   // verilog/uart_rx.v(103[36:51])
    defparam i2307_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i42843_3_lut_4_lut (.I0(baudrate[30]), .I1(baudrate[31]), .I2(baudrate[26]), 
            .I3(baudrate[24]), .O(n59896));
    defparam i42843_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i947_3_lut (.I0(n1266), .I1(n7924[18]), .I2(n294[16]), 
            .I3(GND_net), .O(n1413));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4031_2_lut_4_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n42_adj_5064));   // verilog/uart_rx.v(119[33:55])
    defparam i4031_2_lut_4_lut_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_3_lut_4_lut (.I0(baudrate[30]), .I1(baudrate[31]), .I2(baudrate[27]), 
            .I3(baudrate[24]), .O(n58422));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1038 (.I0(n66095), .I1(baudrate[11]), .I2(n1831), 
            .I3(n58474), .O(n1977));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1038.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_i1044_3_lut (.I0(n1413), .I1(n7950[18]), .I2(n294[15]), 
            .I3(GND_net), .O(n1557));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4202_2_lut_3_lut_4_lut (.I0(n21323), .I1(baudrate[2]), .I2(n962), 
            .I3(baudrate[1]), .O(n42_adj_5065));   // verilog/uart_rx.v(119[33:55])
    defparam i4202_2_lut_3_lut_4_lut.LUT_INIT = 16'hbabb;
    SB_LUT4 div_37_LessThan_2210_i39_4_lut (.I0(n3155), .I1(baudrate[19]), 
            .I2(n8314[19]), .I3(n294[1]), .O(n39_adj_5152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i39_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i41_4_lut (.I0(n3154), .I1(baudrate[20]), 
            .I2(n8314[20]), .I3(n294[1]), .O(n41_adj_5153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i41_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i33_4_lut (.I0(n3158), .I1(baudrate[16]), 
            .I2(n8314[16]), .I3(n294[1]), .O(n33_adj_5154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i33_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_1062_i43_2_lut (.I0(n1554), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2210_i35_4_lut (.I0(n3157), .I1(baudrate[17]), 
            .I2(n8314[17]), .I3(n294[1]), .O(n35_adj_5156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i35_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i42819_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[29]), .I3(baudrate[24]), .O(n59872));
    defparam i42819_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(baudrate[28]), .I1(baudrate[26]), 
            .I2(baudrate[24]), .I3(baudrate[31]), .O(n59212));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2210_i37_4_lut (.I0(n3156), .I1(baudrate[18]), 
            .I2(n8314[18]), .I3(n294[1]), .O(n37_adj_5157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i37_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i29_4_lut (.I0(n3160), .I1(baudrate[14]), 
            .I2(n8314[14]), .I3(n294[1]), .O(n29_adj_5158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i29_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_1062_i39_2_lut (.I0(n1556), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2210_i31_4_lut (.I0(n3159), .I1(baudrate[15]), 
            .I2(n8314[15]), .I3(n294[1]), .O(n31_adj_5160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i31_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i1_2_lut_4_lut_adj_1039 (.I0(baudrate[30]), .I1(baudrate[25]), 
            .I2(baudrate[31]), .I3(baudrate[26]), .O(n59270));
    defparam i1_2_lut_4_lut_adj_1039.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2210_i23_4_lut (.I0(n3163), .I1(baudrate[11]), 
            .I2(n8314[11]), .I3(n294[1]), .O(n23_adj_5161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i23_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i39567_1_lut (.I0(n25199), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56581));
    defparam i39567_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1062_i41_2_lut (.I0(n1555), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2210_i25_4_lut (.I0(n3162), .I1(baudrate[12]), 
            .I2(n8314[12]), .I3(n294[1]), .O(n25_adj_5163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i25_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_1062_i37_2_lut (.I0(n1557), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2210_i7_4_lut (.I0(n3171), .I1(baudrate[3]), 
            .I2(n8314[3]), .I3(n294[1]), .O(n7));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i7_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i49361_2_lut_4_lut (.I0(n66095), .I1(baudrate[11]), .I2(n1831), 
            .I3(n59908), .O(n294[12]));   // verilog/uart_rx.v(119[33:55])
    defparam i49361_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_2210_i45_4_lut (.I0(n3152), .I1(baudrate[22]), 
            .I2(n8314[22]), .I3(n294[1]), .O(n45_adj_5165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i45_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i43_4_lut (.I0(n3153), .I1(baudrate[21]), 
            .I2(n8314[21]), .I3(n294[1]), .O(n43_adj_5166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i43_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i9_4_lut (.I0(n3170), .I1(baudrate[4]), 
            .I2(n8314[4]), .I3(n294[1]), .O(n9));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i9_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i17_4_lut (.I0(n3166), .I1(baudrate[8]), 
            .I2(n8314[8]), .I3(n294[1]), .O(n17_adj_5167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i17_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i19_4_lut (.I0(n3165), .I1(baudrate[9]), 
            .I2(n8314[9]), .I3(n294[1]), .O(n19_adj_5168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i19_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i21_4_lut (.I0(n3164), .I1(baudrate[10]), 
            .I2(n8314[10]), .I3(n294[1]), .O(n21_adj_5169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i21_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i11_4_lut (.I0(n3169), .I1(baudrate[5]), 
            .I2(n8314[5]), .I3(n294[1]), .O(n11));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i11_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i13_4_lut (.I0(n3168), .I1(baudrate[6]), 
            .I2(n8314[6]), .I3(n294[1]), .O(n13));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i13_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i15_4_lut (.I0(n3167), .I1(baudrate[7]), 
            .I2(n8314[7]), .I3(n294[1]), .O(n15));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i15_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 div_37_LessThan_2210_i27_4_lut (.I0(n3161), .I1(baudrate[13]), 
            .I2(n8314[13]), .I3(n294[1]), .O(n27_adj_5170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i27_4_lut.LUT_INIT = 16'h3c66;
    SB_LUT4 i46619_4_lut (.I0(n27_adj_5170), .I1(n15), .I2(n13), .I3(n11), 
            .O(n63681));
    defparam i46619_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46639_4_lut (.I0(n21_adj_5169), .I1(n19_adj_5168), .I2(n17_adj_5167), 
            .I3(n9), .O(n63701));
    defparam i46639_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2210_i16_3_lut (.I0(baudrate[9]), .I1(baudrate[21]), 
            .I2(n43_adj_5166), .I3(GND_net), .O(n16_adj_5171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46591_2_lut (.I0(n43_adj_5166), .I1(n19_adj_5168), .I2(GND_net), 
            .I3(GND_net), .O(n63653));
    defparam i46591_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2210_i8_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n17_adj_5167), .I3(GND_net), .O(n8_adj_5172));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4036_2_lut_3_lut_4_lut_4_lut (.I0(baudrate[2]), .I1(n805), 
            .I2(baudrate[1]), .I3(baudrate[0]), .O(n9620));   // verilog/uart_rx.v(119[33:55])
    defparam i4036_2_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'h0445;
    SB_LUT4 div_37_LessThan_2210_i24_3_lut (.I0(n16_adj_5171), .I1(baudrate[22]), 
            .I2(n45_adj_5165), .I3(GND_net), .O(n24_adj_5173));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2208_3_lut (.I0(n3172), .I1(n8314[2]), .I2(n294[1]), 
            .I3(GND_net), .O(n3274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46660_3_lut (.I0(n7), .I1(n3274), .I2(baudrate[2]), .I3(GND_net), 
            .O(n63722));
    defparam i46660_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 i47626_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n63722), 
            .O(n64688));
    defparam i47626_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i48731_3_lut (.I0(n32_adj_5174), .I1(baudrate[5]), .I2(n39_adj_5159), 
            .I3(GND_net), .O(n65793));   // verilog/uart_rx.v(119[33:55])
    defparam i48731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47618_4_lut (.I0(n19_adj_5168), .I1(n17_adj_5167), .I2(n15), 
            .I3(n64688), .O(n64680));
    defparam i47618_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i48732_3_lut (.I0(n65793), .I1(baudrate[6]), .I2(n41_adj_5162), 
            .I3(GND_net), .O(n65794));   // verilog/uart_rx.v(119[33:55])
    defparam i48732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48833_4_lut (.I0(n25_adj_5163), .I1(n23_adj_5161), .I2(n21_adj_5169), 
            .I3(n64680), .O(n65895));
    defparam i48833_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47220_4_lut (.I0(n41_adj_5162), .I1(n39_adj_5159), .I2(n37_adj_5164), 
            .I3(n63329), .O(n64282));
    defparam i47220_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i48167_4_lut (.I0(n31_adj_5160), .I1(n29_adj_5158), .I2(n27_adj_5170), 
            .I3(n65895), .O(n65229));
    defparam i48167_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_37_LessThan_1922_i14_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2843), .I3(GND_net), .O(n14_adj_5175));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49004_4_lut (.I0(n37_adj_5157), .I1(n35_adj_5156), .I2(n33_adj_5154), 
            .I3(n65229), .O(n66066));
    defparam i49004_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i46865_2_lut_4_lut (.I0(n2838), .I1(baudrate[8]), .I2(n2842), 
            .I3(baudrate[4]), .O(n63927));
    defparam i46865_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i16_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2838), .I3(GND_net), .O(n16_adj_5176));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2210_i12_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n33_adj_5154), .I3(GND_net), .O(n12));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i4_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n58492), .I3(n48_adj_5177), .O(n4_c));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i4_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i48436_3_lut (.I0(n4_c), .I1(baudrate[13]), .I2(n27_adj_5170), 
            .I3(GND_net), .O(n65498));   // verilog/uart_rx.v(119[33:55])
    defparam i48436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i18_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2840), .I3(GND_net), .O(n18_adj_5178));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48437_3_lut (.I0(n65498), .I1(baudrate[14]), .I2(n29_adj_5158), 
            .I3(GND_net), .O(n65499));   // verilog/uart_rx.v(119[33:55])
    defparam i48437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48081_3_lut (.I0(n34_adj_5106), .I1(baudrate[4]), .I2(n37_adj_5164), 
            .I3(GND_net), .O(n65143));   // verilog/uart_rx.v(119[33:55])
    defparam i48081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46826_2_lut_4_lut (.I0(n2830), .I1(baudrate[16]), .I2(n2839), 
            .I3(baudrate[7]), .O(n63888));
    defparam i46826_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1922_i20_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2830), .I3(GND_net), .O(n20_adj_5179));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48479_3_lut (.I0(n65794), .I1(baudrate[7]), .I2(n43_adj_5155), 
            .I3(GND_net), .O(n65541));   // verilog/uart_rx.v(119[33:55])
    defparam i48479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48729_4_lut (.I0(n65541), .I1(n65143), .I2(n43_adj_5155), 
            .I3(n64282), .O(n65791));   // verilog/uart_rx.v(119[33:55])
    defparam i48729_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48730_3_lut (.I0(n65791), .I1(baudrate[8]), .I2(n1553), .I3(GND_net), 
            .O(n65792));   // verilog/uart_rx.v(119[33:55])
    defparam i48730_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46609_2_lut (.I0(n33_adj_5154), .I1(n15), .I2(GND_net), .I3(GND_net), 
            .O(n63671));
    defparam i46609_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_3_lut (.I0(r_SM_Main[0]), .I1(\o_Rx_DV_N_3488[24] ), .I2(n27), 
            .I3(GND_net), .O(n14_adj_5180));
    defparam i5_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i6_4_lut (.I0(n29), .I1(\o_Rx_DV_N_3488[12] ), .I2(n23), .I3(n5225), 
            .O(n15_adj_5181));
    defparam i6_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5181), .I1(\o_Rx_DV_N_3488[8] ), .I2(n14_adj_5180), 
            .I3(n55436), .O(n67140));
    defparam i8_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 div_37_LessThan_2210_i10_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n13), .I3(GND_net), .O(n10));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48481_3_lut (.I0(n65792), .I1(baudrate[9]), .I2(n1552), .I3(GND_net), 
            .O(n48_adj_5182));   // verilog/uart_rx.v(119[33:55])
    defparam i48481_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1341_i28_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1975), .I3(GND_net), .O(n28_adj_5183));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2210_i30_3_lut (.I0(n12), .I1(baudrate[17]), 
            .I2(n35_adj_5156), .I3(GND_net), .O(n30_adj_5184));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46613_4_lut (.I0(n33_adj_5154), .I1(n31_adj_5160), .I2(n29_adj_5158), 
            .I3(n63681), .O(n63675));
    defparam i46613_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46184_2_lut_4_lut (.I0(n1970), .I1(baudrate[8]), .I2(n1974), 
            .I3(baudrate[4]), .O(n63246));
    defparam i46184_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i48943_4_lut (.I0(n30_adj_5184), .I1(n10), .I2(n35_adj_5156), 
            .I3(n63671), .O(n66005));   // verilog/uart_rx.v(119[33:55])
    defparam i48943_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_LessThan_1341_i30_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1970), .I3(GND_net), .O(n30_adj_5185));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47465_3_lut (.I0(n65499), .I1(baudrate[15]), .I2(n31_adj_5160), 
            .I3(GND_net), .O(n64527));   // verilog/uart_rx.v(119[33:55])
    defparam i47465_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49134_4_lut (.I0(n64527), .I1(n66005), .I2(n35_adj_5156), 
            .I3(n63675), .O(n66196));   // verilog/uart_rx.v(119[33:55])
    defparam i49134_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49135_3_lut (.I0(n66196), .I1(baudrate[18]), .I2(n37_adj_5157), 
            .I3(GND_net), .O(n66197));   // verilog/uart_rx.v(119[33:55])
    defparam i49135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2210_i6_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n7), .I3(GND_net), .O(n6_adj_5186));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2210_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48438_3_lut (.I0(n6_adj_5186), .I1(baudrate[10]), .I2(n21_adj_5169), 
            .I3(GND_net), .O(n65500));   // verilog/uart_rx.v(119[33:55])
    defparam i48438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48439_3_lut (.I0(n65500), .I1(baudrate[11]), .I2(n23_adj_5161), 
            .I3(GND_net), .O(n65501));   // verilog/uart_rx.v(119[33:55])
    defparam i48439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46593_4_lut (.I0(n43_adj_5166), .I1(n25_adj_5163), .I2(n23_adj_5161), 
            .I3(n63701), .O(n63655));
    defparam i46593_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48525_4_lut (.I0(n24_adj_5173), .I1(n8_adj_5172), .I2(n45_adj_5165), 
            .I3(n63653), .O(n65587));   // verilog/uart_rx.v(119[33:55])
    defparam i48525_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47463_3_lut (.I0(n65501), .I1(baudrate[12]), .I2(n25_adj_5163), 
            .I3(GND_net), .O(n64525));   // verilog/uart_rx.v(119[33:55])
    defparam i47463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49056_3_lut (.I0(n66197), .I1(baudrate[19]), .I2(n39_adj_5152), 
            .I3(GND_net), .O(n66118));   // verilog/uart_rx.v(119[33:55])
    defparam i49056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46595_4_lut (.I0(n43_adj_5166), .I1(n41_adj_5153), .I2(n39_adj_5152), 
            .I3(n66066), .O(n63657));
    defparam i46595_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48992_4_lut (.I0(n64525), .I1(n65587), .I2(n45_adj_5165), 
            .I3(n63655), .O(n66054));   // verilog/uart_rx.v(119[33:55])
    defparam i48992_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47471_3_lut (.I0(n66118), .I1(baudrate[20]), .I2(n41_adj_5153), 
            .I3(GND_net), .O(n64533));   // verilog/uart_rx.v(119[33:55])
    defparam i47471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i12_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2955), .I3(GND_net), .O(n12_adj_5187));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46804_2_lut_4_lut (.I0(n2950), .I1(baudrate[8]), .I2(n2954), 
            .I3(baudrate[4]), .O(n63866));
    defparam i46804_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1997_i14_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2950), .I3(GND_net), .O(n14_adj_5188));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1040 (.I0(baudrate[25]), .I1(baudrate[31]), .I2(GND_net), 
            .I3(GND_net), .O(n58436));
    defparam i1_2_lut_adj_1040.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_i2187_3_lut (.I0(n3151), .I1(n8314[23]), .I2(n294[1]), 
            .I3(GND_net), .O(n3253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_349_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(98[17:39])
    defparam equal_349_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i48994_4_lut (.I0(n64533), .I1(n66054), .I2(n45_adj_5165), 
            .I3(n63657), .O(n66056));   // verilog/uart_rx.v(119[33:55])
    defparam i48994_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1041 (.I0(n59392), .I1(n59252), .I2(n58436), 
            .I3(n59250), .O(n58444));
    defparam i1_4_lut_adj_1041.LUT_INIT = 16'hfffe;
    SB_LUT4 i49349_4_lut (.I0(n58444), .I1(n66056), .I2(baudrate[23]), 
            .I3(n3253), .O(n57452));   // verilog/uart_rx.v(119[33:55])
    defparam i49349_4_lut.LUT_INIT = 16'h1501;
    SB_LUT4 div_37_LessThan_1997_i16_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2952), .I3(GND_net), .O(n16_adj_5190));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46772_2_lut_4_lut (.I0(n2942), .I1(baudrate[16]), .I2(n2951), 
            .I3(baudrate[7]), .O(n63834));
    defparam i46772_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i42882_1_lut (.I0(n59934), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n56615));
    defparam i42882_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1997_i18_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2942), .I3(GND_net), .O(n18_adj_5191));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2118_3_lut (.I0(n3046), .I1(n8288[23]), .I2(n294[2]), 
            .I3(GND_net), .O(n3151));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2119_3_lut (.I0(n3047), .I1(n8288[22]), .I2(n294[2]), 
            .I3(GND_net), .O(n3152));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1236_3_lut (.I0(n1702), .I1(n8002[14]), .I2(n294[13]), 
            .I3(GND_net), .O(n1840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2120_3_lut (.I0(n3048), .I1(n8288[21]), .I2(n294[2]), 
            .I3(GND_net), .O(n3153));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2121_3_lut (.I0(n3049), .I1(n8288[20]), .I2(n294[2]), 
            .I3(GND_net), .O(n3154));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2122_3_lut (.I0(n3050), .I1(n8288[19]), .I2(n294[2]), 
            .I3(GND_net), .O(n3155));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2125_3_lut (.I0(n3053), .I1(n8288[16]), .I2(n294[2]), 
            .I3(GND_net), .O(n3158));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i33_2_lut (.I0(n3158), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5192));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2126_3_lut (.I0(n3054), .I1(n8288[15]), .I2(n294[2]), 
            .I3(GND_net), .O(n3159));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i31_2_lut (.I0(n3159), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5193));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2123_3_lut (.I0(n3051), .I1(n8288[18]), .I2(n294[2]), 
            .I3(GND_net), .O(n3156));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i37_2_lut (.I0(n3156), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5194));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2124_3_lut (.I0(n3052), .I1(n8288[17]), .I2(n294[2]), 
            .I3(GND_net), .O(n3157));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i35_2_lut (.I0(n3157), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5195));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2130_3_lut (.I0(n3058), .I1(n8288[11]), .I2(n294[2]), 
            .I3(GND_net), .O(n3163));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2131_3_lut (.I0(n3059), .I1(n8288[10]), .I2(n294[2]), 
            .I3(GND_net), .O(n3164));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i21_2_lut (.I0(n3164), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5196));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i23_2_lut (.I0(n3163), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5197));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2137_3_lut (.I0(n3065), .I1(n8288[4]), .I2(n294[2]), 
            .I3(GND_net), .O(n3170));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1327_3_lut (.I0(n1840), .I1(n8028[14]), .I2(n294[12]), 
            .I3(GND_net), .O(n1975));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2138_3_lut (.I0(n3066), .I1(n8288[3]), .I2(n294[2]), 
            .I3(GND_net), .O(n3171));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i9_2_lut (.I0(n3170), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_5198));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2132_3_lut (.I0(n3060), .I1(n8288[9]), .I2(n294[2]), 
            .I3(GND_net), .O(n3165));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2136_3_lut (.I0(n3064), .I1(n8288[5]), .I2(n294[2]), 
            .I3(GND_net), .O(n3169));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i11_2_lut (.I0(n3169), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5199));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i42658_1_lut_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n25199), .I3(baudrate[15]), .O(n56593));
    defparam i42658_1_lut_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i49440_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n25199), .I3(n48_adj_5108), .O(n294[8]));
    defparam i49440_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 div_37_LessThan_2141_i19_2_lut (.I0(n3165), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5200));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2128_3_lut (.I0(n3056), .I1(n8288[13]), .I2(n294[2]), 
            .I3(GND_net), .O(n3161));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2129_3_lut (.I0(n3057), .I1(n8288[12]), .I2(n294[2]), 
            .I3(GND_net), .O(n3162));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i25_2_lut (.I0(n3162), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5201));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i27_2_lut (.I0(n3161), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5202));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i42656_1_lut_2_lut_3_lut (.I0(baudrate[16]), .I1(baudrate[17]), 
            .I2(n25199), .I3(GND_net), .O(n56589));
    defparam i42656_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 div_37_i2127_3_lut (.I0(n3055), .I1(n8288[14]), .I2(n294[2]), 
            .I3(GND_net), .O(n3160));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2133_3_lut (.I0(n3061), .I1(n8288[8]), .I2(n294[2]), 
            .I3(GND_net), .O(n3166));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2134_3_lut (.I0(n3062), .I1(n8288[7]), .I2(n294[2]), 
            .I3(GND_net), .O(n3167));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i10_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3064), .I3(GND_net), .O(n10_adj_5203));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2135_3_lut (.I0(n3063), .I1(n8288[6]), .I2(n294[2]), 
            .I3(GND_net), .O(n3168));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i14_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3061), .I3(GND_net), .O(n14_adj_5204));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i13_2_lut (.I0(n3168), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5205));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i15_2_lut (.I0(n3167), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5206));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2141_i17_2_lut (.I0(n3166), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5207));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46980_2_lut_3_lut (.I0(n25229), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n63061));   // verilog/uart_rx.v(119[33:55])
    defparam i46980_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 div_37_i1416_3_lut (.I0(n1975), .I1(n8054[14]), .I2(n294[11]), 
            .I3(GND_net), .O(n2107));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46717_2_lut_4_lut (.I0(n3051), .I1(baudrate[16]), .I2(n3060), 
            .I3(baudrate[7]), .O(n63779));
    defparam i46717_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i1503_3_lut (.I0(n2107), .I1(n8080[14]), .I2(n294[10]), 
            .I3(GND_net), .O(n2236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i16_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3051), .I3(GND_net), .O(n16_adj_5208));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2141_i29_2_lut (.I0(n3160), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5209));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1588_3_lut (.I0(n2236), .I1(n8106[14]), .I2(n294[9]), 
            .I3(GND_net), .O(n2362));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1042 (.I0(baudrate[26]), .I1(baudrate[30]), .I2(GND_net), 
            .I3(GND_net), .O(n59392));
    defparam i1_2_lut_adj_1042.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1043 (.I0(n59396), .I1(n59398), .I2(n59250), 
            .I3(n59394), .O(n25214));
    defparam i1_4_lut_adj_1043.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2070_i12_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3059), .I3(GND_net), .O(n12_adj_5210));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46750_2_lut_4_lut (.I0(n3059), .I1(baudrate[8]), .I2(n3063), 
            .I3(baudrate[4]), .O(n63812));
    defparam i46750_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i46685_4_lut (.I0(n29_adj_5209), .I1(n17_adj_5207), .I2(n15_adj_5206), 
            .I3(n13_adj_5205), .O(n63747));
    defparam i46685_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47674_4_lut (.I0(n11_adj_5199), .I1(n9_adj_5198), .I2(n3171), 
            .I3(baudrate[2]), .O(n64736));
    defparam i47674_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i48209_4_lut (.I0(n17_adj_5207), .I1(n15_adj_5206), .I2(n13_adj_5205), 
            .I3(n64736), .O(n65271));
    defparam i48209_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48205_4_lut (.I0(n23_adj_5197), .I1(n21_adj_5196), .I2(n19_adj_5200), 
            .I3(n65271), .O(n65267));
    defparam i48205_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i46687_4_lut (.I0(n29_adj_5209), .I1(n27_adj_5202), .I2(n25_adj_5201), 
            .I3(n65267), .O(n63749));
    defparam i46687_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2141_i6_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3172), .I3(GND_net), .O(n6_adj_5211));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48448_3_lut (.I0(n6_adj_5211), .I1(baudrate[13]), .I2(n29_adj_5209), 
            .I3(GND_net), .O(n65510));   // verilog/uart_rx.v(119[33:55])
    defparam i48448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2141_i32_3_lut (.I0(n14_adj_5212), .I1(baudrate[17]), 
            .I2(n37_adj_5194), .I3(GND_net), .O(n32_adj_5213));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48449_3_lut (.I0(n65510), .I1(baudrate[14]), .I2(n31_adj_5193), 
            .I3(GND_net), .O(n65511));   // verilog/uart_rx.v(119[33:55])
    defparam i48449_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46679_4_lut (.I0(n35_adj_5195), .I1(n33_adj_5192), .I2(n31_adj_5193), 
            .I3(n63747), .O(n63741));
    defparam i46679_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48941_4_lut (.I0(n32_adj_5213), .I1(n12_adj_5214), .I2(n37_adj_5194), 
            .I3(n63735), .O(n66003));   // verilog/uart_rx.v(119[33:55])
    defparam i48941_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47451_3_lut (.I0(n65511), .I1(baudrate[15]), .I2(n33_adj_5192), 
            .I3(GND_net), .O(n64513));   // verilog/uart_rx.v(119[33:55])
    defparam i47451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48450_3_lut (.I0(n8_adj_5215), .I1(baudrate[10]), .I2(n23_adj_5197), 
            .I3(GND_net), .O(n65512));   // verilog/uart_rx.v(119[33:55])
    defparam i48450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1044 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(GND_net), 
            .I3(GND_net), .O(n55436));
    defparam i1_2_lut_adj_1044.LUT_INIT = 16'h2222;
    SB_LUT4 i48451_3_lut (.I0(n65512), .I1(baudrate[11]), .I2(n25_adj_5201), 
            .I3(GND_net), .O(n65513));   // verilog/uart_rx.v(119[33:55])
    defparam i48451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47660_4_lut (.I0(n25_adj_5201), .I1(n23_adj_5197), .I2(n21_adj_5196), 
            .I3(n63759), .O(n64722));
    defparam i47660_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i47013_4_lut (.I0(\o_Rx_DV_N_3488[8] ), .I1(\o_Rx_DV_N_3488[12] ), 
            .I2(n5225), .I3(n55436), .O(n62954));
    defparam i47013_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i47009_4_lut (.I0(n62954), .I1(\o_Rx_DV_N_3488[24] ), .I2(n29), 
            .I3(n23), .O(n62951));
    defparam i47009_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i48523_3_lut (.I0(n10_adj_5216), .I1(baudrate[9]), .I2(n21_adj_5196), 
            .I3(GND_net), .O(n65585));   // verilog/uart_rx.v(119[33:55])
    defparam i48523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_4_lut (.I0(r_SM_Main[1]), .I1(n62951), .I2(r_SM_Main[0]), 
            .I3(n27), .O(n27308));
    defparam i14_4_lut.LUT_INIT = 16'h05c5;
    SB_LUT4 i47449_3_lut (.I0(n65513), .I1(baudrate[12]), .I2(n27_adj_5202), 
            .I3(GND_net), .O(n64511));   // verilog/uart_rx.v(119[33:55])
    defparam i47449_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48617_4_lut (.I0(n35_adj_5195), .I1(n33_adj_5192), .I2(n31_adj_5193), 
            .I3(n63749), .O(n65679));
    defparam i48617_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i49132_4_lut (.I0(n64513), .I1(n66003), .I2(n37_adj_5194), 
            .I3(n63741), .O(n66194));   // verilog/uart_rx.v(119[33:55])
    defparam i49132_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48755_4_lut (.I0(n64511), .I1(n65585), .I2(n27_adj_5202), 
            .I3(n64722), .O(n65817));   // verilog/uart_rx.v(119[33:55])
    defparam i48755_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49187_4_lut (.I0(n65817), .I1(n66194), .I2(n37_adj_5194), 
            .I3(n65679), .O(n66249));   // verilog/uart_rx.v(119[33:55])
    defparam i49187_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49188_3_lut (.I0(n66249), .I1(baudrate[18]), .I2(n3155), 
            .I3(GND_net), .O(n66250));   // verilog/uart_rx.v(119[33:55])
    defparam i49188_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49178_3_lut (.I0(n66250), .I1(baudrate[19]), .I2(n3154), 
            .I3(GND_net), .O(n66240));   // verilog/uart_rx.v(119[33:55])
    defparam i49178_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48981_3_lut (.I0(n66240), .I1(baudrate[20]), .I2(n3153), 
            .I3(GND_net), .O(n66043));   // verilog/uart_rx.v(119[33:55])
    defparam i48981_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48982_3_lut (.I0(n66043), .I1(baudrate[21]), .I2(n3152), 
            .I3(GND_net), .O(n66044));   // verilog/uart_rx.v(119[33:55])
    defparam i48982_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i29_2_lut (.I0(n2362), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5090));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47461_3_lut (.I0(n66044), .I1(baudrate[22]), .I2(n3151), 
            .I3(GND_net), .O(n48_adj_5177));   // verilog/uart_rx.v(119[33:55])
    defparam i47461_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2047_3_lut (.I0(n2938), .I1(n8262[23]), .I2(n294[3]), 
            .I3(GND_net), .O(n3046));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2055_3_lut (.I0(n2946), .I1(n8262[15]), .I2(n294[3]), 
            .I3(GND_net), .O(n3054));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2048_3_lut (.I0(n2939), .I1(n8262[22]), .I2(n294[3]), 
            .I3(GND_net), .O(n3047));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2049_3_lut (.I0(n2940), .I1(n8262[21]), .I2(n294[3]), 
            .I3(GND_net), .O(n3048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2050_3_lut (.I0(n2941), .I1(n8262[20]), .I2(n294[3]), 
            .I3(GND_net), .O(n3049));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2053_3_lut (.I0(n2944), .I1(n8262[17]), .I2(n294[3]), 
            .I3(GND_net), .O(n3052));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1045 (.I0(baudrate[27]), .I1(baudrate[28]), .I2(GND_net), 
            .I3(GND_net), .O(n59250));
    defparam i1_2_lut_adj_1045.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2070_i35_2_lut (.I0(n3052), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5217));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2051_3_lut (.I0(n2942), .I1(n8262[19]), .I2(n294[3]), 
            .I3(GND_net), .O(n3050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i39_2_lut (.I0(n3050), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5218));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2054_3_lut (.I0(n2945), .I1(n8262[16]), .I2(n294[3]), 
            .I3(GND_net), .O(n3053));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49461_2_lut_4_lut (.I0(n66044), .I1(baudrate[22]), .I2(n3151), 
            .I3(n25214), .O(n294[1]));
    defparam i49461_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_2070_i33_2_lut (.I0(n3053), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5219));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2052_3_lut (.I0(n2943), .I1(n8262[18]), .I2(n294[3]), 
            .I3(GND_net), .O(n3051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1046 (.I0(n55184), .I1(r_SM_Main[0]), .I2(r_SM_Main[2]), 
            .I3(r_SM_Main[1]), .O(n58594));
    defparam i1_3_lut_4_lut_adj_1046.LUT_INIT = 16'hfdfc;
    SB_LUT4 div_37_LessThan_2070_i37_2_lut (.I0(n3051), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5220));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2056_3_lut (.I0(n2947), .I1(n8262[14]), .I2(n294[3]), 
            .I3(GND_net), .O(n3055));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2057_3_lut (.I0(n2948), .I1(n8262[13]), .I2(n294[3]), 
            .I3(GND_net), .O(n3056));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1047 (.I0(baudrate[13]), .I1(baudrate[14]), .I2(GND_net), 
            .I3(GND_net), .O(n59010));
    defparam i1_2_lut_adj_1047.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2070_i27_2_lut (.I0(n3056), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5221));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i29_2_lut (.I0(n3055), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5222));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2058_3_lut (.I0(n2949), .I1(n8262[12]), .I2(n294[3]), 
            .I3(GND_net), .O(n3057));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2059_3_lut (.I0(n2950), .I1(n8262[11]), .I2(n294[3]), 
            .I3(GND_net), .O(n3058));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i23_2_lut (.I0(n3058), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5223));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i25_2_lut (.I0(n3057), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5224));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2065_3_lut (.I0(n2956), .I1(n8262[5]), .I2(n294[3]), 
            .I3(GND_net), .O(n3064));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2066_3_lut (.I0(n2957), .I1(n8262[4]), .I2(n294[3]), 
            .I3(GND_net), .O(n3065));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i11_2_lut (.I0(n3064), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5225));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2060_3_lut (.I0(n2951), .I1(n8262[10]), .I2(n294[3]), 
            .I3(GND_net), .O(n3059));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2064_3_lut (.I0(n2955), .I1(n8262[6]), .I2(n294[3]), 
            .I3(GND_net), .O(n3063));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1048 (.I0(baudrate[6]), .I1(baudrate[7]), .I2(GND_net), 
            .I3(GND_net), .O(n59232));
    defparam i1_2_lut_adj_1048.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2070_i13_2_lut (.I0(n3063), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5226));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i21_2_lut (.I0(n3059), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5227));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2061_3_lut (.I0(n2952), .I1(n8262[9]), .I2(n294[3]), 
            .I3(GND_net), .O(n3060));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2062_3_lut (.I0(n2953), .I1(n8262[8]), .I2(n294[3]), 
            .I3(GND_net), .O(n3061));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2063_3_lut (.I0(n2954), .I1(n8262[7]), .I2(n294[3]), 
            .I3(GND_net), .O(n3062));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_2070_i15_2_lut (.I0(n3062), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i17_2_lut (.I0(n3061), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5229));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i19_2_lut (.I0(n3060), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5230));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_2070_i31_2_lut (.I0(n3054), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5231));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46733_4_lut (.I0(n31_adj_5231), .I1(n19_adj_5230), .I2(n17_adj_5229), 
            .I3(n15_adj_5228), .O(n63795));
    defparam i46733_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_2_lut_adj_1049 (.I0(baudrate[8]), .I1(baudrate[9]), .I2(GND_net), 
            .I3(GND_net), .O(n59230));
    defparam i1_2_lut_adj_1049.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_2141_i8_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n3170), .I3(GND_net), .O(n8_adj_5215));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1050 (.I0(baudrate[4]), .I1(baudrate[5]), .I2(GND_net), 
            .I3(GND_net), .O(n59170));
    defparam i1_2_lut_adj_1050.LUT_INIT = 16'heeee;
    SB_LUT4 i47724_4_lut (.I0(n13_adj_5226), .I1(n11_adj_5225), .I2(n3065), 
            .I3(baudrate[2]), .O(n64786));
    defparam i47724_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i48231_4_lut (.I0(n19_adj_5230), .I1(n17_adj_5229), .I2(n15_adj_5228), 
            .I3(n64786), .O(n65293));
    defparam i48231_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48229_4_lut (.I0(n25_adj_5224), .I1(n23_adj_5223), .I2(n21_adj_5227), 
            .I3(n65293), .O(n65291));
    defparam i48229_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_1051 (.I0(baudrate[28]), .I1(baudrate[27]), .I2(baudrate[31]), 
            .I3(baudrate[26]), .O(n59148));
    defparam i1_4_lut_adj_1051.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2141_i12_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n3167), .I3(GND_net), .O(n12_adj_5214));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46735_4_lut (.I0(n31_adj_5231), .I1(n29_adj_5222), .I2(n27_adj_5221), 
            .I3(n65291), .O(n63797));
    defparam i46735_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_2070_i8_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n3066), .I3(GND_net), .O(n8_adj_5232));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48456_3_lut (.I0(n8_adj_5232), .I1(baudrate[13]), .I2(n31_adj_5231), 
            .I3(GND_net), .O(n65518));   // verilog/uart_rx.v(119[33:55])
    defparam i48456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46673_2_lut_4_lut (.I0(n3157), .I1(baudrate[16]), .I2(n3166), 
            .I3(baudrate[7]), .O(n63735));
    defparam i46673_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_4_lut_adj_1052 (.I0(n59148), .I1(n59308), .I2(n59252), 
            .I3(n59248), .O(n25205));
    defparam i1_4_lut_adj_1052.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2141_i14_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n3157), .I3(GND_net), .O(n14_adj_5212));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i14_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48457_3_lut (.I0(n65518), .I1(baudrate[14]), .I2(n33_adj_5219), 
            .I3(GND_net), .O(n65519));   // verilog/uart_rx.v(119[33:55])
    defparam i48457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_450_i46_4_lut (.I0(n63061), .I1(baudrate[2]), 
            .I2(n66281), .I3(n48_adj_5031), .O(n46_adj_5233));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i46_4_lut.LUT_INIT = 16'hc0e8;
    SB_LUT4 div_37_LessThan_450_i48_3_lut (.I0(n46_adj_5233), .I1(baudrate[3]), 
            .I2(n56317), .I3(GND_net), .O(n48_adj_5234));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_450_i48_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i1_4_lut_adj_1053 (.I0(n59170), .I1(n59230), .I2(n59232), 
            .I3(n59228), .O(n59182));
    defparam i1_4_lut_adj_1053.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_2141_i10_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n3165), .I3(GND_net), .O(n10_adj_5216));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2141_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_2070_i34_3_lut (.I0(n16_adj_5208), .I1(baudrate[17]), 
            .I2(n39_adj_5218), .I3(GND_net), .O(n34_adj_5235));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i34_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1054 (.I0(n59182), .I1(n25205), .I2(n59174), 
            .I3(n59310), .O(n25152));
    defparam i1_4_lut_adj_1054.LUT_INIT = 16'hfffe;
    SB_LUT4 i42883_2_lut (.I0(baudrate[7]), .I1(n59934), .I2(GND_net), 
            .I3(GND_net), .O(n59936));
    defparam i42883_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i46719_4_lut (.I0(n37_adj_5220), .I1(n35_adj_5217), .I2(n33_adj_5219), 
            .I3(n63795), .O(n63781));
    defparam i46719_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48937_4_lut (.I0(n34_adj_5235), .I1(n14_adj_5204), .I2(n39_adj_5218), 
            .I3(n63779), .O(n65999));   // verilog/uart_rx.v(119[33:55])
    defparam i48937_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47439_3_lut (.I0(n65519), .I1(baudrate[15]), .I2(n35_adj_5217), 
            .I3(GND_net), .O(n64501));   // verilog/uart_rx.v(119[33:55])
    defparam i47439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48458_3_lut (.I0(n10_adj_5203), .I1(baudrate[10]), .I2(n25_adj_5224), 
            .I3(GND_net), .O(n65520));   // verilog/uart_rx.v(119[33:55])
    defparam i48458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48459_3_lut (.I0(n65520), .I1(baudrate[11]), .I2(n27_adj_5221), 
            .I3(GND_net), .O(n65521));   // verilog/uart_rx.v(119[33:55])
    defparam i48459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47706_4_lut (.I0(n27_adj_5221), .I1(n25_adj_5224), .I2(n23_adj_5223), 
            .I3(n63812), .O(n64768));
    defparam i47706_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i46697_2_lut_4_lut (.I0(n3165), .I1(baudrate[8]), .I2(n3169), 
            .I3(baudrate[4]), .O(n63759));
    defparam i46697_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_2070_i20_3_lut (.I0(n12_adj_5210), .I1(baudrate[9]), 
            .I2(n23_adj_5223), .I3(GND_net), .O(n20_adj_5236));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_2070_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47437_3_lut (.I0(n65521), .I1(baudrate[12]), .I2(n29_adj_5222), 
            .I3(GND_net), .O(n64499));   // verilog/uart_rx.v(119[33:55])
    defparam i47437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48627_4_lut (.I0(n37_adj_5220), .I1(n35_adj_5217), .I2(n33_adj_5219), 
            .I3(n63797), .O(n65689));
    defparam i48627_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i49130_4_lut (.I0(n64501), .I1(n65999), .I2(n39_adj_5218), 
            .I3(n63781), .O(n66192));   // verilog/uart_rx.v(119[33:55])
    defparam i49130_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48519_4_lut (.I0(n64499), .I1(n20_adj_5236), .I2(n29_adj_5222), 
            .I3(n64768), .O(n65581));   // verilog/uart_rx.v(119[33:55])
    defparam i48519_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_2_lut_3_lut (.I0(baudrate[26]), .I1(baudrate[30]), .I2(baudrate[23]), 
            .I3(GND_net), .O(n59398));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i49189_4_lut (.I0(n65581), .I1(n66192), .I2(n39_adj_5218), 
            .I3(n65689), .O(n66251));   // verilog/uart_rx.v(119[33:55])
    defparam i49189_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49190_3_lut (.I0(n66251), .I1(baudrate[18]), .I2(n3049), 
            .I3(GND_net), .O(n66252));   // verilog/uart_rx.v(119[33:55])
    defparam i49190_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49180_3_lut (.I0(n66252), .I1(baudrate[19]), .I2(n3048), 
            .I3(GND_net), .O(n66242));   // verilog/uart_rx.v(119[33:55])
    defparam i49180_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48696_3_lut (.I0(n66242), .I1(baudrate[20]), .I2(n3047), 
            .I3(GND_net), .O(n65758));   // verilog/uart_rx.v(119[33:55])
    defparam i48696_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_2_lut_adj_1055 (.I0(baudrate[5]), .I1(baudrate[6]), .I2(GND_net), 
            .I3(GND_net), .O(n59018));
    defparam i1_2_lut_adj_1055.LUT_INIT = 16'heeee;
    SB_LUT4 div_37_LessThan_557_i42_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n805), .I3(GND_net), .O(n42_adj_5237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_557_i42_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49437_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(n59692), .I2(n48_adj_5083), 
            .I3(baudrate[15]), .O(n294[9]));
    defparam i49437_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i42823_2_lut_3_lut_4_lut (.I0(baudrate[16]), .I1(n59692), .I2(n59010), 
            .I3(baudrate[15]), .O(n59876));
    defparam i42823_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48739_3_lut (.I0(n42_adj_5237), .I1(baudrate[2]), .I2(n804), 
            .I3(GND_net), .O(n65801));   // verilog/uart_rx.v(119[33:55])
    defparam i48739_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48740_3_lut (.I0(n65801), .I1(baudrate[3]), .I2(n803), .I3(GND_net), 
            .O(n65802));   // verilog/uart_rx.v(119[33:55])
    defparam i48740_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48463_3_lut (.I0(n65802), .I1(baudrate[4]), .I2(n56321), 
            .I3(GND_net), .O(n48_adj_5238));   // verilog/uart_rx.v(119[33:55])
    defparam i48463_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i42856_1_lut_2_lut (.I0(baudrate[12]), .I1(n59876), .I2(GND_net), 
            .I3(GND_net), .O(n56602));
    defparam i42856_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 div_37_LessThan_1062_i32_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n58472), .I3(n48_adj_5145), .O(n32_adj_5174));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1062_i32_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i1_3_lut_adj_1056 (.I0(n25152), .I1(n48_adj_5234), .I2(baudrate[0]), 
            .I3(GND_net), .O(n805));
    defparam i1_3_lut_adj_1056.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_4_lut_adj_1057 (.I0(n66238), .I1(baudrate[19]), .I2(n2827), 
            .I3(n58486), .O(n2957));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1057.LUT_INIT = 16'h7100;
    SB_LUT4 i49452_2_lut_4_lut (.I0(n66238), .I1(baudrate[19]), .I2(n2827), 
            .I3(n25205), .O(n294[4]));   // verilog/uart_rx.v(119[33:55])
    defparam i49452_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i4194_2_lut (.I0(n962), .I1(baudrate[1]), .I2(GND_net), .I3(GND_net), 
            .O(n40_adj_5239));   // verilog/uart_rx.v(119[33:55])
    defparam i4194_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i49465_2_lut_4_lut (.I0(\r_SM_Main_2__N_3446[1] ), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main[2]), .O(n27312));
    defparam i49465_2_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i1_2_lut_4_lut_adj_1058 (.I0(n66246), .I1(baudrate[20]), .I2(n2938), 
            .I3(n58488), .O(n3066));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1058.LUT_INIT = 16'h7100;
    SB_LUT4 i49455_2_lut_4_lut (.I0(n66246), .I1(baudrate[20]), .I2(n2938), 
            .I3(n59946), .O(n294[3]));   // verilog/uart_rx.v(119[33:55])
    defparam i49455_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i642_4_lut (.I0(n805), .I1(baudrate[1]), .I2(n294[19]), 
            .I3(baudrate[0]), .O(n961));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i642_4_lut.LUT_INIT = 16'h9a6a;
    SB_LUT4 div_37_i745_4_lut (.I0(n961), .I1(n40_adj_5239), .I2(n294[18]), 
            .I3(baudrate[2]), .O(n1114));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i745_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 div_37_i846_3_lut (.I0(n1114), .I1(n7898[20]), .I2(n294[17]), 
            .I3(GND_net), .O(n1264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i945_3_lut (.I0(n1264), .I1(n7924[20]), .I2(n294[16]), 
            .I3(GND_net), .O(n1411));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1042_3_lut (.I0(n1411), .I1(n7950[20]), .I2(n294[15]), 
            .I3(GND_net), .O(n1555));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1974_3_lut (.I0(n2827), .I1(n8236[23]), .I2(n294[4]), 
            .I3(GND_net), .O(n2938));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1981_3_lut (.I0(n2834), .I1(n8236[16]), .I2(n294[4]), 
            .I3(GND_net), .O(n2945));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1975_3_lut (.I0(n2828), .I1(n8236[22]), .I2(n294[4]), 
            .I3(GND_net), .O(n2939));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1976_3_lut (.I0(n2829), .I1(n8236[21]), .I2(n294[4]), 
            .I3(GND_net), .O(n2940));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1979_3_lut (.I0(n2832), .I1(n8236[18]), .I2(n294[4]), 
            .I3(GND_net), .O(n2943));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1980_3_lut (.I0(n2833), .I1(n8236[17]), .I2(n294[4]), 
            .I3(GND_net), .O(n2944));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i35_2_lut (.I0(n2944), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5240));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i37_2_lut (.I0(n2943), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5241));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1977_3_lut (.I0(n2830), .I1(n8236[20]), .I2(n294[4]), 
            .I3(GND_net), .O(n2941));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i41_2_lut (.I0(n2941), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5242));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1978_3_lut (.I0(n2831), .I1(n8236[19]), .I2(n294[4]), 
            .I3(GND_net), .O(n2942));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i39_2_lut (.I0(n2942), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5243));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1982_3_lut (.I0(n2835), .I1(n8236[15]), .I2(n294[4]), 
            .I3(GND_net), .O(n2946));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1983_3_lut (.I0(n2836), .I1(n8236[14]), .I2(n294[4]), 
            .I3(GND_net), .O(n2947));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1059 (.I0(baudrate[6]), .I1(baudrate[7]), 
            .I2(baudrate[8]), .I3(baudrate[9]), .O(n59240));
    defparam i1_2_lut_4_lut_adj_1059.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1997_i29_2_lut (.I0(n2947), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5244));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i31_2_lut (.I0(n2946), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5245));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1984_3_lut (.I0(n2837), .I1(n8236[13]), .I2(n294[4]), 
            .I3(GND_net), .O(n2948));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1985_3_lut (.I0(n2838), .I1(n8236[12]), .I2(n294[4]), 
            .I3(GND_net), .O(n2949));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1986_3_lut (.I0(n2839), .I1(n8236[11]), .I2(n294[4]), 
            .I3(GND_net), .O(n2950));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i23_2_lut (.I0(n2950), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5246));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i25_2_lut (.I0(n2949), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5247));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i27_2_lut (.I0(n2948), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5248));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1990_3_lut (.I0(n2843), .I1(n8236[7]), .I2(n294[4]), 
            .I3(GND_net), .O(n2954));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1991_3_lut (.I0(n2844), .I1(n8236[6]), .I2(n294[4]), 
            .I3(GND_net), .O(n2955));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1992_3_lut (.I0(n2845), .I1(n8236[5]), .I2(n294[4]), 
            .I3(GND_net), .O(n2956));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i13_2_lut (.I0(n2955), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_5249));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i15_2_lut (.I0(n2954), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5250));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1987_3_lut (.I0(n2840), .I1(n8236[10]), .I2(n294[4]), 
            .I3(GND_net), .O(n2951));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1988_3_lut (.I0(n2841), .I1(n8236[9]), .I2(n294[4]), 
            .I3(GND_net), .O(n2952));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1989_3_lut (.I0(n2842), .I1(n8236[8]), .I2(n294[4]), 
            .I3(GND_net), .O(n2953));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i17_2_lut (.I0(n2953), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5251));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i19_2_lut (.I0(n2952), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5252));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i21_2_lut (.I0(n2951), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5253));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1997_i33_2_lut (.I0(n2945), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5254));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46783_4_lut (.I0(n33_adj_5254), .I1(n21_adj_5253), .I2(n19_adj_5252), 
            .I3(n17_adj_5251), .O(n63845));
    defparam i46783_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47765_4_lut (.I0(n15_adj_5250), .I1(n13_adj_5249), .I2(n2956), 
            .I3(baudrate[2]), .O(n64827));
    defparam i47765_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i48253_4_lut (.I0(n21_adj_5253), .I1(n19_adj_5252), .I2(n17_adj_5251), 
            .I3(n64827), .O(n65315));
    defparam i48253_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 div_37_i1137_3_lut (.I0(n1555), .I1(n7976[20]), .I2(n294[14]), 
            .I3(GND_net), .O(n1696));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1060 (.I0(baudrate[10]), .I1(baudrate[11]), 
            .I2(baudrate[12]), .I3(baudrate[13]), .O(n59238));
    defparam i1_2_lut_4_lut_adj_1060.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1230_3_lut (.I0(n1696), .I1(n8002[20]), .I2(n294[13]), 
            .I3(GND_net), .O(n1834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48251_4_lut (.I0(n27_adj_5248), .I1(n25_adj_5247), .I2(n23_adj_5246), 
            .I3(n65315), .O(n65313));
    defparam i48251_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i46785_4_lut (.I0(n33_adj_5254), .I1(n31_adj_5245), .I2(n29_adj_5244), 
            .I3(n65313), .O(n63847));
    defparam i46785_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1997_i10_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2957), .I3(GND_net), .O(n10_adj_5255));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48486_3_lut (.I0(n10_adj_5255), .I1(baudrate[13]), .I2(n33_adj_5254), 
            .I3(GND_net), .O(n65548));   // verilog/uart_rx.v(119[33:55])
    defparam i48486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48487_3_lut (.I0(n65548), .I1(baudrate[14]), .I2(n35_adj_5240), 
            .I3(GND_net), .O(n65549));   // verilog/uart_rx.v(119[33:55])
    defparam i48487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1321_3_lut (.I0(n1834), .I1(n8028[20]), .I2(n294[12]), 
            .I3(GND_net), .O(n1969));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i36_3_lut (.I0(n18_adj_5191), .I1(baudrate[17]), 
            .I2(n41_adj_5242), .I3(GND_net), .O(n36_adj_5256));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i36_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46775_4_lut (.I0(n39_adj_5243), .I1(n37_adj_5241), .I2(n35_adj_5240), 
            .I3(n63845), .O(n63837));
    defparam i46775_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48935_4_lut (.I0(n36_adj_5256), .I1(n16_adj_5190), .I2(n41_adj_5242), 
            .I3(n63834), .O(n65997));   // verilog/uart_rx.v(119[33:55])
    defparam i48935_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47427_3_lut (.I0(n65549), .I1(baudrate[15]), .I2(n37_adj_5241), 
            .I3(GND_net), .O(n64489));   // verilog/uart_rx.v(119[33:55])
    defparam i47427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1997_i22_3_lut (.I0(n14_adj_5188), .I1(baudrate[9]), 
            .I2(n25_adj_5247), .I3(GND_net), .O(n22_adj_5257));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1997_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48929_4_lut (.I0(n22_adj_5257), .I1(n12_adj_5187), .I2(n25_adj_5247), 
            .I3(n63866), .O(n65991));   // verilog/uart_rx.v(119[33:55])
    defparam i48929_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48930_3_lut (.I0(n65991), .I1(baudrate[10]), .I2(n27_adj_5248), 
            .I3(GND_net), .O(n65992));   // verilog/uart_rx.v(119[33:55])
    defparam i48930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48778_3_lut (.I0(n65992), .I1(baudrate[11]), .I2(n29_adj_5244), 
            .I3(GND_net), .O(n65840));   // verilog/uart_rx.v(119[33:55])
    defparam i48778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48635_4_lut (.I0(n39_adj_5243), .I1(n37_adj_5241), .I2(n35_adj_5240), 
            .I3(n63847), .O(n65697));
    defparam i48635_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i49128_4_lut (.I0(n64489), .I1(n65997), .I2(n41_adj_5242), 
            .I3(n63837), .O(n66190));   // verilog/uart_rx.v(119[33:55])
    defparam i49128_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47425_3_lut (.I0(n65840), .I1(baudrate[12]), .I2(n31_adj_5245), 
            .I3(GND_net), .O(n64487));   // verilog/uart_rx.v(119[33:55])
    defparam i47425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49185_4_lut (.I0(n64487), .I1(n66190), .I2(n41_adj_5242), 
            .I3(n65697), .O(n66247));   // verilog/uart_rx.v(119[33:55])
    defparam i49185_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49186_3_lut (.I0(n66247), .I1(baudrate[18]), .I2(n2940), 
            .I3(GND_net), .O(n66248));   // verilog/uart_rx.v(119[33:55])
    defparam i49186_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49184_3_lut (.I0(n66248), .I1(baudrate[19]), .I2(n2939), 
            .I3(GND_net), .O(n66246));   // verilog/uart_rx.v(119[33:55])
    defparam i49184_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1899_3_lut (.I0(n2713), .I1(n8210[23]), .I2(n294[5]), 
            .I3(GND_net), .O(n2827));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i41_2_lut (.I0(n1969), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5258));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1905_3_lut (.I0(n2719), .I1(n8210[17]), .I2(n294[5]), 
            .I3(GND_net), .O(n2833));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1900_3_lut (.I0(n2714), .I1(n8210[22]), .I2(n294[5]), 
            .I3(GND_net), .O(n2828));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1903_3_lut (.I0(n2717), .I1(n8210[19]), .I2(n294[5]), 
            .I3(GND_net), .O(n2831));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i39_2_lut (.I0(n2831), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_5259));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1904_3_lut (.I0(n2718), .I1(n8210[18]), .I2(n294[5]), 
            .I3(GND_net), .O(n2832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i37_2_lut (.I0(n2832), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_5260));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1901_3_lut (.I0(n2715), .I1(n8210[21]), .I2(n294[5]), 
            .I3(GND_net), .O(n2829));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1061 (.I0(n59018), .I1(n59936), .I2(baudrate[0]), 
            .I3(n48_adj_5238), .O(n962));
    defparam i1_3_lut_4_lut_adj_1061.LUT_INIT = 16'h0010;
    SB_LUT4 div_37_LessThan_1922_i43_2_lut (.I0(n2829), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_5261));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1902_3_lut (.I0(n2716), .I1(n8210[20]), .I2(n294[5]), 
            .I3(GND_net), .O(n2830));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i41_2_lut (.I0(n2830), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1341_i27_2_lut (.I0(n1976), .I1(baudrate[2]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5263));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46193_4_lut (.I0(n33_adj_5126), .I1(n31_adj_5124), .I2(n29_adj_5125), 
            .I3(n27_adj_5263), .O(n63255));
    defparam i46193_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i49261_2_lut_3_lut (.I0(n59018), .I1(n59936), .I2(n48_adj_5238), 
            .I3(GND_net), .O(n294[19]));
    defparam i49261_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 div_37_i1906_3_lut (.I0(n2720), .I1(n8210[16]), .I2(n294[5]), 
            .I3(GND_net), .O(n2834));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1907_3_lut (.I0(n2721), .I1(n8210[15]), .I2(n294[5]), 
            .I3(GND_net), .O(n2835));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i31_2_lut (.I0(n2835), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_5264));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1062 (.I0(n65758), .I1(baudrate[21]), .I2(n3046), 
            .I3(n58490), .O(n3172));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1062.LUT_INIT = 16'h7100;
    SB_LUT4 i49458_2_lut_4_lut (.I0(n65758), .I1(baudrate[21]), .I2(n3046), 
            .I3(n25211), .O(n294[2]));   // verilog/uart_rx.v(119[33:55])
    defparam i49458_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1922_i33_2_lut (.I0(n2834), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_5265));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1908_3_lut (.I0(n2722), .I1(n8210[14]), .I2(n294[5]), 
            .I3(GND_net), .O(n2836));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1909_3_lut (.I0(n2723), .I1(n8210[13]), .I2(n294[5]), 
            .I3(GND_net), .O(n2837));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1909_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1910_3_lut (.I0(n2724), .I1(n8210[12]), .I2(n294[5]), 
            .I3(GND_net), .O(n2838));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1910_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i25_2_lut (.I0(n2838), .I1(baudrate[8]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5266));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i27_2_lut (.I0(n2837), .I1(baudrate[9]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5267));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i29_2_lut (.I0(n2836), .I1(baudrate[10]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_5268));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1914_3_lut (.I0(n2728), .I1(n8210[8]), .I2(n294[5]), 
            .I3(GND_net), .O(n2842));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1915_3_lut (.I0(n2729), .I1(n8210[7]), .I2(n294[5]), 
            .I3(GND_net), .O(n2843));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1916_3_lut (.I0(n2730), .I1(n8210[6]), .I2(n294[5]), 
            .I3(GND_net), .O(n2844));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i15_2_lut (.I0(n2843), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5269));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i17_2_lut (.I0(n2842), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_5270));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i1911_3_lut (.I0(n2725), .I1(n8210[11]), .I2(n294[5]), 
            .I3(GND_net), .O(n2839));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1912_3_lut (.I0(n2726), .I1(n8210[10]), .I2(n294[5]), 
            .I3(GND_net), .O(n2840));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1913_3_lut (.I0(n2727), .I1(n8210[9]), .I2(n294[5]), 
            .I3(GND_net), .O(n2841));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1913_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i19_2_lut (.I0(n2841), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_5271));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i21_2_lut (.I0(n2840), .I1(baudrate[6]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_5272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i23_2_lut (.I0(n2839), .I1(baudrate[7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5273));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1922_i35_2_lut (.I0(n2833), .I1(baudrate[13]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_5274));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46846_4_lut (.I0(n35_adj_5274), .I1(n23_adj_5273), .I2(n21_adj_5272), 
            .I3(n19_adj_5271), .O(n63908));
    defparam i46846_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i47819_4_lut (.I0(n17_adj_5270), .I1(n15_adj_5269), .I2(n2844), 
            .I3(baudrate[2]), .O(n64881));
    defparam i47819_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i4200_2_lut_3_lut (.I0(baudrate[2]), .I1(n962), .I2(baudrate[1]), 
            .I3(GND_net), .O(n9784));   // verilog/uart_rx.v(119[33:55])
    defparam i4200_2_lut_3_lut.LUT_INIT = 16'h4545;
    SB_LUT4 i48283_4_lut (.I0(n23_adj_5273), .I1(n21_adj_5272), .I2(n19_adj_5271), 
            .I3(n64881), .O(n65345));
    defparam i48283_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48281_4_lut (.I0(n29_adj_5268), .I1(n27_adj_5267), .I2(n25_adj_5266), 
            .I3(n65345), .O(n65343));
    defparam i48281_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i46848_4_lut (.I0(n35_adj_5274), .I1(n33_adj_5265), .I2(n31_adj_5264), 
            .I3(n65343), .O(n63910));
    defparam i46848_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i5807_2_lut_3_lut (.I0(n805), .I1(baudrate[1]), .I2(baudrate[0]), 
            .I3(GND_net), .O(n21309));   // verilog/uart_rx.v(119[33:55])
    defparam i5807_2_lut_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i42835_2_lut_3_lut (.I0(baudrate[19]), .I1(baudrate[20]), .I2(baudrate[4]), 
            .I3(GND_net), .O(n59888));
    defparam i42835_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_37_LessThan_1922_i12_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n2845), .I3(GND_net), .O(n12_adj_5275));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48527_3_lut (.I0(n12_adj_5275), .I1(baudrate[13]), .I2(n35_adj_5274), 
            .I3(GND_net), .O(n65589));   // verilog/uart_rx.v(119[33:55])
    defparam i48527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i38_3_lut (.I0(n30_adj_5185), .I1(baudrate[9]), 
            .I2(n41_adj_5258), .I3(GND_net), .O(n38_adj_5276));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1341_i26_3_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n1977), .I3(GND_net), .O(n26_adj_5277));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1341_i26_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48719_3_lut (.I0(n26_adj_5277), .I1(baudrate[5]), .I2(n33_adj_5126), 
            .I3(GND_net), .O(n65781));   // verilog/uart_rx.v(119[33:55])
    defparam i48719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i39547_1_lut_4_lut (.I0(n59396), .I1(n59398), .I2(n59250), 
            .I3(n59394), .O(n56561));
    defparam i39547_1_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i48720_3_lut (.I0(n65781), .I1(baudrate[6]), .I2(n35_adj_5127), 
            .I3(GND_net), .O(n65782));   // verilog/uart_rx.v(119[33:55])
    defparam i48720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i38_3_lut (.I0(n20_adj_5179), .I1(baudrate[17]), 
            .I2(n43_adj_5261), .I3(GND_net), .O(n38_adj_5278));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48528_3_lut (.I0(n65589), .I1(baudrate[14]), .I2(n37_adj_5260), 
            .I3(GND_net), .O(n65590));   // verilog/uart_rx.v(119[33:55])
    defparam i48528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46836_4_lut (.I0(n41_adj_5262), .I1(n39_adj_5259), .I2(n37_adj_5260), 
            .I3(n63908), .O(n63898));
    defparam i46836_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46187_4_lut (.I0(n39_adj_5128), .I1(n37_adj_5129), .I2(n35_adj_5127), 
            .I3(n63255), .O(n63249));
    defparam i46187_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48923_4_lut (.I0(n38_adj_5278), .I1(n18_adj_5178), .I2(n43_adj_5261), 
            .I3(n63888), .O(n65985));   // verilog/uart_rx.v(119[33:55])
    defparam i48923_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49043_4_lut (.I0(n38_adj_5276), .I1(n28_adj_5183), .I2(n41_adj_5258), 
            .I3(n63246), .O(n66105));   // verilog/uart_rx.v(119[33:55])
    defparam i49043_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48493_3_lut (.I0(n65782), .I1(baudrate[7]), .I2(n37_adj_5129), 
            .I3(GND_net), .O(n65555));   // verilog/uart_rx.v(119[33:55])
    defparam i48493_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49171_4_lut (.I0(n65555), .I1(n66105), .I2(n41_adj_5258), 
            .I3(n63249), .O(n66233));   // verilog/uart_rx.v(119[33:55])
    defparam i49171_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49172_3_lut (.I0(n66233), .I1(baudrate[10]), .I2(n1968), 
            .I3(GND_net), .O(n66234));   // verilog/uart_rx.v(119[33:55])
    defparam i49172_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i42884_1_lut_2_lut (.I0(baudrate[7]), .I1(n59934), .I2(GND_net), 
            .I3(GND_net), .O(n56619));
    defparam i42884_1_lut_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i47419_3_lut (.I0(n65590), .I1(baudrate[15]), .I2(n39_adj_5259), 
            .I3(GND_net), .O(n64481));   // verilog/uart_rx.v(119[33:55])
    defparam i47419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49127_3_lut (.I0(n66234), .I1(baudrate[11]), .I2(n1967), 
            .I3(GND_net), .O(n66189));   // verilog/uart_rx.v(119[33:55])
    defparam i49127_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49068_3_lut (.I0(n66189), .I1(baudrate[12]), .I2(n1966), 
            .I3(GND_net), .O(n48_adj_5279));   // verilog/uart_rx.v(119[33:55])
    defparam i49068_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i1_3_lut_adj_1063 (.I0(n59876), .I1(n48_adj_5279), .I2(n8054[11]), 
            .I3(GND_net), .O(n2110));
    defparam i1_3_lut_adj_1063.LUT_INIT = 16'h1010;
    SB_LUT4 div_37_i1506_3_lut (.I0(n2110), .I1(n8080[11]), .I2(n294[10]), 
            .I3(GND_net), .O(n2239));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1922_i24_3_lut (.I0(n16_adj_5176), .I1(baudrate[9]), 
            .I2(n27_adj_5267), .I3(GND_net), .O(n24_adj_5280));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1922_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48921_4_lut (.I0(n24_adj_5280), .I1(n14_adj_5175), .I2(n27_adj_5267), 
            .I3(n63927), .O(n65983));   // verilog/uart_rx.v(119[33:55])
    defparam i48921_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i1591_3_lut (.I0(n2239), .I1(n8106[11]), .I2(n294[9]), 
            .I3(GND_net), .O(n2365));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48922_3_lut (.I0(n65983), .I1(baudrate[10]), .I2(n29_adj_5268), 
            .I3(GND_net), .O(n65984));   // verilog/uart_rx.v(119[33:55])
    defparam i48922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48788_3_lut (.I0(n65984), .I1(baudrate[11]), .I2(n31_adj_5264), 
            .I3(GND_net), .O(n65850));   // verilog/uart_rx.v(119[33:55])
    defparam i48788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48647_4_lut (.I0(n41_adj_5262), .I1(n39_adj_5259), .I2(n37_adj_5260), 
            .I3(n63910), .O(n65709));
    defparam i48647_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i49122_4_lut (.I0(n64481), .I1(n65985), .I2(n43_adj_5261), 
            .I3(n63898), .O(n66184));   // verilog/uart_rx.v(119[33:55])
    defparam i49122_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1064 (.I0(n59302), .I1(n59298), .I2(n59300), 
            .I3(n59296), .O(n59282));
    defparam i1_4_lut_adj_1064.LUT_INIT = 16'hfffe;
    SB_LUT4 i47417_3_lut (.I0(n65850), .I1(baudrate[12]), .I2(n33_adj_5265), 
            .I3(GND_net), .O(n64479));   // verilog/uart_rx.v(119[33:55])
    defparam i47417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1065 (.I0(baudrate[30]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n59248));
    defparam i1_2_lut_adj_1065.LUT_INIT = 16'heeee;
    SB_LUT4 i49175_4_lut (.I0(n64479), .I1(n66184), .I2(n43_adj_5261), 
            .I3(n65709), .O(n66237));   // verilog/uart_rx.v(119[33:55])
    defparam i49175_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49176_3_lut (.I0(n66237), .I1(baudrate[18]), .I2(n2828), 
            .I3(GND_net), .O(n66238));   // verilog/uart_rx.v(119[33:55])
    defparam i49176_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1822_3_lut (.I0(n2596), .I1(n8184[23]), .I2(n294[6]), 
            .I3(GND_net), .O(n2713));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1827_3_lut (.I0(n2601), .I1(n8184[18]), .I2(n294[6]), 
            .I3(GND_net), .O(n2718));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1825_3_lut (.I0(n2599), .I1(n8184[20]), .I2(n294[6]), 
            .I3(GND_net), .O(n2716));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i41_2_lut (.I0(n2716), .I1(baudrate[15]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_5014));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i22699_rep_9_2_lut (.I0(n7976[14]), .I1(n294[14]), .I2(GND_net), 
            .I3(GND_net), .O(n56605));   // verilog/uart_rx.v(119[33:55])
    defparam i22699_rep_9_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_37_LessThan_1157_i32_4_lut (.I0(n56605), .I1(baudrate[2]), 
            .I2(n1701), .I3(baudrate[1]), .O(n32_adj_5281));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1157_i32_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i1_2_lut_3_lut_adj_1066 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n58896), .I3(GND_net), .O(n58898));
    defparam i1_2_lut_3_lut_adj_1066.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_37_i2169_1_lut (.I0(baudrate[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1459));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2169_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_adj_1067 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n58932), .I3(GND_net), .O(n58844));
    defparam i1_2_lut_3_lut_adj_1067.LUT_INIT = 16'hf7f7;
    SB_LUT4 i48727_3_lut (.I0(n32_adj_5281), .I1(baudrate[6]), .I2(n39_adj_5130), 
            .I3(GND_net), .O(n65789));   // verilog/uart_rx.v(119[33:55])
    defparam i48727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1068 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n58896), .I3(GND_net), .O(n58970));   // verilog/uart_rx.v(98[17:39])
    defparam i1_2_lut_3_lut_adj_1068.LUT_INIT = 16'hfbfb;
    SB_LUT4 div_37_i1823_3_lut (.I0(n2597), .I1(n8184[22]), .I2(n294[6]), 
            .I3(GND_net), .O(n2714));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i45_2_lut (.I0(n2714), .I1(baudrate[17]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1069 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n58932), .I3(GND_net), .O(n58934));   // verilog/uart_rx.v(98[17:39])
    defparam i1_2_lut_3_lut_adj_1069.LUT_INIT = 16'hfbfb;
    SB_LUT4 i48728_3_lut (.I0(n65789), .I1(baudrate[7]), .I2(n41_adj_5131), 
            .I3(GND_net), .O(n65790));   // verilog/uart_rx.v(119[33:55])
    defparam i48728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47210_4_lut (.I0(n41_adj_5131), .I1(n39_adj_5130), .I2(n37_adj_5132), 
            .I3(n63316), .O(n64272));
    defparam i47210_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i1_2_lut_3_lut_adj_1070 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n58896), .I3(GND_net), .O(n58880));   // verilog/uart_rx.v(98[17:39])
    defparam i1_2_lut_3_lut_adj_1070.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut_adj_1071 (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(n58932), .I3(GND_net), .O(n58952));   // verilog/uart_rx.v(98[17:39])
    defparam i1_2_lut_3_lut_adj_1071.LUT_INIT = 16'hfdfd;
    SB_LUT4 i48083_3_lut (.I0(n34_adj_5100), .I1(baudrate[5]), .I2(n37_adj_5132), 
            .I3(GND_net), .O(n65145));   // verilog/uart_rx.v(119[33:55])
    defparam i48083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1826_3_lut (.I0(n2600), .I1(n8184[19]), .I2(n294[6]), 
            .I3(GND_net), .O(n2717));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48483_3_lut (.I0(n65790), .I1(baudrate[8]), .I2(n43_adj_5133), 
            .I3(GND_net), .O(n65545));   // verilog/uart_rx.v(119[33:55])
    defparam i48483_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1072 (.I0(n59228), .I1(n59908), .I2(n7976[14]), 
            .I3(n48_adj_5182), .O(n1702));
    defparam i1_3_lut_4_lut_adj_1072.LUT_INIT = 16'h0010;
    SB_LUT4 i1_3_lut_4_lut_adj_1073 (.I0(baudrate[28]), .I1(baudrate[25]), 
            .I2(baudrate[26]), .I3(baudrate[29]), .O(n58424));
    defparam i1_3_lut_4_lut_adj_1073.LUT_INIT = 16'hfffe;
    SB_LUT4 i42880_1_lut_2_lut_3_lut (.I0(n59228), .I1(n59908), .I2(baudrate[9]), 
            .I3(GND_net), .O(n56611));
    defparam i42880_1_lut_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i49355_2_lut_3_lut (.I0(n59228), .I1(n59908), .I2(n48_adj_5182), 
            .I3(GND_net), .O(n294[14]));
    defparam i49355_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 div_37_LessThan_1845_i39_2_lut (.I0(n2717), .I1(baudrate[14]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i42881_2_lut_3_lut_4_lut (.I0(n59228), .I1(n59908), .I2(baudrate[8]), 
            .I3(baudrate[9]), .O(n59934));
    defparam i42881_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i49352_2_lut_3_lut_4_lut (.I0(n59228), .I1(n59908), .I2(n48_adj_5145), 
            .I3(baudrate[9]), .O(n294[15]));
    defparam i49352_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i48725_4_lut (.I0(n65545), .I1(n65145), .I2(n43_adj_5133), 
            .I3(n64272), .O(n65787));   // verilog/uart_rx.v(119[33:55])
    defparam i48725_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i1824_3_lut (.I0(n2598), .I1(n8184[21]), .I2(n294[6]), 
            .I3(GND_net), .O(n2715));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48726_3_lut (.I0(n65787), .I1(baudrate[9]), .I2(n1694), .I3(GND_net), 
            .O(n65788));   // verilog/uart_rx.v(119[33:55])
    defparam i48726_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i43_2_lut (.I0(n2715), .I1(baudrate[16]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i2168_1_lut (.I0(baudrate[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1602));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2168_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1250_i30_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n1839), .I3(GND_net), .O(n30_adj_5115));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i30_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46204_2_lut_4_lut (.I0(n1834), .I1(baudrate[8]), .I2(n1838), 
            .I3(baudrate[4]), .O(n63266));
    defparam i46204_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1250_i32_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n1834), .I3(GND_net), .O(n32_adj_5112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1250_i32_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i1828_3_lut (.I0(n2602), .I1(n8184[17]), .I2(n294[6]), 
            .I3(GND_net), .O(n2719));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1829_3_lut (.I0(n2603), .I1(n8184[16]), .I2(n294[6]), 
            .I3(GND_net), .O(n2720));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48485_3_lut (.I0(n65788), .I1(baudrate[10]), .I2(n1693), 
            .I3(GND_net), .O(n48_adj_5282));   // verilog/uart_rx.v(119[33:55])
    defparam i48485_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i33_2_lut (.I0(n2720), .I1(baudrate[11]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1845_i35_2_lut (.I0(n2719), .I1(baudrate[12]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1074 (.I0(n59294), .I1(n59250), .I2(n59252), 
            .I3(baudrate[11]), .O(n59280));
    defparam i1_4_lut_adj_1074.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_i1830_3_lut (.I0(n2604), .I1(n8184[15]), .I2(n294[6]), 
            .I3(GND_net), .O(n2721));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1831_3_lut (.I0(n2605), .I1(n8184[14]), .I2(n294[6]), 
            .I3(GND_net), .O(n2722));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1832_3_lut (.I0(n2606), .I1(n8184[13]), .I2(n294[6]), 
            .I3(GND_net), .O(n2723));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1602_i22_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2365), .I3(GND_net), .O(n22_adj_5095));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47109_2_lut_4_lut (.I0(n2360), .I1(baudrate[8]), .I2(n2364), 
            .I3(baudrate[4]), .O(n64171));
    defparam i47109_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i24_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2360), .I3(GND_net), .O(n24_adj_5093));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1602_i20_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n58476), .I3(n48_adj_5083), .O(n20_adj_5098));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i20_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i1_4_lut_adj_1075 (.I0(n59280), .I1(n59282), .I2(n59270), 
            .I3(n59226), .O(n25178));
    defparam i1_4_lut_adj_1075.LUT_INIT = 16'hfffe;
    SB_LUT4 i46120_2_lut_4_lut (.I0(n2362), .I1(baudrate[6]), .I2(n2363), 
            .I3(baudrate[5]), .O(n63182));
    defparam i46120_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1602_i26_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2362), .I3(GND_net), .O(n26_adj_5091));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2167_1_lut (.I0(baudrate[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1742));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2167_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1076 (.I0(n25178), .I1(n48_adj_5282), .I2(baudrate[0]), 
            .I3(GND_net), .O(n1841));
    defparam i1_3_lut_adj_1076.LUT_INIT = 16'hefef;
    SB_LUT4 div_37_i1328_3_lut (.I0(n1841), .I1(n8028[13]), .I2(n294[12]), 
            .I3(GND_net), .O(n1976));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1417_3_lut (.I0(n1976), .I1(n8054[13]), .I2(n294[11]), 
            .I3(GND_net), .O(n2108));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1504_3_lut (.I0(n2108), .I1(n8080[13]), .I2(n294[10]), 
            .I3(GND_net), .O(n2237));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2166_1_lut (.I0(baudrate[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1879));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2166_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1589_3_lut (.I0(n2237), .I1(n8106[13]), .I2(n294[9]), 
            .I3(GND_net), .O(n2363));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1517_i24_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2238), .I3(GND_net), .O(n24_adj_5079));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46145_2_lut_4_lut (.I0(n2233), .I1(baudrate[8]), .I2(n2237), 
            .I3(baudrate[4]), .O(n63207));
    defparam i46145_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_i2165_1_lut (.I0(baudrate[10]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2013));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2165_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2164_1_lut (.I0(baudrate[11]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2144));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2164_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1517_i26_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2233), .I3(GND_net), .O(n26_adj_5077));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i26_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2163_1_lut (.I0(baudrate[12]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2272));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2163_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_LessThan_1602_i23_2_lut (.I0(n2365), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_5087));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_LessThan_1602_i25_2_lut (.I0(n2364), .I1(baudrate[4]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_5086));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46151_2_lut_4_lut (.I0(n2235), .I1(baudrate[6]), .I2(n2236), 
            .I3(baudrate[5]), .O(n63213));
    defparam i46151_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1517_i28_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2235), .I3(GND_net), .O(n28_adj_5075));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1517_i28_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_i2162_1_lut (.I0(baudrate[13]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2397));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2162_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i49340_2_lut_4_lut (.I0(n66187), .I1(baudrate[13]), .I2(n2098), 
            .I3(n25187), .O(n294[10]));   // verilog/uart_rx.v(119[33:55])
    defparam i49340_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i49413_2_lut_4_lut (.I0(n66189), .I1(baudrate[12]), .I2(n1966), 
            .I3(n59876), .O(n294[11]));
    defparam i49413_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i49337_2_lut_4_lut (.I0(n65788), .I1(baudrate[10]), .I2(n1693), 
            .I3(n25178), .O(n294[13]));   // verilog/uart_rx.v(119[33:55])
    defparam i49337_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 i42833_2_lut_4_lut (.I0(baudrate[5]), .I1(baudrate[6]), .I2(baudrate[7]), 
            .I3(baudrate[8]), .O(n59886));
    defparam i42833_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i49331_2_lut_4_lut (.I0(n65800), .I1(baudrate[5]), .I2(n56323), 
            .I3(n25163), .O(n294[18]));   // verilog/uart_rx.v(119[33:55])
    defparam i49331_2_lut_4_lut.LUT_INIT = 16'h0017;
    SB_LUT4 div_37_LessThan_1602_i27_2_lut (.I0(n2363), .I1(baudrate[5]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5085));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1602_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_37_i743_4_lut (.I0(n959), .I1(baudrate[4]), .I2(n294[18]), 
            .I3(n44_adj_5151), .O(n1112));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i743_4_lut.LUT_INIT = 16'h6a9a;
    SB_LUT4 i1_2_lut_4_lut_adj_1077 (.I0(n65572), .I1(baudrate[16]), .I2(n2476), 
            .I3(n58480), .O(n2612));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1077.LUT_INIT = 16'h7100;
    SB_LUT4 div_37_i844_3_lut (.I0(n1112), .I1(n7898[22]), .I2(n294[17]), 
            .I3(GND_net), .O(n1262));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i943_3_lut (.I0(n1262), .I1(n7924[22]), .I2(n294[16]), 
            .I3(GND_net), .O(n1409));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1040_3_lut (.I0(n1409), .I1(n7950[22]), .I2(n294[15]), 
            .I3(GND_net), .O(n1553));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1135_3_lut (.I0(n1553), .I1(n7976[22]), .I2(n294[14]), 
            .I3(GND_net), .O(n1694));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i2161_1_lut (.I0(baudrate[14]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2519));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2161_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2160_1_lut (.I0(baudrate[15]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2638));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2160_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2175_1_lut (.I0(baudrate[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n538));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2175_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i2174_1_lut (.I0(baudrate[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n858));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2174_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1228_3_lut (.I0(n1694), .I1(n8002[22]), .I2(n294[13]), 
            .I3(GND_net), .O(n1832));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1078 (.I0(n58478), .I1(n48_adj_5108), .I2(GND_net), 
            .I3(GND_net), .O(n2491));
    defparam i1_2_lut_adj_1078.LUT_INIT = 16'h2222;
    SB_LUT4 div_37_i2173_1_lut (.I0(baudrate[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n698));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2173_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_37_i1676_3_lut (.I0(n2367), .I1(n8132[9]), .I2(n294[8]), 
            .I3(GND_net), .O(n2490));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1319_3_lut (.I0(n1832), .I1(n8028[22]), .I2(n294[12]), 
            .I3(GND_net), .O(n1967));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49443_2_lut_4_lut (.I0(n65572), .I1(baudrate[16]), .I2(n2476), 
            .I3(n59692), .O(n294[7]));   // verilog/uart_rx.v(119[33:55])
    defparam i49443_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_i1408_3_lut (.I0(n1967), .I1(n8054[22]), .I2(n294[11]), 
            .I3(GND_net), .O(n2099));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_i1495_3_lut (.I0(n2099), .I1(n8080[22]), .I2(n294[10]), 
            .I3(GND_net), .O(n2228));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i1495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1079 (.I0(baudrate[28]), .I1(baudrate[25]), .I2(GND_net), 
            .I3(GND_net), .O(n58984));
    defparam i1_2_lut_adj_1079.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1080 (.I0(baudrate[22]), .I1(baudrate[23]), .I2(GND_net), 
            .I3(GND_net), .O(n59294));
    defparam i1_2_lut_adj_1080.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1081 (.I0(baudrate[18]), .I1(baudrate[19]), .I2(GND_net), 
            .I3(GND_net), .O(n59298));
    defparam i1_2_lut_adj_1081.LUT_INIT = 16'heeee;
    SB_LUT4 i4207_2_lut_3_lut (.I0(baudrate[3]), .I1(n21323), .I2(n9784), 
            .I3(GND_net), .O(n9791));   // verilog/uart_rx.v(119[33:55])
    defparam i4207_2_lut_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_2_lut_adj_1082 (.I0(baudrate[16]), .I1(baudrate[17]), .I2(GND_net), 
            .I3(GND_net), .O(n59300));
    defparam i1_2_lut_adj_1082.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_adj_1083 (.I0(n66139), .I1(baudrate[17]), .I2(n2596), 
            .I3(n58482), .O(n2730));   // verilog/uart_rx.v(119[33:55])
    defparam i1_2_lut_4_lut_adj_1083.LUT_INIT = 16'h7100;
    SB_LUT4 i49446_2_lut_4_lut (.I0(n66139), .I1(baudrate[17]), .I2(n2596), 
            .I3(n25199), .O(n294[6]));   // verilog/uart_rx.v(119[33:55])
    defparam i49446_2_lut_4_lut.LUT_INIT = 16'h0071;
    SB_LUT4 div_37_LessThan_1685_i20_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2489), .I3(GND_net), .O(n20_adj_5051));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47063_2_lut_4_lut (.I0(n2484), .I1(baudrate[8]), .I2(n2488), 
            .I3(baudrate[4]), .O(n64125));
    defparam i47063_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1685_i22_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2484), .I3(GND_net), .O(n22_adj_5050));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1685_i24_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2486), .I3(GND_net), .O(n24));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i24_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1685_i18_3_lut_4_lut (.I0(baudrate[0]), .I1(baudrate[1]), 
            .I2(n58478), .I3(n48_adj_5108), .O(n18_adj_5048));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1685_i18_3_lut_4_lut.LUT_INIT = 16'hee8e;
    SB_LUT4 i47073_2_lut_4_lut (.I0(n2486), .I1(baudrate[6]), .I2(n2487), 
            .I3(baudrate[5]), .O(n64135));
    defparam i47073_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_3_lut_4_lut_adj_1084 (.I0(n25229), .I1(n48_adj_5031), .I2(baudrate[1]), 
            .I3(baudrate[0]), .O(n44_adj_5052));
    defparam i1_3_lut_4_lut_adj_1084.LUT_INIT = 16'hefff;
    SB_LUT4 div_37_LessThan_1766_i18_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2610), .I3(GND_net), .O(n18_adj_5033));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47006_2_lut_4_lut (.I0(n2605), .I1(baudrate[8]), .I2(n2609), 
            .I3(baudrate[4]), .O(n64068));
    defparam i47006_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1430_i27_2_lut (.I0(n2108), .I1(baudrate[3]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_5283));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49322_2_lut_4_lut (.I0(n46_adj_5233), .I1(baudrate[3]), .I2(n56317), 
            .I3(n25152), .O(n294[20]));   // verilog/uart_rx.v(119[33:55])
    defparam i49322_2_lut_4_lut.LUT_INIT = 16'h0017;
    SB_LUT4 i46173_4_lut (.I0(n33_adj_5136), .I1(n31_adj_5134), .I2(n29_adj_5135), 
            .I3(n27_adj_5283), .O(n63235));
    defparam i46173_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_37_LessThan_1766_i20_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2605), .I3(GND_net), .O(n20_adj_5032));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1766_i22_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2607), .I3(GND_net), .O(n22_adj_5030));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1766_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i47025_2_lut_4_lut (.I0(n2607), .I1(baudrate[6]), .I2(n2608), 
            .I3(baudrate[5]), .O(n64087));
    defparam i47025_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i46322_2_lut_3_lut (.I0(baudrate[1]), .I1(n48_adj_5031), .I2(n25229), 
            .I3(GND_net), .O(n63384));   // verilog/uart_rx.v(119[33:55])
    defparam i46322_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 div_37_LessThan_1430_i38_3_lut (.I0(n30_adj_5147), .I1(baudrate[10]), 
            .I2(n41), .I3(GND_net), .O(n38_adj_5284));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i38_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22703_rep_8_2_lut (.I0(n8054[11]), .I1(n294[11]), .I2(GND_net), 
            .I3(GND_net), .O(n56596));   // verilog/uart_rx.v(119[33:55])
    defparam i22703_rep_8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1085 (.I0(baudrate[12]), .I1(baudrate[13]), 
            .I2(baudrate[14]), .I3(baudrate[15]), .O(n59174));
    defparam i1_2_lut_4_lut_adj_1085.LUT_INIT = 16'hfffe;
    SB_LUT4 div_37_LessThan_1430_i26_4_lut (.I0(n56596), .I1(baudrate[2]), 
            .I2(n2109), .I3(baudrate[1]), .O(n26_adj_5285));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1430_i26_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i48709_3_lut (.I0(n26_adj_5285), .I1(baudrate[6]), .I2(n33_adj_5136), 
            .I3(GND_net), .O(n65771));   // verilog/uart_rx.v(119[33:55])
    defparam i48709_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48710_3_lut (.I0(n65771), .I1(baudrate[7]), .I2(n35_adj_5137), 
            .I3(GND_net), .O(n65772));   // verilog/uart_rx.v(119[33:55])
    defparam i48710_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_37_LessThan_1845_i16_3_lut_3_lut (.I0(baudrate[2]), .I1(baudrate[3]), 
            .I2(n2728), .I3(GND_net), .O(n16));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46169_4_lut (.I0(n39_adj_5138), .I1(n37), .I2(n35_adj_5137), 
            .I3(n63235), .O(n63231));
    defparam i46169_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46935_2_lut_4_lut (.I0(n2723), .I1(baudrate[8]), .I2(n2727), 
            .I3(baudrate[4]), .O(n63997));
    defparam i46935_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1845_i18_3_lut_3_lut (.I0(baudrate[4]), .I1(baudrate[8]), 
            .I2(n2723), .I3(GND_net), .O(n18));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i18_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_37_LessThan_1845_i20_3_lut_3_lut (.I0(baudrate[5]), .I1(baudrate[6]), 
            .I2(n2725), .I3(GND_net), .O(n20));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i20_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46888_2_lut_4_lut (.I0(n2715), .I1(baudrate[16]), .I2(n2724), 
            .I3(baudrate[7]), .O(n63950));
    defparam i46888_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 div_37_LessThan_1845_i22_3_lut_3_lut (.I0(baudrate[7]), .I1(baudrate[16]), 
            .I2(n2715), .I3(GND_net), .O(n22));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_LessThan_1845_i22_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i49045_4_lut (.I0(n38_adj_5284), .I1(n28_adj_5146), .I2(n41), 
            .I3(n63229), .O(n66107));   // verilog/uart_rx.v(119[33:55])
    defparam i49045_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_37_i2172_1_lut (.I0(baudrate[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n856));   // verilog/uart_rx.v(119[33:55])
    defparam div_37_i2172_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (GND_net, enable_slow_N_4213, clk16MHz, \state_7__N_4110[0] , 
            n29153, ID, n29152, n29143, n29142, n29141, n29140, 
            n29139, n29138, baudrate, n29137, n29136, n29135, n29134, 
            n29133, n29132, n29131, n29130, n29129, n29128, n29127, 
            n29126, n29125, n29124, n29123, n29114, n29113, n29112, 
            n29111, n29110, n29109, n29108, n29107, data_ready, 
            n28925, n55526, n55533, \state_7__N_3918[0] , data, n55524, 
            n57999, n25095, VCC_net, n38386, scl_enable, \state[0] , 
            n29156, scl, sda_enable, sda_out, n29812, n29811, n29810, 
            n29809, n29808, n29806, n29586, n6, n6715, n10, \state_7__N_4126[3] , 
            n38223, n38221, n4, n25100, n4_adj_3) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input GND_net;
    output enable_slow_N_4213;
    input clk16MHz;
    output \state_7__N_4110[0] ;
    input n29153;
    output [7:0]ID;
    input n29152;
    input n29143;
    input n29142;
    input n29141;
    input n29140;
    input n29139;
    input n29138;
    output [31:0]baudrate;
    input n29137;
    input n29136;
    input n29135;
    input n29134;
    input n29133;
    input n29132;
    input n29131;
    input n29130;
    input n29129;
    input n29128;
    input n29127;
    input n29126;
    input n29125;
    input n29124;
    input n29123;
    input n29114;
    input n29113;
    input n29112;
    input n29111;
    input n29110;
    input n29109;
    input n29108;
    input n29107;
    output data_ready;
    input n28925;
    output n55526;
    output n55533;
    input \state_7__N_3918[0] ;
    output [7:0]data;
    output n55524;
    output n57999;
    output n25095;
    input VCC_net;
    output n38386;
    output scl_enable;
    output \state[0] ;
    input n29156;
    output scl;
    output sda_enable;
    output sda_out;
    input n29812;
    input n29811;
    input n29810;
    input n29809;
    input n29808;
    input n29806;
    input n29586;
    input n6;
    output n6715;
    output n10;
    input \state_7__N_4126[3] ;
    output n38223;
    output n38221;
    output n4;
    output n25100;
    output n4_adj_3;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(41[6:14])
    wire [7:0]state;   // verilog/eeprom.v(27[11:16])
    
    wire n4_c, n55527, ready_prev, n21231;
    wire [0:0]n5935;
    
    wire enable;
    wire [15:0]delay_counter_15__N_3956;
    
    wire n27282;
    wire [15:0]delay_counter;   // verilog/eeprom.v(28[12:25])
    
    wire n46759, n6940, n28654, n6942, n6943, n6944, n6945, n6946, 
        enable_slow_N_4212, n38662, n38470, n24974;
    wire [15:0]n5401;
    
    wire n46760;
    wire [2:0]byte_counter;   // verilog/eeprom.v(30[11:23])
    
    wire n66273, n63170;
    wire [7:0]state_7__N_3885;
    
    wire n57974, n50413, n27467, n28892;
    wire [2:0]n17;
    
    wire n29122, n29121, n29120, n29119, n29118, n29117, n29116, 
        n29115, n48526, n48525, n48524, n48523, n48522, n48521, 
        n48520, n48519, n48518, n48517, n48516, n48515, n48514, 
        n48513, n48512, n29813, n54857, n54655, rw, n54799, n4_adj_5008, 
        n63165, n46782, n16, n22, n57940, n20, n24, n49865, 
        n59722;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n55019, n12, n63163, n4_adj_5009, n55531;
    
    SB_LUT4 i1_2_lut (.I0(state[2]), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n4_c));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_4_lut (.I0(n55527), .I1(state[1]), .I2(ready_prev), .I3(n4_c), 
            .O(n21231));
    defparam i2_4_lut.LUT_INIT = 16'hfffb;
    SB_DFF ready_prev_59 (.Q(ready_prev), .C(clk16MHz), .D(enable_slow_N_4213));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFSR enable_58 (.Q(enable), .C(clk16MHz), .D(n5935[0]), .R(state[2]));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(clk16MHz), .E(n27282), 
            .D(delay_counter_15__N_3956[1]), .R(n46759));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(clk16MHz), .E(n27282), 
            .D(delay_counter_15__N_3956[2]), .R(n46759));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(clk16MHz), .E(n27282), 
            .D(delay_counter_15__N_3956[3]), .R(n46759));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(clk16MHz), .E(n27282), 
            .D(n6940), .S(n28654));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(clk16MHz), .E(n27282), 
            .D(delay_counter_15__N_3956[5]), .R(n46759));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(clk16MHz), .E(n27282), 
            .D(n6942), .S(n28654));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(clk16MHz), .E(n27282), 
            .D(n6943), .S(n28654));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(clk16MHz), .E(n27282), 
            .D(n6944), .S(n28654));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(clk16MHz), .E(n27282), 
            .D(n6945), .S(n28654));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(clk16MHz), 
            .E(n27282), .D(n6946), .S(n28654));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i49421_2_lut (.I0(\state_7__N_4110[0] ), .I1(enable_slow_N_4213), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4212));
    defparam i49421_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i22729_2_lut (.I0(state[2]), .I1(n38662), .I2(GND_net), .I3(GND_net), 
            .O(n38470));
    defparam i22729_2_lut.LUT_INIT = 16'h7777;
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(clk16MHz), 
            .E(n27282), .D(delay_counter_15__N_3956[11]), .R(n46759));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(clk16MHz), 
            .E(n27282), .D(delay_counter_15__N_3956[12]), .R(n46759));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(clk16MHz), 
            .E(n27282), .D(delay_counter_15__N_3956[13]), .R(n46759));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(clk16MHz), 
            .E(n27282), .D(delay_counter_15__N_3956[14]), .R(n46759));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i49269_2_lut (.I0(n24974), .I1(enable_slow_N_4213), .I2(GND_net), 
            .I3(GND_net), .O(n5401[9]));
    defparam i49269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_980 (.I0(state[0]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n46760));   // verilog/eeprom.v(35[8] 81[4])
    defparam i1_2_lut_adj_980.LUT_INIT = 16'heeee;
    SB_LUT4 i22917_3_lut (.I0(byte_counter[0]), .I1(byte_counter[2]), .I2(byte_counter[1]), 
            .I3(GND_net), .O(n38662));
    defparam i22917_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i49211_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n66273));   // verilog/eeprom.v(27[11:16])
    defparam i49211_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut (.I0(n46759), .I1(n66273), .I2(n63170), .I3(state[2]), 
            .O(n27282));   // verilog/eeprom.v(27[11:16])
    defparam i1_4_lut.LUT_INIT = 16'hafee;
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(clk16MHz), 
            .E(n27282), .D(delay_counter_15__N_3956[15]), .R(n46759));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFE state_i1 (.Q(state[1]), .C(clk16MHz), .E(n57974), .D(state_7__N_3885[1]));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR byte_counter_2047__i0 (.Q(byte_counter[0]), .C(clk16MHz), 
            .E(n27467), .D(n50413), .R(n28892));   // verilog/eeprom.v(68[25:39])
    SB_DFF bytes_0___i2 (.Q(ID[1]), .C(clk16MHz), .D(n29153));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i3 (.Q(ID[2]), .C(clk16MHz), .D(n29152));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR byte_counter_2047__i2 (.Q(byte_counter[2]), .C(clk16MHz), 
            .E(n27467), .D(n17[2]), .R(n28892));   // verilog/eeprom.v(68[25:39])
    SB_DFFESR byte_counter_2047__i1 (.Q(byte_counter[1]), .C(clk16MHz), 
            .E(n27467), .D(n17[1]), .R(n28892));   // verilog/eeprom.v(68[25:39])
    SB_DFF bytes_0___i4 (.Q(ID[3]), .C(clk16MHz), .D(n29143));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i5 (.Q(ID[4]), .C(clk16MHz), .D(n29142));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i6 (.Q(ID[5]), .C(clk16MHz), .D(n29141));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i7 (.Q(ID[6]), .C(clk16MHz), .D(n29140));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i8 (.Q(ID[7]), .C(clk16MHz), .D(n29139));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i9 (.Q(baudrate[0]), .C(clk16MHz), .D(n29138));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i10 (.Q(baudrate[1]), .C(clk16MHz), .D(n29137));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i11 (.Q(baudrate[2]), .C(clk16MHz), .D(n29136));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i12 (.Q(baudrate[3]), .C(clk16MHz), .D(n29135));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i13 (.Q(baudrate[4]), .C(clk16MHz), .D(n29134));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i14 (.Q(baudrate[5]), .C(clk16MHz), .D(n29133));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i15 (.Q(baudrate[6]), .C(clk16MHz), .D(n29132));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i16 (.Q(baudrate[7]), .C(clk16MHz), .D(n29131));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i17 (.Q(baudrate[8]), .C(clk16MHz), .D(n29130));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i18 (.Q(baudrate[9]), .C(clk16MHz), .D(n29129));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i19 (.Q(baudrate[10]), .C(clk16MHz), .D(n29128));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i20 (.Q(baudrate[11]), .C(clk16MHz), .D(n29127));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i21 (.Q(baudrate[12]), .C(clk16MHz), .D(n29126));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i22 (.Q(baudrate[13]), .C(clk16MHz), .D(n29125));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i23 (.Q(baudrate[14]), .C(clk16MHz), .D(n29124));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i24 (.Q(baudrate[15]), .C(clk16MHz), .D(n29123));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i25 (.Q(baudrate[16]), .C(clk16MHz), .D(n29122));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i26 (.Q(baudrate[17]), .C(clk16MHz), .D(n29121));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i27 (.Q(baudrate[18]), .C(clk16MHz), .D(n29120));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i28 (.Q(baudrate[19]), .C(clk16MHz), .D(n29119));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i29 (.Q(baudrate[20]), .C(clk16MHz), .D(n29118));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i30 (.Q(baudrate[21]), .C(clk16MHz), .D(n29117));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i31 (.Q(baudrate[22]), .C(clk16MHz), .D(n29116));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i32 (.Q(baudrate[23]), .C(clk16MHz), .D(n29115));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i33 (.Q(baudrate[24]), .C(clk16MHz), .D(n29114));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i34 (.Q(baudrate[25]), .C(clk16MHz), .D(n29113));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i35 (.Q(baudrate[26]), .C(clk16MHz), .D(n29112));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i36 (.Q(baudrate[27]), .C(clk16MHz), .D(n29111));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i37 (.Q(baudrate[28]), .C(clk16MHz), .D(n29110));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i38 (.Q(baudrate[29]), .C(clk16MHz), .D(n29109));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i39 (.Q(baudrate[30]), .C(clk16MHz), .D(n29108));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i40 (.Q(baudrate[31]), .C(clk16MHz), .D(n29107));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(clk16MHz), .E(n27282), 
            .D(delay_counter_15__N_3956[0]), .R(n46759));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 add_1198_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n5401[9]), 
            .I3(n48526), .O(delay_counter_15__N_3956[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1198_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n5401[9]), 
            .I3(n48525), .O(delay_counter_15__N_3956[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_16 (.CI(n48525), .I0(delay_counter[14]), .I1(n5401[9]), 
            .CO(n48526));
    SB_LUT4 add_1198_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n5401[9]), 
            .I3(n48524), .O(delay_counter_15__N_3956[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_15 (.CI(n48524), .I0(delay_counter[13]), .I1(n5401[9]), 
            .CO(n48525));
    SB_LUT4 add_1198_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n5401[9]), 
            .I3(n48523), .O(delay_counter_15__N_3956[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_14 (.CI(n48523), .I0(delay_counter[12]), .I1(n5401[9]), 
            .CO(n48524));
    SB_LUT4 add_1198_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n5401[9]), 
            .I3(n48522), .O(delay_counter_15__N_3956[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_13 (.CI(n48522), .I0(delay_counter[11]), .I1(n5401[9]), 
            .CO(n48523));
    SB_LUT4 add_1198_12_lut (.I0(n38470), .I1(delay_counter[10]), .I2(n5401[9]), 
            .I3(n48521), .O(n6946)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_12 (.CI(n48521), .I0(delay_counter[10]), .I1(n5401[9]), 
            .CO(n48522));
    SB_LUT4 add_1198_11_lut (.I0(n38470), .I1(delay_counter[9]), .I2(n5401[9]), 
            .I3(n48520), .O(n6945)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_11 (.CI(n48520), .I0(delay_counter[9]), .I1(n5401[9]), 
            .CO(n48521));
    SB_LUT4 add_1198_10_lut (.I0(n38470), .I1(delay_counter[8]), .I2(n5401[9]), 
            .I3(n48519), .O(n6944)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_10 (.CI(n48519), .I0(delay_counter[8]), .I1(n5401[9]), 
            .CO(n48520));
    SB_LUT4 add_1198_9_lut (.I0(n38470), .I1(delay_counter[7]), .I2(n5401[9]), 
            .I3(n48518), .O(n6943)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_9 (.CI(n48518), .I0(delay_counter[7]), .I1(n5401[9]), 
            .CO(n48519));
    SB_LUT4 add_1198_8_lut (.I0(n38470), .I1(delay_counter[6]), .I2(n5401[9]), 
            .I3(n48517), .O(n6942)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_8 (.CI(n48517), .I0(delay_counter[6]), .I1(n5401[9]), 
            .CO(n48518));
    SB_LUT4 add_1198_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n5401[9]), 
            .I3(n48516), .O(delay_counter_15__N_3956[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_7 (.CI(n48516), .I0(delay_counter[5]), .I1(n5401[9]), 
            .CO(n48517));
    SB_LUT4 add_1198_6_lut (.I0(n38470), .I1(delay_counter[4]), .I2(n5401[9]), 
            .I3(n48515), .O(n6940)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1198_6 (.CI(n48515), .I0(delay_counter[4]), .I1(n5401[9]), 
            .CO(n48516));
    SB_LUT4 add_1198_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n5401[9]), 
            .I3(n48514), .O(delay_counter_15__N_3956[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_5 (.CI(n48514), .I0(delay_counter[3]), .I1(n5401[9]), 
            .CO(n48515));
    SB_LUT4 add_1198_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n5401[9]), 
            .I3(n48513), .O(delay_counter_15__N_3956[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_4 (.CI(n48513), .I0(delay_counter[2]), .I1(n5401[9]), 
            .CO(n48514));
    SB_LUT4 add_1198_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n5401[9]), 
            .I3(n48512), .O(delay_counter_15__N_3956[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_3 (.CI(n48512), .I0(delay_counter[1]), .I1(n5401[9]), 
            .CO(n48513));
    SB_LUT4 add_1198_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n5401[9]), 
            .I3(GND_net), .O(delay_counter_15__N_3956[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1198_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1198_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n5401[9]), 
            .CO(n48512));
    SB_DFF state_i2 (.Q(state[2]), .C(clk16MHz), .D(n29813));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF state_i0 (.Q(state[0]), .C(clk16MHz), .D(n54857));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF rw_64 (.Q(rw), .C(clk16MHz), .D(n54655));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF data_ready_61 (.Q(data_ready), .C(clk16MHz), .D(n54799));   // verilog/eeprom.v(35[8] 81[4])
    SB_DFF bytes_0___i1 (.Q(ID[0]), .C(clk16MHz), .D(n28925));   // verilog/eeprom.v(35[8] 81[4])
    SB_LUT4 i32374_2_lut_3_lut_4_lut (.I0(ready_prev), .I1(enable_slow_N_4213), 
            .I2(byte_counter[0]), .I3(byte_counter[1]), .O(n17[1]));   // verilog/eeprom.v(68[25:39])
    defparam i32374_2_lut_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(byte_counter[0]), .I1(n21231), .I2(byte_counter[1]), 
            .I3(byte_counter[2]), .O(n55526));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_981 (.I0(byte_counter[1]), .I1(byte_counter[2]), 
            .I2(n21231), .I3(byte_counter[0]), .O(n55533));   // verilog/eeprom.v(66[9:28])
    defparam i1_2_lut_3_lut_4_lut_adj_981.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_4_lut_adj_982 (.I0(state[2]), .I1(state[1]), .I2(\state_7__N_3918[0] ), 
            .I3(state[0]), .O(n4_adj_5008));
    defparam i1_4_lut_adj_982.LUT_INIT = 16'hbbba;
    SB_LUT4 i47070_3_lut (.I0(n55527), .I1(n24974), .I2(state[1]), .I3(GND_net), 
            .O(n63165));
    defparam i47070_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i2_4_lut_adj_983 (.I0(n63165), .I1(n4_adj_5008), .I2(n46782), 
            .I3(state[0]), .O(n57974));
    defparam i2_4_lut_adj_983.LUT_INIT = 16'hcfee;
    SB_LUT4 i3_2_lut (.I0(delay_counter[7]), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(GND_net), .O(n16));   // verilog/eeprom.v(55[12:28])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut (.I0(delay_counter[1]), .I1(delay_counter[6]), .I2(delay_counter[2]), 
            .I3(delay_counter[12]), .O(n22));   // verilog/eeprom.v(55[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut (.I0(delay_counter[9]), .I1(delay_counter[14]), .I2(delay_counter[11]), 
            .I3(delay_counter[15]), .O(n57940));   // verilog/eeprom.v(55[12:28])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6668_4_lut (.I0(state[1]), .I1(n38662), .I2(state[2]), .I3(state[0]), 
            .O(state_7__N_3885[1]));   // verilog/eeprom.v(38[3] 80[10])
    defparam i6668_4_lut.LUT_INIT = 16'ha5ba;
    SB_LUT4 i7_3_lut (.I0(delay_counter[8]), .I1(delay_counter[4]), .I2(delay_counter[13]), 
            .I3(GND_net), .O(n20));   // verilog/eeprom.v(55[12:28])
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n57940), .I1(n22), .I2(n16), .I3(delay_counter[0]), 
            .O(n24));   // verilog/eeprom.v(55[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(delay_counter[5]), .I1(n24), .I2(n20), .I3(delay_counter[10]), 
            .O(n24974));   // verilog/eeprom.v(55[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(state[0]), .I1(n24974), .I2(enable_slow_N_4213), 
            .I3(GND_net), .O(n49865));
    defparam i2_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i13_4_lut (.I0(data_ready), .I1(state[2]), .I2(n46760), .I3(n38662), 
            .O(n54799));   // verilog/eeprom.v(27[11:16])
    defparam i13_4_lut.LUT_INIT = 16'haca8;
    SB_LUT4 i42673_3_lut (.I0(state[2]), .I1(n49865), .I2(state[1]), .I3(GND_net), 
            .O(n59722));
    defparam i42673_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_4_lut_adj_984 (.I0(rw), .I1(saved_addr[0]), .I2(n55527), 
            .I3(\state_7__N_4110[0] ), .O(n55019));   // verilog/i2c_controller.v(33[12:17])
    defparam i1_4_lut_adj_984.LUT_INIT = 16'hcacc;
    SB_LUT4 i30_4_lut (.I0(\state_7__N_3918[0] ), .I1(n24974), .I2(state[1]), 
            .I3(n55527), .O(n12));
    defparam i30_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i29_4_lut (.I0(n12), .I1(n63163), .I2(state[0]), .I3(state[2]), 
            .O(n54857));
    defparam i29_4_lut.LUT_INIT = 16'hf0ca;
    SB_LUT4 i1_4_lut_adj_985 (.I0(state[1]), .I1(state[0]), .I2(n46782), 
            .I3(state[2]), .O(n29813));
    defparam i1_4_lut_adj_985.LUT_INIT = 16'hee08;
    SB_LUT4 i47068_2_lut_3_lut (.I0(ready_prev), .I1(enable_slow_N_4213), 
            .I2(state[1]), .I3(GND_net), .O(n63163));
    defparam i47068_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i11_4_lut_4_lut (.I0(rw), .I1(state[1]), .I2(state[0]), .I3(n59722), 
            .O(n54655));   // verilog/eeprom.v(27[11:16])
    defparam i11_4_lut_4_lut.LUT_INIT = 16'haace;
    SB_LUT4 i19670_3_lut_4_lut (.I0(state[0]), .I1(n24974), .I2(enable_slow_N_4213), 
            .I3(state[1]), .O(n5935[0]));   // verilog/eeprom.v(27[11:16])
    defparam i19670_3_lut_4_lut.LUT_INIT = 16'h10aa;
    SB_LUT4 i13270_3_lut_4_lut (.I0(n4_adj_5009), .I1(n55531), .I2(data[7]), 
            .I3(baudrate[23]), .O(n29115));
    defparam i13270_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13271_3_lut_4_lut (.I0(n4_adj_5009), .I1(n55531), .I2(data[6]), 
            .I3(baudrate[22]), .O(n29116));
    defparam i13271_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_4_lut (.I0(state[0]), .I1(n38662), .I2(state[2]), 
            .I3(state[1]), .O(n46759));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h001a;
    SB_LUT4 i12810_2_lut_4_lut (.I0(state[0]), .I1(n38662), .I2(state[2]), 
            .I3(n27282), .O(n28654));
    defparam i12810_2_lut_4_lut.LUT_INIT = 16'h3a00;
    SB_LUT4 i13272_3_lut_4_lut (.I0(n4_adj_5009), .I1(n55531), .I2(data[5]), 
            .I3(baudrate[21]), .O(n29117));
    defparam i13272_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13273_3_lut_4_lut (.I0(n4_adj_5009), .I1(n55531), .I2(data[4]), 
            .I3(baudrate[20]), .O(n29118));
    defparam i13273_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13274_3_lut_4_lut (.I0(n4_adj_5009), .I1(n55531), .I2(data[3]), 
            .I3(baudrate[19]), .O(n29119));
    defparam i13274_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13275_3_lut_4_lut (.I0(n4_adj_5009), .I1(n55531), .I2(data[2]), 
            .I3(baudrate[18]), .O(n29120));
    defparam i13275_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13276_3_lut_4_lut (.I0(n4_adj_5009), .I1(n55531), .I2(data[1]), 
            .I3(baudrate[17]), .O(n29121));
    defparam i13276_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13277_3_lut_4_lut (.I0(n4_adj_5009), .I1(n55531), .I2(data[0]), 
            .I3(baudrate[16]), .O(n29122));
    defparam i13277_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut (.I0(ready_prev), .I1(enable_slow_N_4213), .I2(byte_counter[0]), 
            .I3(GND_net), .O(n50413));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hb4b4;
    SB_LUT4 i1_4_lut_4_lut_adj_986 (.I0(state[2]), .I1(\state_7__N_3918[0] ), 
            .I2(state[0]), .I3(state[1]), .O(n27467));
    defparam i1_4_lut_4_lut_adj_986.LUT_INIT = 16'h5004;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state_7__N_3918[0] ), .I1(state[0]), .I2(state[1]), 
            .I3(state[2]), .O(n28892));   // verilog/eeprom.v(68[25:39])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i47084_2_lut_3_lut (.I0(n38662), .I1(state[0]), .I2(state[1]), 
            .I3(GND_net), .O(n63170));   // verilog/eeprom.v(27[11:16])
    defparam i47084_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 equal_323_i4_2_lut (.I0(byte_counter[1]), .I1(byte_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5009));   // verilog/eeprom.v(66[9:28])
    defparam equal_323_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_987 (.I0(byte_counter[1]), .I1(byte_counter[2]), 
            .I2(n21231), .I3(byte_counter[0]), .O(n55524));   // verilog/eeprom.v(66[9:28])
    defparam i1_2_lut_3_lut_4_lut_adj_987.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_988 (.I0(byte_counter[0]), .I1(n21231), .I2(byte_counter[2]), 
            .I3(byte_counter[1]), .O(n57999));
    defparam i2_3_lut_4_lut_adj_988.LUT_INIT = 16'hffef;
    SB_LUT4 i32381_3_lut_4_lut (.I0(n46782), .I1(byte_counter[0]), .I2(byte_counter[1]), 
            .I3(byte_counter[2]), .O(n17[2]));   // verilog/eeprom.v(68[25:39])
    defparam i32381_3_lut_4_lut.LUT_INIT = 16'hbf40;
    SB_LUT4 i1_2_lut_adj_989 (.I0(n21231), .I1(byte_counter[0]), .I2(GND_net), 
            .I3(GND_net), .O(n55531));
    defparam i1_2_lut_adj_989.LUT_INIT = 16'hbbbb;
    i2c_controller i2c (.n25095(n25095), .GND_net(GND_net), .VCC_net(VCC_net), 
            .n38386(n38386), .clk16MHz(clk16MHz), .scl_enable(scl_enable), 
            .enable_slow_N_4212(enable_slow_N_4212), .\state_7__N_4110[0] (\state_7__N_4110[0] ), 
            .\state[0] (\state[0] ), .n29156(n29156), .data({data}), .scl(scl), 
            .sda_enable(sda_enable), .sda_out(sda_out), .n29812(n29812), 
            .n29811(n29811), .n29810(n29810), .n29809(n29809), .n29808(n29808), 
            .n29806(n29806), .n29586(n29586), .n6(n6), .n55019(n55019), 
            .\saved_addr[0] (saved_addr[0]), .n6715(n6715), .n10(n10), 
            .ready_prev(ready_prev), .enable_slow_N_4213(enable_slow_N_4213), 
            .n46782(n46782), .\state_7__N_4126[3] (\state_7__N_4126[3] ), 
            .enable(enable), .n38223(n38223), .n38221(n38221), .n4(n4), 
            .n25100(n25100), .n4_adj_2(n4_adj_3), .n55527(n55527)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(83[16] 97[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (n25095, GND_net, VCC_net, n38386, clk16MHz, 
            scl_enable, enable_slow_N_4212, \state_7__N_4110[0] , \state[0] , 
            n29156, data, scl, sda_enable, sda_out, n29812, n29811, 
            n29810, n29809, n29808, n29806, n29586, n6, n55019, 
            \saved_addr[0] , n6715, n10, ready_prev, enable_slow_N_4213, 
            n46782, \state_7__N_4126[3] , enable, n38223, n38221, 
            n4, n25100, n4_adj_2, n55527) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output n25095;
    input GND_net;
    input VCC_net;
    output n38386;
    input clk16MHz;
    output scl_enable;
    input enable_slow_N_4212;
    output \state_7__N_4110[0] ;
    output \state[0] ;
    input n29156;
    output [7:0]data;
    output scl;
    output sda_enable;
    output sda_out;
    input n29812;
    input n29811;
    input n29810;
    input n29809;
    input n29808;
    input n29806;
    input n29586;
    input n6;
    input n55019;
    output \saved_addr[0] ;
    output n6715;
    output n10;
    input ready_prev;
    output enable_slow_N_4213;
    output n46782;
    input \state_7__N_4126[3] ;
    input enable;
    output n38223;
    output n38221;
    output n4;
    output n25100;
    output n4_adj_2;
    output n55527;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(41[6:14])
    
    wire n15;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n49287, n49286, n49285, n49284, n49283, i2c_clk_N_4199, 
        scl_enable_N_4200, n27356, n28648;
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    wire n58134, n27336, n54735, n57461, n27334, sda_out_adj_4998;
    wire [7:0]n119;
    
    wire n27393, n28597, n48533, n48532, n48531, n48530, n48529, 
        n48528, n48527, n5, n38677, n38524, n38675, n58283, n57985, 
        n58196, n6708, n63164, n56496, n28, n66283, n11, n56380;
    wire [1:0]n6784;
    
    wire n10_adj_4999, n11_adj_5000, n11_adj_5001, n4_c, n11_adj_5002, 
        n10_adj_5003, n11_adj_5004, state_7__N_4109, n15_adj_5007;
    
    SB_LUT4 i1_2_lut (.I0(n15), .I1(counter[0]), .I2(GND_net), .I3(GND_net), 
            .O(n25095));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 counter2_2057_2058_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n49287), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_2057_2058_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n49286), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_6 (.CI(n49286), .I0(GND_net), .I1(counter2[4]), 
            .CO(n49287));
    SB_LUT4 counter2_2057_2058_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n49285), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_5 (.CI(n49285), .I0(GND_net), .I1(counter2[3]), 
            .CO(n49286));
    SB_LUT4 counter2_2057_2058_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n49284), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_4 (.CI(n49284), .I0(GND_net), .I1(counter2[2]), 
            .CO(n49285));
    SB_LUT4 counter2_2057_2058_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n49283), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2057_2058_add_4_3 (.CI(n49283), .I0(GND_net), .I1(counter2[1]), 
            .CO(n49284));
    SB_LUT4 counter2_2057_2058_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2057_2058_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22645_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n38386));
    defparam i22645_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter2_2057_2058_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n49283));
    SB_DFF i2c_clk_122 (.Q(i2c_clk), .C(clk16MHz), .D(i2c_clk_N_4199));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_124 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4200));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_DFFE enable_slow_121 (.Q(\state_7__N_4110[0] ), .C(clk16MHz), .E(n27356), 
            .D(enable_slow_N_4212));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFSR counter2_2057_2058__i1 (.Q(counter2[0]), .C(clk16MHz), .D(n29[0]), 
            .R(n28648));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 i22602_3_lut_4_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(state[2]), 
            .I3(state[3]), .O(scl_enable_N_4200));   // verilog/i2c_controller.v(44[32:47])
    defparam i22602_3_lut_4_lut_4_lut.LUT_INIT = 16'hfefc;
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n29156));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i22537_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i22537_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFNESS write_enable_132 (.Q(sda_enable), .C(i2c_clk), .E(n27336), 
            .D(n58134), .S(n54735));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFNESS sda_out_133 (.Q(sda_out_adj_4998), .C(i2c_clk), .E(n27334), 
            .D(n57461), .S(n54735));   // verilog/i2c_controller.v(180[12] 218[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n27393), .D(n119[0]), 
            .S(n28597));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i2555_2_lut (.I0(sda_out_adj_4998), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n48533), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n48532), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n48532), .I0(counter[6]), .I1(VCC_net), 
            .CO(n48533));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n48531), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n48531), .I0(counter[5]), .I1(VCC_net), 
            .CO(n48532));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n48530), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n48530), .I0(counter[4]), .I1(VCC_net), 
            .CO(n48531));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n48529), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n48529), .I0(counter[3]), .I1(VCC_net), 
            .CO(n48530));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n48528), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n48528), .I0(counter[2]), .I1(VCC_net), 
            .CO(n48529));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n48527), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n48527), .I0(counter[1]), .I1(VCC_net), 
            .CO(n48528));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n48527));
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n29812));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n29811));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n29810));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n29809));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n29808));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n29806));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n29586));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n6));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n55019));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n27393), .D(n119[1]), 
            .S(n28597));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n27393), .D(n119[2]), 
            .S(n28597));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n27393), .D(n119[3]), 
            .R(n28597));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n27393), .D(n119[4]), 
            .R(n28597));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n27393), .D(n119[5]), 
            .R(n28597));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n27393), .D(n119[6]), 
            .R(n28597));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n27393), .D(n119[7]), 
            .R(n28597));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i1 (.Q(state[1]), .C(i2c_clk), .E(n6715), .D(n5), 
            .S(n38677));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(state[2]), .C(i2c_clk), .E(n6715), .D(n38524), 
            .S(n38675));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(state[3]), .C(i2c_clk), .E(n6715), .D(n58283), 
            .S(n57985));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_2057_2058__i2 (.Q(counter2[1]), .C(clk16MHz), .D(n29[1]), 
            .R(n28648));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i3 (.Q(counter2[2]), .C(clk16MHz), .D(n29[2]), 
            .R(n28648));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i4 (.Q(counter2[3]), .C(clk16MHz), .D(n29[3]), 
            .R(n28648));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i5 (.Q(counter2[4]), .C(clk16MHz), .D(n29[4]), 
            .R(n28648));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2057_2058__i6 (.Q(counter2[5]), .C(clk16MHz), .D(n29[5]), 
            .R(n28648));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(n10), .I1(counter[5]), .I2(counter[3]), .I3(counter[4]), 
            .O(n58196));   // verilog/i2c_controller.v(110[10:22])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n58196), .I2(counter[7]), .I3(counter[0]), 
            .O(n6708));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_967 (.I0(n27393), .I1(\state[0] ), .I2(state[2]), 
            .I3(state[3]), .O(n28597));
    defparam i3_4_lut_adj_967.LUT_INIT = 16'h0008;
    SB_LUT4 i1_4_lut (.I0(state[3]), .I1(n63164), .I2(n56496), .I3(\state[0] ), 
            .O(n27393));
    defparam i1_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i1_4_lut_adj_968 (.I0(state[3]), .I1(state[1]), .I2(\state[0] ), 
            .I3(state[2]), .O(n28));
    defparam i1_4_lut_adj_968.LUT_INIT = 16'h5110;
    SB_LUT4 i49221_2_lut (.I0(state[3]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(n66283));
    defparam i49221_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_969 (.I0(n11), .I1(n66283), .I2(n28), .I3(n56380), 
            .O(n27334));
    defparam i1_4_lut_adj_969.LUT_INIT = 16'ha0a8;
    SB_LUT4 mux_1830_Mux_1_i7_4_lut (.I0(counter[1]), .I1(counter[0]), .I2(counter[2]), 
            .I3(\saved_addr[0] ), .O(n6784[1]));   // verilog/i2c_controller.v(201[28:35])
    defparam mux_1830_Mux_1_i7_4_lut.LUT_INIT = 16'hc1c0;
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_adj_4999));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_adj_4999), .I2(counter2[0]), 
            .I3(GND_net), .O(n28648));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_970 (.I0(i2c_clk), .I1(n28648), .I2(GND_net), 
            .I3(GND_net), .O(i2c_clk_N_4199));
    defparam i1_2_lut_adj_970.LUT_INIT = 16'h6666;
    SB_LUT4 i39373_2_lut (.I0(state[2]), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n56380));
    defparam i39373_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_971 (.I0(n11), .I1(n56380), .I2(state[3]), .I3(state[1]), 
            .O(n54735));
    defparam i3_4_lut_adj_971.LUT_INIT = 16'h0020;
    SB_LUT4 i1_4_lut_adj_972 (.I0(n11), .I1(state[1]), .I2(state[3]), 
            .I3(n56380), .O(n27336));
    defparam i1_4_lut_adj_972.LUT_INIT = 16'h0a22;
    SB_LUT4 state_7__I_0_142_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(state[3]), .I3(state[2]), .O(n11_adj_5000));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_142_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_2_lut_adj_973 (.I0(ready_prev), .I1(enable_slow_N_4213), 
            .I2(GND_net), .I3(GND_net), .O(n46782));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i1_2_lut_adj_973.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_4_lut_adj_974 (.I0(\state_7__N_4126[3] ), .I1(n11_adj_5001), 
            .I2(n11), .I3(enable), .O(n4_c));
    defparam i1_4_lut_adj_974.LUT_INIT = 16'h2a2f;
    SB_LUT4 i49342_3_lut (.I0(n6715), .I1(n15), .I2(n11_adj_5000), .I3(GND_net), 
            .O(n38675));
    defparam i49342_3_lut.LUT_INIT = 16'h2a2a;
    SB_LUT4 i49358_2_lut (.I0(\state_7__N_4126[3] ), .I1(n11_adj_5001), 
            .I2(GND_net), .I3(GND_net), .O(n38524));
    defparam i49358_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_4_lut_adj_975 (.I0(n11_adj_5002), .I1(n11_adj_5001), .I2(\saved_addr[0] ), 
            .I3(\state_7__N_4126[3] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_975.LUT_INIT = 16'h5575;
    SB_LUT4 i1_2_lut_adj_976 (.I0(state[3]), .I1(state[2]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_5003));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_976.LUT_INIT = 16'hdddd;
    SB_LUT4 i22483_2_lut (.I0(n11_adj_5004), .I1(n11_adj_5000), .I2(GND_net), 
            .I3(GND_net), .O(n38223));
    defparam i22483_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49237_4_lut (.I0(state_7__N_4109), .I1(n6708), .I2(n11_adj_5004), 
            .I3(n38221), .O(n6715));
    defparam i49237_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 equal_355_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_355_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_977 (.I0(counter[0]), .I1(n15), .I2(GND_net), 
            .I3(GND_net), .O(n25100));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i1_2_lut_adj_977.LUT_INIT = 16'heeee;
    SB_LUT4 equal_353_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_2));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_353_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i49344_3_lut_4_lut (.I0(n6715), .I1(n15_adj_5007), .I2(n11_adj_5004), 
            .I3(n11_adj_5000), .O(n38677));
    defparam i49344_3_lut_4_lut.LUT_INIT = 16'h2aaa;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[3]), .I1(state[1]), .I2(state[2]), 
            .I3(\state[0] ), .O(n58134));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h1110;
    SB_LUT4 i2_3_lut_4_lut_adj_978 (.I0(\state[0] ), .I1(state[1]), .I2(n10_adj_5003), 
            .I3(n4_c), .O(n58283));   // verilog/i2c_controller.v(151[5:14])
    defparam i2_3_lut_4_lut_adj_978.LUT_INIT = 16'hff04;
    SB_LUT4 state_7__I_0_144_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(state[2]), .I3(state[3]), .O(n15));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_144_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 i49334_3_lut_4_lut (.I0(state[3]), .I1(state[2]), .I2(n6715), 
            .I3(state[1]), .O(n57985));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i49334_3_lut_4_lut.LUT_INIT = 16'h0040;
    SB_LUT4 i22884_2_lut_3_lut (.I0(state[3]), .I1(state[2]), .I2(\state[0] ), 
            .I3(GND_net), .O(n38221));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i22884_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 equal_276_i11_2_lut_3_lut_4_lut (.I0(state[2]), .I1(state[3]), 
            .I2(state[1]), .I3(\state[0] ), .O(n15_adj_5007));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam equal_276_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_3_lut_4_lut_adj_979 (.I0(state[2]), .I1(state[3]), .I2(n6784[1]), 
            .I3(state[1]), .O(n57461));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i2_3_lut_4_lut_adj_979.LUT_INIT = 16'h1000;
    SB_LUT4 i49429_2_lut_3_lut_4_lut (.I0(state[2]), .I1(state[3]), .I2(state[1]), 
            .I3(\state[0] ), .O(enable_slow_N_4213));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam i49429_2_lut_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 state_7__I_0_140_i11_2_lut_3_lut_4_lut (.I0(state[2]), .I1(state[3]), 
            .I2(\state[0] ), .I3(state[1]), .O(n11_adj_5001));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam state_7__I_0_140_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(state[2]), .I1(state[3]), 
            .I2(state[1]), .I3(\state[0] ), .O(n11_adj_5004));   // verilog/i2c_controller.v(181[4] 217[11])
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i39365_3_lut_4_lut (.I0(state[2]), .I1(state[1]), .I2(\state[0] ), 
            .I3(state[3]), .O(n55527));
    defparam i39365_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47069_2_lut_3_lut (.I0(state[2]), .I1(state[1]), .I2(n6708), 
            .I3(GND_net), .O(n63164));
    defparam i47069_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i22882_3_lut_4_lut (.I0(state[1]), .I1(\state[0] ), .I2(state[2]), 
            .I3(state[3]), .O(state_7__N_4109));
    defparam i22882_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 equal_1562_i11_2_lut_3_lut_4_lut (.I0(state[1]), .I1(\state[0] ), 
            .I2(state[2]), .I3(state[3]), .O(n11));
    defparam equal_1562_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut (.I0(enable), .I1(\state_7__N_4110[0] ), .I2(enable_slow_N_4213), 
            .I3(GND_net), .O(n27356));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 state_7__I_0_145_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), 
            .I2(state[2]), .I3(state[3]), .O(n11_adj_5002));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_145_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i39488_3_lut_4_lut (.I0(\state[0] ), .I1(state[1]), .I2(\state_7__N_4126[3] ), 
            .I3(state[2]), .O(n56496));   // verilog/i2c_controller.v(77[27:43])
    defparam i39488_3_lut_4_lut.LUT_INIT = 16'hffd0;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (n2882, pwm_out, clk32MHz, GND_net, VCC_net, pwm_setpoint, 
            reset) /* synthesis syn_module_defined=1 */ ;
    input n2882;
    output pwm_out;
    input clk32MHz;
    input GND_net;
    input VCC_net;
    input [23:0]pwm_setpoint;
    input reset;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(41[16:24])
    
    wire pwm_out_N_577, n53897;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n49141, n48, n53939, n49140, n53967, n49139, n54001, 
        n49138, n54043, n49137, n54085, n49136, n54117, n49135, 
        n54153, n49134, n54189, n49133, n54225, n49132, n54253, 
        n49131, n54289, n49130, n54325, n49129, n54369, n49128, 
        n54415, n49127, n54459, n49126, n54513, n49125, n54567, 
        n49124, n54699, n49123, n54841, n49122, n54963, n49121, 
        n54961, n49120, n54959, n49119, n54939, n41, n39, n45, 
        n37, n43, n29, n31, n23, n25, n35, n33, n11, n13, 
        n15, n27, n9, n17, n19, n21, n63920, n63894, n12, 
        n30, n63965, n64899, n64887, n65933, n65327, n66070, n6, 
        n65663, n65664, n16, n24, n63622, n8, n63614, n65453, 
        n64306, n4, n65667, n65668, n63789, n10, n63739, n65937, 
        n64302, n66202, n66203, n66112, n63661, n65775, n65456, 
        n66015, n57984, n22, n15_adj_4995, n20, n24_adj_4996, n19_adj_4997;
    
    SB_DFFE pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .E(n2882), .D(pwm_out_N_577));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 pwm_counter_2040_add_4_25_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n49141), .O(n53897)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 pwm_counter_2040_add_4_24_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n49140), .O(n53939)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_24 (.CI(n49140), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n49141));
    SB_LUT4 pwm_counter_2040_add_4_23_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n49139), .O(n53967)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_23 (.CI(n49139), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n49140));
    SB_LUT4 pwm_counter_2040_add_4_22_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n49138), .O(n54001)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_22 (.CI(n49138), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n49139));
    SB_LUT4 pwm_counter_2040_add_4_21_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n49137), .O(n54043)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_21 (.CI(n49137), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n49138));
    SB_LUT4 pwm_counter_2040_add_4_20_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n49136), .O(n54085)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_20 (.CI(n49136), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n49137));
    SB_LUT4 pwm_counter_2040_add_4_19_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n49135), .O(n54117)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_19 (.CI(n49135), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n49136));
    SB_LUT4 pwm_counter_2040_add_4_18_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n49134), .O(n54153)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_18 (.CI(n49134), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n49135));
    SB_LUT4 pwm_counter_2040_add_4_17_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n49133), .O(n54189)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_17 (.CI(n49133), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n49134));
    SB_LUT4 pwm_counter_2040_add_4_16_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n49132), .O(n54225)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_16 (.CI(n49132), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n49133));
    SB_LUT4 pwm_counter_2040_add_4_15_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n49131), .O(n54253)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_15 (.CI(n49131), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n49132));
    SB_LUT4 pwm_counter_2040_add_4_14_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n49130), .O(n54289)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_14 (.CI(n49130), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n49131));
    SB_LUT4 pwm_counter_2040_add_4_13_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n49129), .O(n54325)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_13 (.CI(n49129), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n49130));
    SB_LUT4 pwm_counter_2040_add_4_12_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n49128), .O(n54369)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_12 (.CI(n49128), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n49129));
    SB_LUT4 pwm_counter_2040_add_4_11_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n49127), .O(n54415)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_11 (.CI(n49127), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n49128));
    SB_LUT4 pwm_counter_2040_add_4_10_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n49126), .O(n54459)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_10 (.CI(n49126), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n49127));
    SB_LUT4 pwm_counter_2040_add_4_9_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n49125), .O(n54513)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_9 (.CI(n49125), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n49126));
    SB_LUT4 pwm_counter_2040_add_4_8_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n49124), .O(n54567)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_8 (.CI(n49124), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n49125));
    SB_LUT4 pwm_counter_2040_add_4_7_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n49123), .O(n54699)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_7 (.CI(n49123), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n49124));
    SB_LUT4 pwm_counter_2040_add_4_6_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n49122), .O(n54841)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_6 (.CI(n49122), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n49123));
    SB_LUT4 pwm_counter_2040_add_4_5_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n49121), .O(n54963)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_5 (.CI(n49121), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n49122));
    SB_LUT4 pwm_counter_2040_add_4_4_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n49120), .O(n54961)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_4 (.CI(n49120), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n49121));
    SB_LUT4 pwm_counter_2040_add_4_3_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n49119), .O(n54959)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_3 (.CI(n49119), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n49120));
    SB_LUT4 pwm_counter_2040_add_4_2_lut (.I0(n48), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n54939)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2040_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY pwm_counter_2040_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n49119));
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(pwm_counter[22]), .I1(pwm_setpoint[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46858_4_lut (.I0(n21), .I1(n19), .I2(n17), .I3(n9), .O(n63920));
    defparam i46858_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46832_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11), .O(n63894));
    defparam i46832_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47837_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n63965), 
            .O(n64899));
    defparam i47837_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i47825_4_lut (.I0(n19), .I1(n17), .I2(n15), .I3(n64899), 
            .O(n64887));
    defparam i47825_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i48871_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n64887), 
            .O(n65933));
    defparam i48871_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48265_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n65933), 
            .O(n65327));
    defparam i48265_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i49008_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n65327), 
            .O(n66070));
    defparam i49008_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48601_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n65663));   // verilog/pwm.v(21[8:24])
    defparam i48601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48602_3_lut (.I0(n65663), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n65664));   // verilog/pwm.v(21[8:24])
    defparam i48602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46560_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n63920), 
            .O(n63622));
    defparam i46560_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48391_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n63614), 
            .O(n65453));   // verilog/pwm.v(21[8:24])
    defparam i48391_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47244_3_lut (.I0(n65664), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n64306));   // verilog/pwm.v(21[8:24])
    defparam i47244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_counter[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_setpoint[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i48605_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n65667));   // verilog/pwm.v(21[8:24])
    defparam i48605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48606_3_lut (.I0(n65667), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n65668));   // verilog/pwm.v(21[8:24])
    defparam i48606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46727_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n63894), 
            .O(n63789));
    defparam i46727_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48875_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n63739), 
            .O(n65937));   // verilog/pwm.v(21[8:24])
    defparam i48875_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47240_3_lut (.I0(n65668), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n64302));   // verilog/pwm.v(21[8:24])
    defparam i47240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49140_4_lut (.I0(n64302), .I1(n65937), .I2(n35), .I3(n63789), 
            .O(n66202));   // verilog/pwm.v(21[8:24])
    defparam i49140_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49141_3_lut (.I0(n66202), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n66203));   // verilog/pwm.v(21[8:24])
    defparam i49141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49050_3_lut (.I0(n66203), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n66112));   // verilog/pwm.v(21[8:24])
    defparam i49050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46599_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n66070), 
            .O(n63661));
    defparam i46599_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48713_4_lut (.I0(n64306), .I1(n65453), .I2(n45), .I3(n63622), 
            .O(n65775));   // verilog/pwm.v(21[8:24])
    defparam i48713_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48394_3_lut (.I0(n66112), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n65456));   // verilog/pwm.v(21[8:24])
    defparam i48394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48953_4_lut (.I0(n65456), .I1(n65775), .I2(n45), .I3(n63661), 
            .O(n66015));   // verilog/pwm.v(21[8:24])
    defparam i48953_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48954_3_lut (.I0(n66015), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_577));   // verilog/pwm.v(21[8:24])
    defparam i48954_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFR pwm_counter_2040__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n54939), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n54959), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n54961), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n54963), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n54841), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n54699), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n54567), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n54513), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n54459), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n54415), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n54369), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n54325), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n54289), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n54253), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n54225), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n54189), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n54153), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n54117), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n54085), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n54043), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n54001), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n53967), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n53939), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_DFFR pwm_counter_2040__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n53897), 
            .R(reset));   // verilog/pwm.v(17[20:33])
    SB_LUT4 i46903_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n63965));   // verilog/pwm.v(21[8:24])
    defparam i46903_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n57984));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_4_lut (.I0(pwm_counter[22]), .I1(pwm_counter[15]), .I2(pwm_counter[18]), 
            .I3(pwm_counter[16]), .O(n22));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n57984), .I1(pwm_counter[12]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n15_adj_4995));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i7_3_lut (.I0(pwm_counter[17]), .I1(pwm_counter[21]), .I2(pwm_counter[11]), 
            .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n15_adj_4995), .I1(n22), .I2(pwm_counter[20]), 
            .I3(pwm_counter[13]), .O(n24_adj_4996));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(pwm_counter[19]), .I1(pwm_counter[14]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4997));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(pwm_counter[23]), .I1(n19_adj_4997), .I2(n24_adj_4996), 
            .I3(n20), .O(n48));   // verilog/pwm.v(17[20:33])
    defparam i1_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46552_2_lut_4_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n63614));
    defparam i46552_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[21]), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46677_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n63739));
    defparam i46677_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, \Ki[2] , n335, setpoint, deadband, \Ki[3] , 
            \Kp[7] , IntegralLimit, \Kp[1] , \Kp[0] , \Ki[4] , \Ki[5] , 
            \Kp[2] , \Kp[3] , \Kp[4] , \Kp[5] , \Kp[6] , \Kp[8] , 
            \Kp[9] , \Kp[10] , \Kp[11] , \Kp[12] , \Kp[13] , \Kp[14] , 
            \Ki[6] , \Kp[15] , \encoder1_position_scaled[0] , n15, n62934, 
            n15_adj_1, \encoder1_position_scaled[1] , n62948, \motor_state[9] , 
            control_update, duty, clk16MHz, reset, \motor_state[8] , 
            \Ki[1] , \Ki[0] , PWMLimit, \Ki[7] , \Ki[8] , \Ki[9] , 
            \motor_state[7] , VCC_net, \motor_state[6] , \Ki[10] , \Ki[11] , 
            \Ki[12] , \Ki[13] , \motor_state[5] , \Ki[14] , \Ki[15] , 
            \motor_state[4] , \motor_state[10] , \motor_state[3] , n3, 
            control_mode, n55181, n105, n7064, n38638, n29778, \PID_CONTROLLER.integral , 
            n29777, n29776, n29775, n29774, n29773, n29772, n29771, 
            n29770, n29769, n29768, n29767, n29766, n29765, n29764, 
            n29763, n29762, n29761, n29760, n29759, n29758, n29757, 
            n29754, n28910, \motor_state[23] , \motor_state[22] , \motor_state[21] , 
            \motor_state[20] , \motor_state[19] , \motor_state[18] , \motor_state[17] , 
            \motor_state[16] , \motor_state[15] , n9, \motor_state[13] , 
            \motor_state[12] , \motor_state[11] , n38659, n24981, n38328, 
            n21, n25, n36, n33833, n40, n33791) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input \Ki[2] ;
    output [23:0]n335;
    input [23:0]setpoint;
    input [23:0]deadband;
    input \Ki[3] ;
    input \Kp[7] ;
    input [23:0]IntegralLimit;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Kp[2] ;
    input \Kp[3] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input \Kp[6] ;
    input \Kp[8] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Kp[13] ;
    input \Kp[14] ;
    input \Ki[6] ;
    input \Kp[15] ;
    input \encoder1_position_scaled[0] ;
    input n15;
    input n62934;
    input n15_adj_1;
    input \encoder1_position_scaled[1] ;
    input n62948;
    input \motor_state[9] ;
    output control_update;
    output [23:0]duty;
    input clk16MHz;
    input reset;
    input \motor_state[8] ;
    input \Ki[1] ;
    input \Ki[0] ;
    input [23:0]PWMLimit;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Ki[9] ;
    input \motor_state[7] ;
    input VCC_net;
    input \motor_state[6] ;
    input \Ki[10] ;
    input \Ki[11] ;
    input \Ki[12] ;
    input \Ki[13] ;
    input \motor_state[5] ;
    input \Ki[14] ;
    input \Ki[15] ;
    input \motor_state[4] ;
    input \motor_state[10] ;
    input \motor_state[3] ;
    input n3;
    input [7:0]control_mode;
    output n55181;
    output n105;
    input n7064;
    input n38638;
    input n29778;
    output [23:0]\PID_CONTROLLER.integral ;
    input n29777;
    input n29776;
    input n29775;
    input n29774;
    input n29773;
    input n29772;
    input n29771;
    input n29770;
    input n29769;
    input n29768;
    input n29767;
    input n29766;
    input n29765;
    input n29764;
    input n29763;
    input n29762;
    input n29761;
    input n29760;
    input n29759;
    input n29758;
    input n29757;
    input n29754;
    input n28910;
    input \motor_state[23] ;
    input \motor_state[22] ;
    input \motor_state[21] ;
    input \motor_state[20] ;
    input \motor_state[19] ;
    input \motor_state[18] ;
    input \motor_state[17] ;
    input \motor_state[16] ;
    input \motor_state[15] ;
    input n9;
    input \motor_state[13] ;
    input \motor_state[12] ;
    input \motor_state[11] ;
    output n38659;
    input n24981;
    output n38328;
    input n21;
    input n25;
    output n36;
    input n33833;
    output n40;
    input n33791;
    
    wire clk16MHz /* synthesis SET_AS_NETWORK=clk16MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(41[6:14])
    
    wire n6;
    wire [23:0]n455;
    
    wire n21_c, n65191, n159, n9972, n63174, n4744, n67071;
    wire [23:0]n535;
    
    wire n67074, n43;
    wire [13:0]n18600;
    wire [12:0]n18990;
    
    wire n977, n49311, n23, n65192, n49312, n904, n49310;
    wire [12:0]n18825;
    wire [11:0]n19186;
    
    wire n542, n48668, n48669, n63173, n67065, n67068, n37, n63172, 
        n67059, n67062, n469_adj_4430, n48667, n831, n49309, n758, 
        n49308, n685, n49307, n396, n48666, n612, n49306, n539, 
        n49305, n466, n49304, n17, n8, n393, n49303, n323, n48665, 
        n320, n49302, n247, n49301, n174, n49300, n35, n250, 
        n48664, n63168, n67053, n232;
    wire [23:0]n207;
    
    wire n524, n67056, n32, n101;
    wire [11:0]n19326;
    
    wire n980, n49299, n907, n49298, n29, n177, n48663, n16, 
        n45, n24, n43_adj_4431, n25_c, n63616, n63552, n63167, 
        n67047, n834, n49297, n67050, n761, n49296, n688, n49295, 
        n35_adj_4432, n104, n615, n49294, n262, n150;
    wire [23:0]n233;
    
    wire n41, n33, n223_adj_4433, n77, n31, n8_adj_4434, n335_c, 
        n39, n296, n63160, n67041, n369, n150_adj_4435, n223_adj_4436, 
        n296_adj_4437, n67044, n45_adj_4438, n369_adj_4439, n442, 
        n515, n588, n661, n734, n807, n880, n953, n1026, n43_adj_4440, 
        n29_adj_4441, n31_adj_4442, n597, n408, n442_adj_4443, n1099;
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(290[22:33])
    
    wire n23_adj_4445, n25_adj_4446, n37_adj_4447, n35_adj_4448, n33_adj_4449, 
        n48292, n542_adj_4450, n49293, n469_adj_4451, n49292, n48293, 
        n67014, counter_31__N_3714, n63549, n65480, n48291;
    wire [23:0]n28;
    
    wire n63709, n396_adj_4452, n49291, n323_adj_4453, n49290, n250_adj_4454, 
        n49289, n177_adj_4455, n49288, n35_adj_4456, n104_adj_4457, 
        n9_c;
    wire [23:0]n285;
    
    wire n284;
    wire [23:0]n310;
    
    wire n258, n64678, n17_adj_4458, n74, n63142, n67029, n5, 
        n147, n220, n64372, n481, n19, n4, n21_adj_4460, n554_adj_4461, 
        n515_adj_4462, n11, n627, n700, n13, n588_adj_4463, n74_adj_4464, 
        n5_adj_4465, n27, n65189, n29_adj_4467, n65190, n110, n41_adj_4469, 
        n67220, n15_adj_4471, n33_adj_4472, n31_adj_4473, n63596, 
        n63586, n67032, n293, n27_adj_4474;
    wire [10:0]n19495;
    
    wire n910, n48653, n837, n48652, n147_adj_4475, n220_adj_4476, 
        n293_adj_4477, n764, n48651, n64658, n691, n48650, n64027, 
        n64016, n670, n305, n67215, n378;
    wire [0:0]n10361;
    wire [21:0]n10958;
    
    wire n48917;
    wire [47:0]n34;
    
    wire n48916, n183, n618, n48649, n366, n743, n366_adj_4478, 
        n451, n524_adj_4479, n256_adj_4480, n545, n48648;
    wire [13:0]n61;
    wire [31:0]counter;   // verilog/motorControl.v(22[11:18])
    
    wire n49223, n48915, n48914, n472_adj_4481, n48647, n399, n48646, 
        n12, n49222, n49221, n329, n49220, n48913, n49219, n816, 
        n48290, n326, n48645, n597_adj_4482, n49218, n49217, n49216, 
        n49215, n253_adj_4483, n48644, n49214, n48912, n49213, n49212, 
        n439, n49211, n48911, n180, n48643, n48910, n38, n107;
    wire [6:0]n20336;
    wire [5:0]n20432;
    
    wire n560, n48642, n1096, n48909, n487, n48641, n414, n48640, 
        n1023, n48908, n341, n48639, n950, n48907, n268, n48638, 
        n877, n48906, n195, n48637, n889, n30, n10, n35_adj_4486, 
        n63577, n65869, n64374, n53, n122, n66090, n37_adj_4487, 
        n66091, n804, n48905;
    wire [9:0]n19756;
    
    wire n840, n48636, n10_adj_4489, n30_adj_4490, n670_adj_4491, 
        n731, n48904, n767, n48635, n402, n694, n48634, n64043, 
        n64963, n64955, n658, n48903, n621, n48633, n63697, n65947, 
        n48289, n585, n48902, n548, n48632, n65385, n743_adj_4492, 
        n66086, n962, n512, n816_adj_4493, n475_adj_4494, n64670, 
        n16_adj_4495, n889_adj_4496, n48631, n962_adj_4497, n1035, 
        n48901, n6_adj_4498, n65651, n65652, n48630, n48288, n1035_adj_4499, 
        n1108, n8_adj_4500, n48900, n48629, n67235, n48628, n48899, 
        n24_adj_4501, n48627, n48287, n63941, n1108_adj_4502, n63935, 
        n65472, n39_adj_4503, n66065, n64332, n4_adj_4504, n48898, 
        n65647, n65648, n119, n64000, n50, n63990, n65965, n64334, 
        n64666, n67230, n48897, n66176, n63118, n66741, n48896, 
        n66177, n192, n41_adj_4507, n66060, n63555, n265, n66149, 
        n48294, n48286, n48285, n48284, n338, n16_adj_4508, n411, 
        n63140, n67017, n67020, n63646, n484_adj_4509, n63139, n67011, 
        n439_adj_4510, n63954, n65807, n8_adj_4511, n24_adj_4512, 
        n63716, n67228, n63713, n67256, n66021, n64340, n66023, 
        n41_adj_4513, n39_adj_4514, n45_adj_4515, n43_adj_4516, n66744, 
        n37_adj_4517, n29_adj_4518, n31_adj_4519, n23_adj_4520, n25_adj_4521, 
        n35_adj_4522, n33_adj_4523, n11_adj_4524, n13_adj_4525, n15_adj_4526, 
        n27_adj_4527, n9_adj_4529, n17_adj_4530, n19_adj_4531, n21_adj_4532, 
        n65247, n63900, n63886, n12_adj_4533, n10_adj_4534, n30_adj_4535, 
        n63931, n64863, n64855, n557_adj_4536, n65931, n64380, n66037, 
        n45_adj_4537, n37_adj_4538, n41_adj_4540, n43_adj_4541;
    wire [8:0]n19973;
    
    wire n770, n48611, n29_adj_4543, n67253, n31_adj_4544, n33_adj_4545, 
        n697, n48610, n39_adj_4546, n35_adj_4548, n65319, n6_adj_4549, 
        n66080, n64674, n630, n16_adj_4550, n624, n48609, n25015, 
        n21_adj_4551, n19_adj_4552, n17_adj_4553, n9_adj_4554, n64127, 
        n6_adj_4555, n65643, n27_adj_4556, n15_adj_4557, n13_adj_4558, 
        n11_adj_4559, n64108, n12_adj_4560, n10_adj_4561, n30_adj_4562, 
        n65644;
    wire [20:0]n12488;
    
    wire n48883, n83, n48882, n64177, n65043, n65027, n8_adj_4563, 
        n25_adj_4564, n23_adj_4565, n65957, n24_adj_4566;
    wire [10:0]n19612;
    
    wire n910_adj_4567, n49108, n551_adj_4568, n48608, n837_adj_4569, 
        n49107, n48881, n478_adj_4570, n48607, n764_adj_4571, n49106, 
        n691_adj_4572, n49105, n65413, n618_adj_4573, n49104, n545_adj_4574, 
        n49103, n472_adj_4575, n49102, n399_adj_4576, n49101, n66088, 
        n16_adj_4577, n14, n512_adj_4578, n65673, n83_adj_4579, n14_adj_4580, 
        n326_adj_4581, n49100, n405, n48606, n332, n48605, n48880, 
        n253_adj_4582, n49099, n180_adj_4583, n49098, n259, n48604, 
        n38_adj_4584, n107_adj_4585, n6_adj_4586, n65659, n48879, 
        n63822, n186, n48603, n48878, n44, n113, n63818, n65474, 
        n64342, n156, n229, n63687, n67218, n65233, n67247, n48877, 
        n4_adj_4587, n1099_adj_4588, n48876, n65889, n65660, n67209, 
        n65641, n66154, n1026_adj_4591, n48875, n156_adj_4592, n953_adj_4593, 
        n48874, n65642, n880_adj_4594, n48873, n57914, n490_adj_4595, 
        n48596, n63876, n63872, n65967, n302_adj_4596;
    wire [4:0]n20502;
    
    wire n417, n48595, n67206, n63117, n66735, n8_adj_4597, n27_adj_4598, 
        n15_adj_4599, n13_adj_4600, n11_adj_4601, n63783, n229_adj_4602, 
        n807_adj_4603, n48872, n64344, n585_adj_4604, n344_adj_4605, 
        n48594, n375, n66178, n271, n48593, n66179, n658_adj_4606, 
        n731_adj_4607, n734_adj_4608, n48871, n198, n48592, n661_adj_4609, 
        n48870, n66738, n66147, n63826, n12_adj_4610, n448_adj_4611, 
        n24_adj_4612, n63116, n66729, n66732, n63115, n66723, n66726, 
        n10_adj_4613;
    wire [0:0]n11041;
    wire [21:0]n11500;
    
    wire n49492;
    wire [43:0]n360;
    
    wire n49491, n30_adj_4614, n49490, n49489, n49488, n49487, n49486, 
        n64052, n49485, n302_adj_4615, n1096_adj_4616, n49484, n1023_adj_4617, 
        n49483, n950_adj_4618, n49482, n877_adj_4619, n49481, n66025, 
        n56, n125, n804_adj_4621, n49480, n49479, n49478, n49477, 
        n49476, n64350, n49475, n9_adj_4623, n63814, n64770, n19_adj_4624, 
        n17_adj_4625, n64764, n63114, n66705, n66708, n25_adj_4626, 
        n23_adj_4627, n21_adj_4628, n65913, n65277, n49474, n49473, 
        n64046, n65470, n49472, n49471, n48869, n66027, n63546;
    wire [7:0]n20150;
    
    wire n48591, n48590, n66074;
    wire [20:0]n12999;
    
    wire n49470, n49469, n48868, n64322, n4_adj_4631, n65657, n65658, 
        n64089, n48589, n64076, n65963, n6_adj_4632, n49468, n64324, 
        n66174, n66175, n66153, n64056, n66017, n49467, n64330, 
        n66019, n37_adj_4633, n45_adj_4634, n41_adj_4635, n49466, 
        n43_adj_4636, n35_adj_4637, n16_adj_4638, n49465, n48588, 
        n63644, n63111, n66687, n49464, n39_adj_4639, n31_adj_4640, 
        n521, n33_adj_4641, n27_adj_4642, n29_adj_4643, n7062, n24983, 
        n49463, n48867, n594, n48587, n49462, n49461, n49460, 
        n6_adj_4644, n49459, n49458, n49457, n49456, n49455, n49454, 
        n49453, n49452, n375_adj_4645, n49451, n667, n49450, n48866, 
        n48865, n48586, n448_adj_4646, n48864, n48863, n48585;
    wire [19:0]n14310;
    
    wire n49449, n8_adj_4647, n77_adj_4648, n49448, n189, n48584;
    wire [19:0]n13844;
    
    wire n48862, n49447, n47, n116, n15_adj_4649, n13_adj_4650, 
        n11_adj_4651, n63510, n8_adj_4652, n12_adj_4653, n49446, n48861, 
        n48860, n48859, n49445, n48858, n49444, n48857, n45_adj_4654, 
        n24_adj_4655, n66690, n1102, n48856, n1102_adj_4656, n49443, 
        n10_adj_4657, n30_adj_4658, n9_adj_4659, n64548, n19_adj_4660, 
        n17_adj_4661, n64542, n25_adj_4662, n23_adj_4663, n21_adj_4664, 
        n65847, n65149, n66047, n65179, n65180, n16_adj_4665, n1029, 
        n48855, n1029_adj_4666, n49442, n956, n48854, n66852, n883, 
        n48853, n956_adj_4667, n49441, n810, n48852, n883_adj_4668, 
        n49440, n737, n48851, n664, n48850, n810_adj_4669, n49439, 
        n591, n48849, n737_adj_4670, n49438, n664_adj_4671, n49437, 
        n65637, n518, n48848, n445_adj_4672, n48847, n372, n48846, 
        n591_adj_4673, n49436, n518_adj_4674, n49435, n445_adj_4675, 
        n49434, n299_adj_4676, n48845, n226_adj_4677, n48844, n372_adj_4678, 
        n49433, n299_adj_4679, n49432, n226_adj_4680, n49431, n153, 
        n48843, n153_adj_4681, n49430, n11_adj_4682, n80, n11_adj_4683, 
        n80_adj_4684;
    wire [9:0]n19852;
    wire [8:0]n20050;
    
    wire n770_adj_4685, n48842, n697_adj_4686, n48841;
    wire [18:0]n15476;
    
    wire n49429, n624_adj_4687, n48840, n49428, n551_adj_4688, n48839, 
        n49427, n478_adj_4689, n48838, n49426, n405_adj_4690, n48837, 
        n332_adj_4691, n48836, n63055, n66681, n66684, n49425, n259_adj_4692, 
        n48835, n186_adj_4693, n48834, n44_adj_4694, n113_adj_4695, 
        n1105, n49424;
    wire [18:0]n15053;
    
    wire n48833, n48832, n1032, n49423, n48831, n959, n49422, 
        n48830, n886, n49421, n48829, n1105_adj_4696, n48828, n813, 
        n49420, n740, n49419, n1032_adj_4697, n48827, n667_adj_4698, 
        n49418, n959_adj_4699, n48826, n886_adj_4700, n48825, n813_adj_4701, 
        n48824, n594_adj_4702, n49417, n521_adj_4703, n49416, n740_adj_4704, 
        n48823, n49415, n48822, n49414, n48821, n48820, n49413, 
        n48819, n48818, n49412, n48817, n49411, n66666, n66660, 
        n66570, n67098, n67092, n67086, n67080, n48816, n48815;
    wire [6:0]n20291;
    
    wire n49410, n49409, n65638, n49408, n49407, n63793, n49406, 
        n48352, n49405, n48351, n48350, n63724, n63718, n65476, 
        n64352, n62983, n4_adj_4705, n65629, n49404, n48349, n48348, 
        n48347;
    wire [17:0]n16401;
    
    wire n49403, n48346, n49402, n48345, n48344;
    wire [17:0]n16054;
    
    wire n48802, n48801, n49401, n49400, n48800, n48799, n48343, 
        n49399, n48342, n48798, n48797, n49398, n48796, n65630, 
        n48341, n48795, n48794, n49397, n48340, n48793, n48339, 
        n8_adj_4706, n24_adj_4707, n48792, n48338, n49396, n48337, 
        n48791, n49395, n48790, n48789, n48336, n63521, n63474, 
        n63464, n65482, n64382, n48335, n49394, n48788, n48015, 
        n59388, n48787, n48334, n49393, n48333, n49392, n39_adj_4708, 
        n49391, n48786, n63178, n67095, n48785, n48332, n12_adj_4709, 
        n48331, n17_adj_4710, n86;
    wire [23:0]n1_adj_4992;
    
    wire n48498, n48330, n451_adj_4711, n49390, n48497, n48496, 
        n48329, n48328, n378_adj_4714, n49389, n48495, n48327, n305_adj_4716, 
        n49388, n48494, n48493, n232_adj_4718, n49387, n48326, n159_adj_4719, 
        n49386, n48492, n17_adj_4721, n86_adj_4722;
    wire [16:0]n17048;
    
    wire n49385, n48491;
    wire [3:0]n20550;
    
    wire n4_adj_4724, n49384, n63669, n49383, n1111, n49382;
    wire [16:0]n16763;
    
    wire n48773, n48772, n1038, n49381, n48771, n1111_adj_4725, 
        n48770, n67241, n1038_adj_4726, n48769, n965, n49380, n965_adj_4727, 
        n48768, n892, n48767, n48490, n892_adj_4729, n49379, n819, 
        n48766, n746, n48765, n48489, n819_adj_4731, n49378, n673, 
        n48764, n48488, n746_adj_4733, n49377, n600, n48763, n673_adj_4734, 
        n49376, n600_adj_4735, n49375, n63177, n67089, n527, n48762, 
        n527_adj_4736, n49374, n48487, n454, n49373, n454_adj_4738, 
        n48761, n381, n48760, n381_adj_4739, n49372, n308_adj_4740, 
        n48759, n308_adj_4741, n49371, n235_adj_4742, n48758, n162, 
        n48757, n20, n89, n235_adj_4743, n49370;
    wire [15:0]n17373;
    
    wire n48756, n48755, n48486, n162_adj_4745, n49369, n1114, n48754, 
        n1041, n48753, n20_adj_4746, n89_adj_4747, n968, n48752;
    wire [15:0]n17625;
    
    wire n49368, n895, n48751, n49367, n822, n48750, n749, n48749, 
        n1114_adj_4748, n49366, n676, n48748, n603, n48747, n530, 
        n48746, n1041_adj_4749, n49365, n457_adj_4750, n48745, n384_adj_4751, 
        n48744, n968_adj_4752, n49364, n311_adj_4753, n48743, n10_adj_4754, 
        n238_adj_4755, n48742, n895_adj_4756, n49363, n165, n48741, 
        n23_adj_4757, n92, n48485, n822_adj_4759, n49362;
    wire [14:0]n17931;
    
    wire n48740, n1117, n48739, n749_adj_4760, n49361, n48484, n1044, 
        n48738, n676_adj_4762, n49360, n971, n48737, n898, n48736, 
        n825, n48735, n603_adj_4763, n49359, n752, n48734, n48483, 
        n63176, n67083, n840_adj_4765, n48972, n48325, n530_adj_4766, 
        n49358, n48482, n48324, n679, n48733, n48481, n457_adj_4768, 
        n49357, n48480, n606, n48732, n48479, n48478, n48323, 
        n533, n48731, n48477, n48322, n384_adj_4772, n49356, n767_adj_4773, 
        n48971, n311_adj_4774, n49355, n460_adj_4775, n48730, n30_adj_4776, 
        n48476, n387_adj_4778, n48729, n47_adj_4780;
    wire [23:0]n1_adj_4993;
    
    wire n48475, n238_adj_4782, n49354, n314, n48728, n48474, n694_adj_4784, 
        n48970, n241_adj_4785, n48727, n48473, n168, n48726, n48472, 
        n165_adj_4788, n49353, n48471, n26, n95, n48470, n48469;
    wire [7:0]n20210;
    
    wire n700_adj_4792, n48725, n48468, n48321, n23_adj_4794, n92_adj_4795, 
        n627_adj_4796, n48724, n48467, n48466, n63677, n554_adj_4799, 
        n48723, n48465, n48320, n48464, n48319;
    wire [5:0]n20400;
    
    wire n560_adj_4802, n49352, n481_adj_4803, n48722, n48463, n48318, 
        n48462, n48317, n487_adj_4806, n49351, n408_adj_4807, n48721, 
        n48461, n48316, n414_adj_4809, n49350, n48460, n48459, n48315, 
        n621_adj_4812, n48969, n341_adj_4813, n49349, n335_adj_4814, 
        n48720, n48458, n262_adj_4816, n48719, n48457, n268_adj_4818, 
        n49348, n548_adj_4819, n48968, n475_adj_4820, n48967, n48314, 
        n189_adj_4821, n48718, n48456, n48313, n48455, n48312, n195_adj_4825, 
        n49347, n47_adj_4826, n116_adj_4827, n48454, n402_adj_4829, 
        n48966, n329_adj_4830, n48965, n53_adj_4831, n122_adj_4832, 
        n256_adj_4833, n48964, n48453, n48311;
    wire [14:0]n18152;
    
    wire n49346, n1117_adj_4835, n49345, n48310, n38672;
    wire [23:0]n1_adj_4994;
    
    wire n48452, n48451, n183_adj_4839, n48963, n1044_adj_4840, n49344, 
        n41_adj_4841, n110_adj_4842, n48309, n971_adj_4843, n49343, 
        n48450, n48308, n48449, n898_adj_4846, n49342, n48448, n347_adj_4848, 
        n48447, n48446, n48445, n825_adj_4852, n49341, n48444, n6_adj_4854, 
        n55858, n752_adj_4855, n49340, n48443, n48442, n48441, n48307, 
        n679_adj_4859, n49339;
    wire [13:0]n18408;
    
    wire n1120, n48708, n48440, n1047, n48707, n48439, n974, n48706, 
        n48438, n901, n48705, n606_adj_4863, n49338, n828, n48704, 
        n48437, n48436, n533_adj_4866, n49337, n755, n48703, n48435, 
        n48434, n460_adj_4869, n49336, n682, n48702, n48433, n48432, 
        n609, n48701, n48431, n387_adj_4873, n49335, n536_adj_4874, 
        n48700, n48430, n59384, n463_adj_4877, n48699, n314_adj_4878, 
        n49334, n48306, n48305, n48304, n390_adj_4879, n48698, n48303, 
        n317, n48697, n48302, n241_adj_4880, n49333, n168_adj_4881, 
        n49332, n244_adj_4882, n48696, n26_adj_4883, n95_adj_4884, 
        n171, n48695, n29_adj_4885, n98, n48301, n48300, n1120_adj_4886, 
        n49331, n1047_adj_4887, n49330, n48299, n974_adj_4888, n49329, 
        n1050, n48694, n977_adj_4889, n48693, n48298, n901_adj_4890, 
        n49328, n904_adj_4891, n48692, n48297, n48296, n831_adj_4893, 
        n48691, n828_adj_4894, n49327, n755_adj_4895, n49326, n758_adj_4896, 
        n48690, n48295, n685_adj_4897, n48689, n682_adj_4898, n49325, 
        n609_adj_4899, n49324, n612_adj_4900, n48688, n536_adj_4901, 
        n49323, n463_adj_4902, n49322, n68_adj_4903, n63175, n67077, 
        n539_adj_4904, n48687, n390_adj_4905, n49321, n466_adj_4906, 
        n48686, n393_adj_4907, n48685, n320_adj_4908, n48684, n317_adj_4909, 
        n49320, n247_adj_4910, n48683, n244_adj_4911, n49319, n174_adj_4912, 
        n48682, n32_adj_4913, n101_adj_4914, n171_adj_4915, n49318, 
        n630_adj_4916, n48681, n557_adj_4917, n48680, n29_adj_4918, 
        n98_adj_4919, n484_adj_4920, n48679, n411_adj_4921, n48678, 
        n57863, n490_adj_4922, n49317;
    wire [4:0]n20481;
    
    wire n417_adj_4923, n49316, n338_adj_4924, n48677, n344_adj_4925, 
        n49315, n265_adj_4926, n48676, n192_adj_4927, n48675, n50_adj_4928, 
        n119_adj_4929, n271_adj_4930, n49314, n198_adj_4931, n49313, 
        n980_adj_4932, n48674, n907_adj_4933, n48673, n834_adj_4934, 
        n48672, n56_adj_4935, n125_adj_4936, n761_adj_4937, n48671, 
        n688_adj_4938, n48670, n1050_adj_4939, n615_adj_4940, n48010, 
        n49517, n59374, n67502, n59378, n65971, n8_adj_4941, n6_adj_4942, 
        n9_adj_4943, n11_adj_4944, n13_adj_4945, n15_adj_4946, n19_adj_4947, 
        n64364;
    wire [3:0]n20538;
    
    wire n6_adj_4949, n66182, n4_adj_4951, n65177, n66183, n65178;
    wire [1:0]n20596;
    
    wire n47985;
    wire [2:0]n20575;
    
    wire n66143, n59342, n59346, n59344, n63492, n47955, n59352, 
        n4_adj_4953, n8_adj_4954, n6_adj_4955, n6_adj_4956, n6_adj_4957, 
        n63239, n8_adj_4958, n10_adj_4959, n65631, n63488, n65865, 
        n63259, n65632, n64384, n63649, n66092, n66093, n67204, 
        n65478, n64362, n66063, n63476, n63651, n63132, n66849, 
        n65809, n66033, n64390, n64370, n66035, n4_adj_4965, n65635, 
        n66039, n65636, n4_adj_4966, n57934, n63761, n63757, n65969, 
        n25017, n64354, n66180, n66181, n62945, n66145, n63019, 
        n41_adj_4967, n63737, n63054, n66029, n66663, n64360, n66036, 
        n66031, n66657, n58117, n18_adj_4968, n20_adj_4969, n7_adj_4970, 
        n4_adj_4972, n48038, n4_adj_4973, n48119, n10_adj_4974, n31_adj_4975, 
        n29_adj_4976, n27_adj_4977, n19_adj_4978, n23_adj_4979, n15_adj_4980, 
        n17_adj_4981, n7_adj_4982, n9_adj_4983, n11_adj_4984, n13_adj_4985, 
        n5_adj_4986, n63268, n63253, n65441, n4_adj_4988, n65490, 
        n65491, n64202, n65103, n65464, n16_adj_4989, n66099, n66100, 
        n66008, n66567, n64204, n65488, n65806, n66041, n66042, 
        n65486, n65487, n12_adj_4991, n64616, n64608, n65871, n65181;
    
    SB_LUT4 i48129_3_lut (.I0(n6), .I1(n455[10]), .I2(n21_c), .I3(GND_net), 
            .O(n65191));   // verilog/motorControl.v(63[16:31])
    defparam i48129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i108_2_lut (.I0(\Ki[2] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9972_bdd_4_lut_49919 (.I0(n9972), .I1(n63174), .I2(setpoint[8]), 
            .I3(n4744), .O(n67071));
    defparam n9972_bdd_4_lut_49919.LUT_INIT = 16'he4aa;
    SB_LUT4 n67071_bdd_4_lut (.I0(n67071), .I1(n535[8]), .I2(n455[8]), 
            .I3(n4744), .O(n67074));
    defparam n67071_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_26_i43_2_lut (.I0(deadband[21]), .I1(n455[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4930_14_lut (.I0(GND_net), .I1(n18990[11]), .I2(n977), 
            .I3(n49311), .O(n18600[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4930_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48130_3_lut (.I0(n65191), .I1(n455[11]), .I2(n23), .I3(GND_net), 
            .O(n65192));   // verilog/motorControl.v(63[16:31])
    defparam i48130_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4930_14 (.CI(n49311), .I0(n18990[11]), .I1(n977), .CO(n49312));
    SB_LUT4 add_4930_13_lut (.I0(GND_net), .I1(n18990[10]), .I2(n904), 
            .I3(n49310), .O(n18600[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4930_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4945_8_lut (.I0(GND_net), .I1(n19186[5]), .I2(n542), .I3(n48668), 
            .O(n18825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4945_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4930_13 (.CI(n49310), .I0(n18990[10]), .I1(n904), .CO(n49311));
    SB_CARRY add_4945_8 (.CI(n48668), .I0(n19186[5]), .I1(n542), .CO(n48669));
    SB_LUT4 n9972_bdd_4_lut_49914 (.I0(n9972), .I1(n63173), .I2(setpoint[7]), 
            .I3(n4744), .O(n67065));
    defparam n9972_bdd_4_lut_49914.LUT_INIT = 16'he4aa;
    SB_LUT4 n67065_bdd_4_lut (.I0(n67065), .I1(n535[7]), .I2(n455[7]), 
            .I3(n4744), .O(n67068));
    defparam n67065_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_26_i37_2_lut (.I0(deadband[18]), .I1(n455[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n9972_bdd_4_lut_49909 (.I0(n9972), .I1(n63172), .I2(setpoint[6]), 
            .I3(n4744), .O(n67059));
    defparam n9972_bdd_4_lut_49909.LUT_INIT = 16'he4aa;
    SB_LUT4 n67059_bdd_4_lut (.I0(n67059), .I1(n535[6]), .I2(n455[6]), 
            .I3(n4744), .O(n67062));
    defparam n67059_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_4945_7_lut (.I0(GND_net), .I1(n19186[4]), .I2(n469_adj_4430), 
            .I3(n48667), .O(n18825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4945_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4930_12_lut (.I0(GND_net), .I1(n18990[9]), .I2(n831), 
            .I3(n49309), .O(n18600[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4930_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4930_12 (.CI(n49309), .I0(n18990[9]), .I1(n831), .CO(n49310));
    SB_CARRY add_4945_7 (.CI(n48667), .I0(n19186[4]), .I1(n469_adj_4430), 
            .CO(n48668));
    SB_LUT4 add_4930_11_lut (.I0(GND_net), .I1(n18990[8]), .I2(n758), 
            .I3(n49308), .O(n18600[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4930_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4930_11 (.CI(n49308), .I0(n18990[8]), .I1(n758), .CO(n49309));
    SB_LUT4 add_4930_10_lut (.I0(GND_net), .I1(n18990[7]), .I2(n685), 
            .I3(n49307), .O(n18600[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4930_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4930_10 (.CI(n49307), .I0(n18990[7]), .I1(n685), .CO(n49308));
    SB_LUT4 add_4945_6_lut (.I0(GND_net), .I1(n19186[3]), .I2(n396), .I3(n48666), 
            .O(n18825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4945_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4930_9_lut (.I0(GND_net), .I1(n18990[6]), .I2(n612), .I3(n49306), 
            .O(n18600[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4930_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4930_9 (.CI(n49306), .I0(n18990[6]), .I1(n612), .CO(n49307));
    SB_LUT4 add_4930_8_lut (.I0(GND_net), .I1(n18990[5]), .I2(n539), .I3(n49305), 
            .O(n18600[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4930_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4945_6 (.CI(n48666), .I0(n19186[3]), .I1(n396), .CO(n48667));
    SB_CARRY add_4930_8 (.CI(n49305), .I0(n18990[5]), .I1(n539), .CO(n49306));
    SB_LUT4 add_4930_7_lut (.I0(GND_net), .I1(n18990[4]), .I2(n466), .I3(n49304), 
            .O(n18600[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4930_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_30_i8_3_lut (.I0(n455[4]), .I1(n455[8]), .I2(n17), 
            .I3(GND_net), .O(n8));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4930_7 (.CI(n49304), .I0(n18990[4]), .I1(n466), .CO(n49305));
    SB_LUT4 add_4930_6_lut (.I0(GND_net), .I1(n18990[3]), .I2(n393), .I3(n49303), 
            .O(n18600[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4930_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4945_5_lut (.I0(GND_net), .I1(n19186[2]), .I2(n323), .I3(n48665), 
            .O(n18825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4945_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4930_6 (.CI(n49303), .I0(n18990[3]), .I1(n393), .CO(n49304));
    SB_CARRY add_4945_5 (.CI(n48665), .I0(n19186[2]), .I1(n323), .CO(n48666));
    SB_LUT4 add_4930_5_lut (.I0(GND_net), .I1(n18990[2]), .I2(n320), .I3(n49302), 
            .O(n18600[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4930_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4930_5 (.CI(n49302), .I0(n18990[2]), .I1(n320), .CO(n49303));
    SB_LUT4 add_4930_4_lut (.I0(GND_net), .I1(n18990[1]), .I2(n247), .I3(n49301), 
            .O(n18600[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4930_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4930_4 (.CI(n49301), .I0(n18990[1]), .I1(n247), .CO(n49302));
    SB_LUT4 add_4930_3_lut (.I0(GND_net), .I1(n18990[0]), .I2(n174), .I3(n49300), 
            .O(n18600[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4930_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_26_i35_2_lut (.I0(deadband[17]), .I1(n455[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4945_4_lut (.I0(GND_net), .I1(n19186[1]), .I2(n250), .I3(n48664), 
            .O(n18825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4945_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9972_bdd_4_lut_49904 (.I0(n9972), .I1(n63168), .I2(setpoint[5]), 
            .I3(n4744), .O(n67053));
    defparam n9972_bdd_4_lut_49904.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_24_i157_2_lut (.I0(\Ki[3] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i157_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4930_3 (.CI(n49300), .I0(n18990[0]), .I1(n174), .CO(n49301));
    SB_LUT4 mult_23_i353_2_lut (.I0(\Kp[7] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n67053_bdd_4_lut (.I0(n67053), .I1(n535[5]), .I2(n455[5]), 
            .I3(n4744), .O(n67056));
    defparam n67053_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_4930_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n18600[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4930_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4930_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n49300));
    SB_CARRY add_4945_4 (.CI(n48664), .I0(n19186[1]), .I1(n250), .CO(n48665));
    SB_LUT4 add_4956_14_lut (.I0(GND_net), .I1(n19326[11]), .I2(n980), 
            .I3(n49299), .O(n18990[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4956_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4956_13_lut (.I0(GND_net), .I1(n19326[10]), .I2(n907), 
            .I3(n49298), .O(n18990[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4956_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_26_i29_2_lut (.I0(deadband[14]), .I1(n455[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4945_3_lut (.I0(GND_net), .I1(n19186[0]), .I2(n177), .I3(n48663), 
            .O(n18825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4945_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4956_13 (.CI(n49298), .I0(n19326[10]), .I1(n907), .CO(n49299));
    SB_LUT4 LessThan_30_i24_3_lut (.I0(n16), .I1(n455[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46490_4_lut (.I0(n43_adj_4431), .I1(n25_c), .I2(n23), .I3(n63616), 
            .O(n63552));
    defparam i46490_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 n9972_bdd_4_lut_49899 (.I0(n9972), .I1(n63167), .I2(setpoint[4]), 
            .I3(n4744), .O(n67047));
    defparam n9972_bdd_4_lut_49899.LUT_INIT = 16'he4aa;
    SB_LUT4 add_4956_12_lut (.I0(GND_net), .I1(n19326[9]), .I2(n834), 
            .I3(n49297), .O(n18990[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4956_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4945_3 (.CI(n48663), .I0(n19186[0]), .I1(n177), .CO(n48664));
    SB_CARRY add_4956_12 (.CI(n49297), .I0(n19326[9]), .I1(n834), .CO(n49298));
    SB_LUT4 n67047_bdd_4_lut (.I0(n67047), .I1(n535[4]), .I2(n455[4]), 
            .I3(n4744), .O(n67050));
    defparam n67047_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_4956_11_lut (.I0(GND_net), .I1(n19326[8]), .I2(n761), 
            .I3(n49296), .O(n18990[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4956_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4956_11 (.CI(n49296), .I0(n19326[8]), .I1(n761), .CO(n49297));
    SB_LUT4 add_4956_10_lut (.I0(GND_net), .I1(n19326[7]), .I2(n688), 
            .I3(n49295), .O(n18990[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4956_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4956_10 (.CI(n49295), .I0(n19326[7]), .I1(n688), .CO(n49296));
    SB_LUT4 add_4945_2_lut (.I0(GND_net), .I1(n35_adj_4432), .I2(n104), 
            .I3(GND_net), .O(n18825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4945_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4956_9_lut (.I0(GND_net), .I1(n19326[6]), .I2(n615), .I3(n49294), 
            .O(n18990[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4956_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4956_9 (.CI(n49294), .I0(n19326[6]), .I1(n615), .CO(n49295));
    SB_LUT4 mult_24_i177_2_lut (.I0(\Ki[3] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i102_2_lut (.I0(\Ki[2] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i41_2_lut (.I0(IntegralLimit[20]), .I1(n233[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i33_2_lut (.I0(deadband[16]), .I1(n455[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i151_2_lut (.I0(\Ki[3] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4433));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i53_2_lut (.I0(\Kp[1] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_26_i31_2_lut (.I0(deadband[15]), .I1(n455[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i6_2_lut (.I0(\Kp[0] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4434));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i226_2_lut (.I0(\Ki[4] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335_c));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i39_2_lut (.I0(IntegralLimit[19]), .I1(n233[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i200_2_lut (.I0(\Ki[4] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9972_bdd_4_lut_49894 (.I0(n9972), .I1(n63160), .I2(setpoint[3]), 
            .I3(n4744), .O(n67041));
    defparam n9972_bdd_4_lut_49894.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_24_i249_2_lut (.I0(\Ki[5] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i102_2_lut (.I0(\Kp[2] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4435));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i151_2_lut (.I0(\Kp[3] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4436));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i200_2_lut (.I0(\Kp[4] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n296_adj_4437));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n67041_bdd_4_lut (.I0(n67041), .I1(n535[3]), .I2(n455[3]), 
            .I3(n4744), .O(n67044));
    defparam n67041_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_17_i45_2_lut (.I0(IntegralLimit[22]), .I1(n233[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4438));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i249_2_lut (.I0(\Kp[5] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n369_adj_4439));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i298_2_lut (.I0(\Kp[6] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n442));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i347_2_lut (.I0(\Kp[7] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i396_2_lut (.I0(\Kp[8] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n588));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i445_2_lut (.I0(\Kp[9] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n661));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i494_2_lut (.I0(\Kp[10] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i543_2_lut (.I0(\Kp[11] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i592_2_lut (.I0(\Kp[12] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i641_2_lut (.I0(\Kp[13] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i690_2_lut (.I0(\Kp[14] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1026));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i43_2_lut (.I0(IntegralLimit[21]), .I1(n233[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4440));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i29_2_lut (.I0(IntegralLimit[14]), .I1(n233[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4441));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i31_2_lut (.I0(IntegralLimit[15]), .I1(n233[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4442));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i402_2_lut (.I0(\Kp[8] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i275_2_lut (.I0(\Ki[5] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i298_2_lut (.I0(\Ki[6] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442_adj_4443));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i298_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4945_2 (.CI(GND_net), .I0(n35_adj_4432), .I1(n104), .CO(n48663));
    SB_LUT4 mult_23_i739_2_lut (.I0(\Kp[15] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1099));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49249_4_lut (.I0(\encoder1_position_scaled[0] ), .I1(n15), 
            .I2(n62934), .I3(n15_adj_1), .O(motor_state[0]));   // verilog/motorControl.v(53[17:33])
    defparam i49249_4_lut.LUT_INIT = 16'h3f77;
    SB_LUT4 LessThan_17_i23_2_lut (.I0(IntegralLimit[11]), .I1(n233[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4445));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i25_2_lut (.I0(IntegralLimit[12]), .I1(n233[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4446));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i37_2_lut (.I0(IntegralLimit[18]), .I1(n233[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4447));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i49272_4_lut (.I0(\encoder1_position_scaled[1] ), .I1(n15), 
            .I2(n62948), .I3(n15_adj_1), .O(motor_state[1]));   // verilog/motorControl.v(53[17:33])
    defparam i49272_4_lut.LUT_INIT = 16'h3f77;
    SB_LUT4 LessThan_17_i35_2_lut (.I0(IntegralLimit[17]), .I1(n233[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4448));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i33_2_lut (.I0(IntegralLimit[16]), .I1(n233[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4449));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_15_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(\motor_state[9] ), 
            .I3(n48292), .O(n207[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4956_8_lut (.I0(GND_net), .I1(n19326[5]), .I2(n542_adj_4450), 
            .I3(n49293), .O(n18990[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4956_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4956_8 (.CI(n49293), .I0(n19326[5]), .I1(n542_adj_4450), 
            .CO(n49294));
    SB_LUT4 add_4956_7_lut (.I0(GND_net), .I1(n19326[4]), .I2(n469_adj_4451), 
            .I3(n49292), .O(n18990[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4956_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_11 (.CI(n48292), .I0(setpoint[9]), .I1(\motor_state[9] ), 
            .CO(n48293));
    SB_DFFER result_i0_i0 (.Q(duty[0]), .C(clk16MHz), .E(control_update), 
            .D(n67014), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFF control_update_46 (.Q(control_update), .C(clk16MHz), .D(counter_31__N_3714));   // verilog/motorControl.v(24[10] 31[6])
    SB_LUT4 i48418_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n63549), 
            .O(n65480));   // verilog/motorControl.v(63[16:31])
    defparam i48418_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 sub_15_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(\motor_state[8] ), 
            .I3(n48291), .O(n207[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46647_4_lut (.I0(n455[6]), .I1(n455[5]), .I2(n28[6]), .I3(n28[5]), 
            .O(n63709));
    defparam i46647_4_lut.LUT_INIT = 16'h7bde;
    SB_CARRY add_4956_7 (.CI(n49292), .I0(n19326[4]), .I1(n469_adj_4451), 
            .CO(n49293));
    SB_LUT4 add_4956_6_lut (.I0(GND_net), .I1(n19326[3]), .I2(n396_adj_4452), 
            .I3(n49291), .O(n18990[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4956_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4956_6 (.CI(n49291), .I0(n19326[3]), .I1(n396_adj_4452), 
            .CO(n49292));
    SB_LUT4 add_4956_5_lut (.I0(GND_net), .I1(n19326[2]), .I2(n323_adj_4453), 
            .I3(n49290), .O(n18990[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4956_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4956_5 (.CI(n49290), .I0(n19326[2]), .I1(n323_adj_4453), 
            .CO(n49291));
    SB_LUT4 add_4956_4_lut (.I0(GND_net), .I1(n19326[1]), .I2(n250_adj_4454), 
            .I3(n49289), .O(n18990[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4956_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4956_4 (.CI(n49289), .I0(n19326[1]), .I1(n250_adj_4454), 
            .CO(n49290));
    SB_LUT4 add_4956_3_lut (.I0(GND_net), .I1(n19326[0]), .I2(n177_adj_4455), 
            .I3(n49288), .O(n18990[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4956_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4956_3 (.CI(n49288), .I0(n19326[0]), .I1(n177_adj_4455), 
            .CO(n49289));
    SB_LUT4 add_4956_2_lut (.I0(GND_net), .I1(n35_adj_4456), .I2(n104_adj_4457), 
            .I3(GND_net), .O(n18990[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4956_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4956_2 (.CI(GND_net), .I0(n35_adj_4456), .I1(n104_adj_4457), 
            .CO(n49288));
    SB_LUT4 LessThan_17_i9_2_lut (.I0(IntegralLimit[4]), .I1(n233[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_c));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_21_i2_3_lut (.I0(n233[1]), .I1(n285[1]), .I2(n284), .I3(GND_net), 
            .O(n310[1]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i2_3_lut (.I0(n310[1]), .I1(IntegralLimit[1]), .I2(n258), 
            .I3(GND_net), .O(n335[1]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47616_3_lut (.I0(n455[7]), .I1(n63709), .I2(n28[7]), .I3(GND_net), 
            .O(n64678));
    defparam i47616_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 LessThan_17_i17_2_lut (.I0(IntegralLimit[8]), .I1(n233[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4458));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i51_2_lut (.I0(\Ki[1] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9972_bdd_4_lut_49889 (.I0(n9972), .I1(n63142), .I2(setpoint[2]), 
            .I3(n4744), .O(n67029));
    defparam n9972_bdd_4_lut_49889.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_24_i4_2_lut (.I0(\Ki[0] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i100_2_lut (.I0(\Ki[2] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i149_2_lut (.I0(\Ki[3] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47310_3_lut (.I0(n65192), .I1(n455[12]), .I2(n25_c), .I3(GND_net), 
            .O(n64372));   // verilog/motorControl.v(63[16:31])
    defparam i47310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i324_2_lut (.I0(\Ki[6] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i19_2_lut (.I0(IntegralLimit[9]), .I1(n233[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i4_4_lut (.I0(n455[0]), .I1(n455[1]), .I2(PWMLimit[1]), 
            .I3(PWMLimit[0]), .O(n4));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 LessThan_17_i21_2_lut (.I0(IntegralLimit[10]), .I1(n233[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4460));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i373_2_lut (.I0(\Ki[7] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4461));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i347_2_lut (.I0(\Ki[7] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515_adj_4462));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i11_2_lut (.I0(IntegralLimit[5]), .I1(n233[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i422_2_lut (.I0(\Ki[8] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i471_2_lut (.I0(\Ki[9] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i13_2_lut (.I0(IntegralLimit[6]), .I1(n233[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i396_2_lut (.I0(\Ki[8] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_4463));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i51_2_lut (.I0(\Kp[1] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4464));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i4_2_lut (.I0(\Kp[0] ), .I1(n207[5]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4465));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48127_3_lut (.I0(n4), .I1(n455[13]), .I2(n27), .I3(GND_net), 
            .O(n65189));   // verilog/motorControl.v(63[16:31])
    defparam i48127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48128_3_lut (.I0(n65189), .I1(n455[14]), .I2(n29_adj_4467), 
            .I3(GND_net), .O(n65190));   // verilog/motorControl.v(63[16:31])
    defparam i48128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i14_3_lut (.I0(n233[13]), .I1(n285[13]), .I2(n284), 
            .I3(GND_net), .O(n310[13]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i14_3_lut (.I0(n310[13]), .I1(IntegralLimit[13]), .I2(n258), 
            .I3(GND_net), .O(n335[13]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i75_2_lut (.I0(\Ki[1] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i28_2_lut (.I0(\Ki[0] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4469));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_28_i27_rep_74_2_lut (.I0(n455[13]), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n67220));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i27_rep_74_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_17_i15_2_lut (.I0(IntegralLimit[7]), .I1(n233[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4471));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46524_4_lut (.I0(n33_adj_4472), .I1(n31_adj_4473), .I2(n29_adj_4467), 
            .I3(n63596), .O(n63586));
    defparam i46524_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 n67029_bdd_4_lut (.I0(n67029), .I1(n535[2]), .I2(n455[2]), 
            .I3(n4744), .O(n67032));
    defparam n67029_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mult_24_i198_2_lut (.I0(\Ki[4] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i27_2_lut (.I0(IntegralLimit[13]), .I1(n233[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4474));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4970_13_lut (.I0(GND_net), .I1(n19495[10]), .I2(n910), 
            .I3(n48653), .O(n19186[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4970_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4970_12_lut (.I0(GND_net), .I1(n19495[9]), .I2(n837), 
            .I3(n48652), .O(n19186[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4970_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i100_2_lut (.I0(\Kp[2] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4475));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i149_2_lut (.I0(\Kp[3] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n220_adj_4476));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i198_2_lut (.I0(\Kp[4] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n293_adj_4477));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i198_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4970_12 (.CI(n48652), .I0(n19495[9]), .I1(n837), .CO(n48653));
    SB_LUT4 add_4970_11_lut (.I0(GND_net), .I1(n19495[8]), .I2(n764), 
            .I3(n48651), .O(n19186[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4970_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_10 (.CI(n48291), .I0(setpoint[8]), .I1(\motor_state[8] ), 
            .CO(n48292));
    SB_LUT4 i47596_4_lut (.I0(n455[14]), .I1(n67220), .I2(n28[14]), .I3(n64678), 
            .O(n64658));
    defparam i47596_4_lut.LUT_INIT = 16'hdeff;
    SB_CARRY add_4970_11 (.CI(n48651), .I0(n19495[8]), .I1(n764), .CO(n48652));
    SB_LUT4 add_4970_10_lut (.I0(GND_net), .I1(n19495[7]), .I2(n691), 
            .I3(n48650), .O(n19186[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4970_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4970_10 (.CI(n48650), .I0(n19495[7]), .I1(n691), .CO(n48651));
    SB_LUT4 i46965_4_lut (.I0(n21_adj_4460), .I1(n19), .I2(n17_adj_4458), 
            .I3(n9_c), .O(n64027));
    defparam i46965_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46954_4_lut (.I0(n27_adj_4474), .I1(n15_adj_4471), .I2(n13), 
            .I3(n11), .O(n64016));
    defparam i46954_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_i451_2_lut (.I0(\Kp[9] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i206_2_lut (.I0(\Ki[4] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_28_i31_rep_69_2_lut (.I0(n455[15]), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n67215));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i31_rep_69_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i255_2_lut (.I0(\Ki[5] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_add_1225_24_lut (.I0(n335[23]), .I1(n10958[21]), .I2(GND_net), 
            .I3(n48917), .O(n10361[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_24_add_1225_23_lut (.I0(GND_net), .I1(n10958[20]), .I2(GND_net), 
            .I3(n48916), .O(n34[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i124_2_lut (.I0(\Ki[2] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4970_9_lut (.I0(GND_net), .I1(n19495[6]), .I2(n618), .I3(n48649), 
            .O(n19186[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4970_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i247_2_lut (.I0(\Kp[5] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n366));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i500_2_lut (.I0(\Kp[10] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i247_2_lut (.I0(\Ki[5] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366_adj_4478));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i247_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_24_add_1225_23 (.CI(n48916), .I0(n10958[20]), .I1(GND_net), 
            .CO(n48917));
    SB_LUT4 mult_24_i304_2_lut (.I0(\Ki[6] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i304_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4970_9 (.CI(n48649), .I0(n19495[6]), .I1(n618), .CO(n48650));
    SB_LUT4 mult_24_i353_2_lut (.I0(\Ki[7] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524_adj_4479));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i173_2_lut (.I0(\Ki[3] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4480));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4970_8_lut (.I0(GND_net), .I1(n19495[5]), .I2(n545), .I3(n48648), 
            .O(n19186[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4970_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2045_2046_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[13]), .I3(n49223), .O(n61[13])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_22_lut (.I0(GND_net), .I1(n10958[19]), .I2(GND_net), 
            .I3(n48915), .O(n34[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_22 (.CI(n48915), .I0(n10958[19]), .I1(GND_net), 
            .CO(n48916));
    SB_CARRY add_4970_8 (.CI(n48648), .I0(n19495[5]), .I1(n545), .CO(n48649));
    SB_LUT4 mult_24_add_1225_21_lut (.I0(GND_net), .I1(n10958[18]), .I2(GND_net), 
            .I3(n48914), .O(n34[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4970_7_lut (.I0(GND_net), .I1(n19495[4]), .I2(n472_adj_4481), 
            .I3(n48647), .O(n19186[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4970_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4970_7 (.CI(n48647), .I0(n19495[4]), .I1(n472_adj_4481), 
            .CO(n48648));
    SB_LUT4 add_4970_6_lut (.I0(GND_net), .I1(n19495[3]), .I2(n399), .I3(n48646), 
            .O(n19186[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4970_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i12_3_lut (.I0(n233[7]), .I1(n233[16]), .I2(n33_adj_4449), 
            .I3(GND_net), .O(n12));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 counter_2045_2046_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[12]), .I3(n49222), .O(n61[12])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_14 (.CI(n49222), .I0(GND_net), .I1(counter[12]), 
            .CO(n49223));
    SB_LUT4 counter_2045_2046_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[11]), .I3(n49221), .O(n61[11])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_13 (.CI(n49221), .I0(GND_net), .I1(counter[11]), 
            .CO(n49222));
    SB_CARRY add_4970_6 (.CI(n48646), .I0(n19495[3]), .I1(n399), .CO(n48647));
    SB_LUT4 mult_24_i222_2_lut (.I0(\Ki[4] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2045_2046_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[10]), .I3(n49220), .O(n61[10])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_12 (.CI(n49220), .I0(GND_net), .I1(counter[10]), 
            .CO(n49221));
    SB_CARRY mult_24_add_1225_21 (.CI(n48914), .I0(n10958[18]), .I1(GND_net), 
            .CO(n48915));
    SB_LUT4 mult_24_add_1225_20_lut (.I0(GND_net), .I1(n10958[17]), .I2(GND_net), 
            .I3(n48913), .O(n34[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2045_2046_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[9]), .I3(n49219), .O(n61[9])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_20 (.CI(n48913), .I0(n10958[17]), .I1(GND_net), 
            .CO(n48914));
    SB_LUT4 mult_23_i549_2_lut (.I0(\Kp[11] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n816));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_15_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(\motor_state[7] ), 
            .I3(n48290), .O(n207[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4970_5_lut (.I0(GND_net), .I1(n19495[2]), .I2(n326), .I3(n48645), 
            .O(n19186[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4970_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i402_2_lut (.I0(\Ki[8] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597_adj_4482));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i402_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY counter_2045_2046_add_4_11 (.CI(n49219), .I0(GND_net), .I1(counter[9]), 
            .CO(n49220));
    SB_LUT4 counter_2045_2046_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter[8]), .I3(n49218), .O(n61[8])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_10 (.CI(n49218), .I0(GND_net), .I1(counter[8]), 
            .CO(n49219));
    SB_LUT4 counter_2045_2046_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(counter[7]), 
            .I3(n49217), .O(n61[7])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_9 (.CI(n49217), .I0(GND_net), .I1(counter[7]), 
            .CO(n49218));
    SB_LUT4 counter_2045_2046_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(counter[6]), 
            .I3(n49216), .O(n61[6])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_8 (.CI(n49216), .I0(GND_net), .I1(counter[6]), 
            .CO(n49217));
    SB_LUT4 counter_2045_2046_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(counter[5]), 
            .I3(n49215), .O(n61[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4970_5 (.CI(n48645), .I0(n19495[2]), .I1(n326), .CO(n48646));
    SB_LUT4 add_4970_4_lut (.I0(GND_net), .I1(n19495[1]), .I2(n253_adj_4483), 
            .I3(n48644), .O(n19186[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4970_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_7 (.CI(n49215), .I0(GND_net), .I1(counter[5]), 
            .CO(n49216));
    SB_LUT4 counter_2045_2046_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n49214), .O(n61[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_19_lut (.I0(GND_net), .I1(n10958[16]), .I2(GND_net), 
            .I3(n48912), .O(n34[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_6 (.CI(n49214), .I0(GND_net), .I1(counter[4]), 
            .CO(n49215));
    SB_LUT4 counter_2045_2046_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n49213), .O(n61[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_5 (.CI(n49213), .I0(GND_net), .I1(counter[3]), 
            .CO(n49214));
    SB_CARRY sub_15_add_2_9 (.CI(n48290), .I0(setpoint[7]), .I1(\motor_state[7] ), 
            .CO(n48291));
    SB_LUT4 counter_2045_2046_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n49212), .O(n61[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_4 (.CI(n49212), .I0(GND_net), .I1(counter[2]), 
            .CO(n49213));
    SB_LUT4 mult_24_i296_2_lut (.I0(\Ki[6] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 counter_2045_2046_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n49211), .O(n61[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_3 (.CI(n49211), .I0(GND_net), .I1(counter[1]), 
            .CO(n49212));
    SB_CARRY mult_24_add_1225_19 (.CI(n48912), .I0(n10958[16]), .I1(GND_net), 
            .CO(n48913));
    SB_LUT4 counter_2045_2046_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n61[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2045_2046_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4970_4 (.CI(n48644), .I0(n19495[1]), .I1(n253_adj_4483), 
            .CO(n48645));
    SB_LUT4 mult_24_add_1225_18_lut (.I0(GND_net), .I1(n10958[15]), .I2(GND_net), 
            .I3(n48911), .O(n34[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2045_2046_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n49211));
    SB_LUT4 add_4970_3_lut (.I0(GND_net), .I1(n19495[0]), .I2(n180), .I3(n48643), 
            .O(n19186[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4970_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_18 (.CI(n48911), .I0(n10958[15]), .I1(GND_net), 
            .CO(n48912));
    SB_LUT4 mult_24_add_1225_17_lut (.I0(GND_net), .I1(n10958[14]), .I2(GND_net), 
            .I3(n48910), .O(n34[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4970_3 (.CI(n48643), .I0(n19495[0]), .I1(n180), .CO(n48644));
    SB_CARRY mult_24_add_1225_17 (.CI(n48910), .I0(n10958[14]), .I1(GND_net), 
            .CO(n48911));
    SB_LUT4 add_4970_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n19186[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4970_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4970_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n48643));
    SB_LUT4 add_5070_8_lut (.I0(GND_net), .I1(n20432[5]), .I2(n560), .I3(n48642), 
            .O(n20336[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_16_lut (.I0(GND_net), .I1(n10958[13]), .I2(n1096), 
            .I3(n48909), .O(n34[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5070_7_lut (.I0(GND_net), .I1(n20432[4]), .I2(n487), .I3(n48641), 
            .O(n20336[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_7 (.CI(n48641), .I0(n20432[4]), .I1(n487), .CO(n48642));
    SB_CARRY mult_24_add_1225_16 (.CI(n48909), .I0(n10958[13]), .I1(n1096), 
            .CO(n48910));
    SB_LUT4 add_5070_6_lut (.I0(GND_net), .I1(n20432[3]), .I2(n414), .I3(n48640), 
            .O(n20336[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_15_lut (.I0(GND_net), .I1(n10958[12]), .I2(n1023), 
            .I3(n48908), .O(n34[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_6 (.CI(n48640), .I0(n20432[3]), .I1(n414), .CO(n48641));
    SB_CARRY mult_24_add_1225_15 (.CI(n48908), .I0(n10958[12]), .I1(n1023), 
            .CO(n48909));
    SB_LUT4 add_5070_5_lut (.I0(GND_net), .I1(n20432[2]), .I2(n341), .I3(n48639), 
            .O(n20336[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_14_lut (.I0(GND_net), .I1(n10958[11]), .I2(n950), 
            .I3(n48907), .O(n34[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_14 (.CI(n48907), .I0(n10958[11]), .I1(n950), 
            .CO(n48908));
    SB_CARRY add_5070_5 (.CI(n48639), .I0(n20432[2]), .I1(n341), .CO(n48640));
    SB_LUT4 add_5070_4_lut (.I0(GND_net), .I1(n20432[1]), .I2(n268), .I3(n48638), 
            .O(n20336[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_4 (.CI(n48638), .I0(n20432[1]), .I1(n268), .CO(n48639));
    SB_LUT4 mult_24_add_1225_13_lut (.I0(GND_net), .I1(n10958[10]), .I2(n877), 
            .I3(n48906), .O(n34[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5070_3_lut (.I0(GND_net), .I1(n20432[0]), .I2(n195), .I3(n48637), 
            .O(n20336[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_3 (.CI(n48637), .I0(n20432[0]), .I1(n195), .CO(n48638));
    SB_LUT4 mult_23_i598_2_lut (.I0(\Kp[12] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i598_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_24_add_1225_13 (.CI(n48906), .I0(n10958[10]), .I1(n877), 
            .CO(n48907));
    SB_LUT4 i48807_4_lut (.I0(n30), .I1(n10), .I2(n35_adj_4486), .I3(n63577), 
            .O(n65869));   // verilog/motorControl.v(63[16:31])
    defparam i48807_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47312_3_lut (.I0(n65190), .I1(n455[15]), .I2(n31_adj_4473), 
            .I3(GND_net), .O(n64374));   // verilog/motorControl.v(63[16:31])
    defparam i47312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5070_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n20336[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49028_4_lut (.I0(n64374), .I1(n65869), .I2(n35_adj_4486), 
            .I3(n63586), .O(n66090));   // verilog/motorControl.v(63[16:31])
    defparam i49028_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49029_3_lut (.I0(n66090), .I1(n455[18]), .I2(n37_adj_4487), 
            .I3(GND_net), .O(n66091));   // verilog/motorControl.v(63[16:31])
    defparam i49029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_add_1225_12_lut (.I0(GND_net), .I1(n10958[9]), .I2(n804), 
            .I3(n48905), .O(n34[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n48637));
    SB_LUT4 add_4993_12_lut (.I0(GND_net), .I1(n19756[9]), .I2(n840), 
            .I3(n48636), .O(n19495[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4993_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_17_i10_3_lut (.I0(n233[5]), .I1(n233[6]), .I2(n13), 
            .I3(GND_net), .O(n10_adj_4489));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_17_i30_3_lut (.I0(n12), .I1(n233[17]), .I2(n35_adj_4448), 
            .I3(GND_net), .O(n30_adj_4490));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_24_add_1225_12 (.CI(n48905), .I0(n10958[9]), .I1(n804), 
            .CO(n48906));
    SB_LUT4 mult_24_i451_2_lut (.I0(\Ki[9] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670_adj_4491));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_add_1225_11_lut (.I0(GND_net), .I1(n10958[8]), .I2(n731), 
            .I3(n48904), .O(n34[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4993_11_lut (.I0(GND_net), .I1(n19756[8]), .I2(n767), 
            .I3(n48635), .O(n19495[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4993_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i271_2_lut (.I0(\Ki[5] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i271_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4993_11 (.CI(n48635), .I0(n19756[8]), .I1(n767), .CO(n48636));
    SB_LUT4 add_4993_10_lut (.I0(GND_net), .I1(n19756[7]), .I2(n694), 
            .I3(n48634), .O(n19495[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4993_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47901_4_lut (.I0(n13), .I1(n11), .I2(n9_c), .I3(n64043), 
            .O(n64963));
    defparam i47901_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i47893_4_lut (.I0(n19), .I1(n17_adj_4458), .I2(n15_adj_4471), 
            .I3(n64963), .O(n64955));
    defparam i47893_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY mult_24_add_1225_11 (.CI(n48904), .I0(n10958[8]), .I1(n731), 
            .CO(n48905));
    SB_LUT4 mult_24_add_1225_10_lut (.I0(GND_net), .I1(n10958[7]), .I2(n658), 
            .I3(n48903), .O(n34[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4993_10 (.CI(n48634), .I0(n19756[7]), .I1(n694), .CO(n48635));
    SB_LUT4 add_4993_9_lut (.I0(GND_net), .I1(n19756[6]), .I2(n621), .I3(n48633), 
            .O(n19495[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4993_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_10 (.CI(n48903), .I0(n10958[7]), .I1(n658), 
            .CO(n48904));
    SB_LUT4 i46635_4_lut (.I0(n455[8]), .I1(n455[4]), .I2(n28[8]), .I3(n28[4]), 
            .O(n63697));
    defparam i46635_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i48885_4_lut (.I0(n25_adj_4446), .I1(n23_adj_4445), .I2(n21_adj_4460), 
            .I3(n64955), .O(n65947));
    defparam i48885_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_15_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(\motor_state[6] ), 
            .I3(n48289), .O(n207[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4993_9 (.CI(n48633), .I0(n19756[6]), .I1(n621), .CO(n48634));
    SB_LUT4 mult_24_add_1225_9_lut (.I0(GND_net), .I1(n10958[6]), .I2(n585), 
            .I3(n48902), .O(n34[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4993_8_lut (.I0(GND_net), .I1(n19756[5]), .I2(n548), .I3(n48632), 
            .O(n19495[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4993_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48323_4_lut (.I0(n31_adj_4442), .I1(n29_adj_4441), .I2(n27_adj_4474), 
            .I3(n65947), .O(n65385));
    defparam i48323_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_24_i500_2_lut (.I0(\Ki[10] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_4492));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i500_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_15_add_2_8 (.CI(n48289), .I0(setpoint[6]), .I1(\motor_state[6] ), 
            .CO(n48290));
    SB_LUT4 i49024_4_lut (.I0(n37_adj_4447), .I1(n35_adj_4448), .I2(n33_adj_4449), 
            .I3(n65385), .O(n66086));
    defparam i49024_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_23_i647_2_lut (.I0(\Kp[13] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i647_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_24_add_1225_9 (.CI(n48902), .I0(n10958[6]), .I1(n585), 
            .CO(n48903));
    SB_LUT4 mult_24_i345_2_lut (.I0(\Ki[7] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i549_2_lut (.I0(\Ki[11] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_4493));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i549_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4993_8 (.CI(n48632), .I0(n19756[5]), .I1(n548), .CO(n48633));
    SB_LUT4 mult_24_i320_2_lut (.I0(\Ki[6] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4494));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47608_3_lut (.I0(n455[9]), .I1(n63697), .I2(n28[9]), .I3(GND_net), 
            .O(n64670));
    defparam i47608_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 LessThan_17_i16_3_lut (.I0(n233[9]), .I1(n233[21]), .I2(n43_adj_4440), 
            .I3(GND_net), .O(n16_adj_4495));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i598_2_lut (.I0(\Ki[12] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_4496));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4993_7_lut (.I0(GND_net), .I1(n19756[4]), .I2(n475_adj_4494), 
            .I3(n48631), .O(n19495[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4993_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i647_2_lut (.I0(\Ki[13] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962_adj_4497));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i696_2_lut (.I0(\Kp[14] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_add_1225_8_lut (.I0(GND_net), .I1(n10958[5]), .I2(n512), 
            .I3(n48901), .O(n34[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48589_3_lut (.I0(n6_adj_4498), .I1(n233[10]), .I2(n21_adj_4460), 
            .I3(GND_net), .O(n65651));   // verilog/motorControl.v(56[14:36])
    defparam i48589_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4993_7 (.CI(n48631), .I0(n19756[4]), .I1(n475_adj_4494), 
            .CO(n48632));
    SB_LUT4 i48590_3_lut (.I0(n65651), .I1(n233[11]), .I2(n23_adj_4445), 
            .I3(GND_net), .O(n65652));   // verilog/motorControl.v(56[14:36])
    defparam i48590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4993_6_lut (.I0(GND_net), .I1(n19756[3]), .I2(n402), .I3(n48630), 
            .O(n19495[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4993_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(\motor_state[5] ), 
            .I3(n48288), .O(n207[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4993_6 (.CI(n48630), .I0(n19756[3]), .I1(n402), .CO(n48631));
    SB_LUT4 mult_24_i696_2_lut (.I0(\Ki[14] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_4499));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i696_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_24_add_1225_8 (.CI(n48901), .I0(n10958[5]), .I1(n512), 
            .CO(n48902));
    SB_LUT4 mult_24_i745_2_lut (.I0(\Ki[15] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i8_3_lut (.I0(n233[4]), .I1(n233[8]), .I2(n17_adj_4458), 
            .I3(GND_net), .O(n8_adj_4500));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_add_1225_7_lut (.I0(GND_net), .I1(n10958[4]), .I2(n439), 
            .I3(n48900), .O(n34[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4993_5_lut (.I0(GND_net), .I1(n19756[2]), .I2(n329), .I3(n48629), 
            .O(n19495[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4993_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_28_i21_rep_89_2_lut (.I0(n455[10]), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n67235));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i21_rep_89_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_24_add_1225_7 (.CI(n48900), .I0(n10958[4]), .I1(n439), 
            .CO(n48901));
    SB_CARRY add_4993_5 (.CI(n48629), .I0(n19756[2]), .I1(n329), .CO(n48630));
    SB_LUT4 add_4993_4_lut (.I0(GND_net), .I1(n19756[1]), .I2(n256_adj_4480), 
            .I3(n48628), .O(n19495[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4993_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_add_1225_6_lut (.I0(GND_net), .I1(n10958[3]), .I2(n366_adj_4478), 
            .I3(n48899), .O(n34[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4993_4 (.CI(n48628), .I0(n19756[1]), .I1(n256_adj_4480), 
            .CO(n48629));
    SB_LUT4 LessThan_17_i24_3_lut (.I0(n16_adj_4495), .I1(n233[22]), .I2(n45_adj_4438), 
            .I3(GND_net), .O(n24_adj_4501));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_24_add_1225_6 (.CI(n48899), .I0(n10958[3]), .I1(n366_adj_4478), 
            .CO(n48900));
    SB_LUT4 add_4993_3_lut (.I0(GND_net), .I1(n19756[0]), .I2(n183), .I3(n48627), 
            .O(n19495[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4993_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_7 (.CI(n48288), .I0(setpoint[5]), .I1(\motor_state[5] ), 
            .CO(n48289));
    SB_LUT4 sub_15_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(\motor_state[4] ), 
            .I3(n48287), .O(n207[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46879_4_lut (.I0(n43_adj_4440), .I1(n25_adj_4446), .I2(n23_adj_4445), 
            .I3(n64027), .O(n63941));
    defparam i46879_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_i745_2_lut (.I0(\Kp[15] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_4502));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48410_4_lut (.I0(n24_adj_4501), .I1(n8_adj_4500), .I2(n45_adj_4438), 
            .I3(n63935), .O(n65472));   // verilog/motorControl.v(56[14:36])
    defparam i48410_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49003_3_lut (.I0(n66091), .I1(n455[19]), .I2(n39_adj_4503), 
            .I3(GND_net), .O(n66065));   // verilog/motorControl.v(63[16:31])
    defparam i49003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47270_3_lut (.I0(n65652), .I1(n233[12]), .I2(n25_adj_4446), 
            .I3(GND_net), .O(n64332));   // verilog/motorControl.v(56[14:36])
    defparam i47270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i369_2_lut (.I0(\Ki[7] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i4_4_lut (.I0(n233[0]), .I1(n233[1]), .I2(IntegralLimit[1]), 
            .I3(IntegralLimit[0]), .O(n4_adj_4504));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 mux_21_i17_3_lut (.I0(n233[16]), .I1(n285[16]), .I2(n284), 
            .I3(GND_net), .O(n310[16]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i17_3_lut (.I0(n310[16]), .I1(IntegralLimit[16]), .I2(n258), 
            .I3(GND_net), .O(n335[16]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_add_1225_5_lut (.I0(GND_net), .I1(n10958[2]), .I2(n293), 
            .I3(n48898), .O(n34[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4993_3 (.CI(n48627), .I0(n19756[0]), .I1(n183), .CO(n48628));
    SB_LUT4 mult_24_i394_2_lut (.I0(\Ki[8] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48585_3_lut (.I0(n4_adj_4504), .I1(n233[13]), .I2(n27_adj_4474), 
            .I3(GND_net), .O(n65647));   // verilog/motorControl.v(56[14:36])
    defparam i48585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48586_3_lut (.I0(n65647), .I1(n233[14]), .I2(n29_adj_4441), 
            .I3(GND_net), .O(n65648));   // verilog/motorControl.v(56[14:36])
    defparam i48586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i81_2_lut (.I0(\Ki[1] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46938_4_lut (.I0(n33_adj_4449), .I1(n31_adj_4442), .I2(n29_adj_4441), 
            .I3(n64016), .O(n64000));
    defparam i46938_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i34_2_lut (.I0(\Ki[0] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48903_4_lut (.I0(n30_adj_4490), .I1(n10_adj_4489), .I2(n35_adj_4448), 
            .I3(n63990), .O(n65965));   // verilog/motorControl.v(56[14:36])
    defparam i48903_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47272_3_lut (.I0(n65648), .I1(n233[15]), .I2(n31_adj_4442), 
            .I3(GND_net), .O(n64334));   // verilog/motorControl.v(56[14:36])
    defparam i47272_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4993_2_lut (.I0(GND_net), .I1(n41_adj_4469), .I2(n110), 
            .I3(GND_net), .O(n19495[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4993_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_6 (.CI(n48287), .I0(setpoint[4]), .I1(\motor_state[4] ), 
            .CO(n48288));
    SB_CARRY mult_24_add_1225_5 (.CI(n48898), .I0(n10958[2]), .I1(n293), 
            .CO(n48899));
    SB_CARRY add_4993_2 (.CI(GND_net), .I0(n41_adj_4469), .I1(n110), .CO(n48627));
    SB_LUT4 i47604_4_lut (.I0(n455[11]), .I1(n67235), .I2(n28[11]), .I3(n64670), 
            .O(n64666));
    defparam i47604_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 LessThan_28_i25_rep_84_2_lut (.I0(n455[12]), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n67230));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i25_rep_84_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_add_1225_4_lut (.I0(GND_net), .I1(n10958[1]), .I2(n220), 
            .I3(n48897), .O(n34[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_4 (.CI(n48897), .I0(n10958[1]), .I1(n220), 
            .CO(n48898));
    SB_LUT4 mult_24_i418_2_lut (.I0(\Ki[8] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i443_2_lut (.I0(\Ki[9] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49114_4_lut (.I0(n64334), .I1(n65965), .I2(n35_adj_4448), 
            .I3(n64000), .O(n66176));   // verilog/motorControl.v(56[14:36])
    defparam i49114_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 n9972_bdd_4_lut_49731 (.I0(n9972), .I1(n63118), .I2(setpoint[22]), 
            .I3(n4744), .O(n66741));
    defparam n9972_bdd_4_lut_49731.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_24_add_1225_3_lut (.I0(GND_net), .I1(n10958[0]), .I2(n147), 
            .I3(n48896), .O(n34[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_24_add_1225_3 (.CI(n48896), .I0(n10958[0]), .I1(n147), 
            .CO(n48897));
    SB_LUT4 i49115_3_lut (.I0(n66176), .I1(n233[18]), .I2(n37_adj_4447), 
            .I3(GND_net), .O(n66177));   // verilog/motorControl.v(56[14:36])
    defparam i49115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i467_2_lut (.I0(\Ki[9] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_add_1225_2_lut (.I0(GND_net), .I1(n5), .I2(n74), .I3(GND_net), 
            .O(n34[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_24_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i130_2_lut (.I0(\Ki[2] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i516_2_lut (.I0(\Ki[10] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i492_2_lut (.I0(\Ki[10] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46493_4_lut (.I0(n43_adj_4431), .I1(n41_adj_4507), .I2(n39_adj_4503), 
            .I3(n66060), .O(n63555));
    defparam i46493_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_24_i179_2_lut (.I0(\Ki[3] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i179_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_24_add_1225_2 (.CI(GND_net), .I0(n5), .I1(n74), .CO(n48896));
    SB_LUT4 i49087_3_lut (.I0(n66177), .I1(n233[19]), .I2(n39), .I3(GND_net), 
            .O(n66149));   // verilog/motorControl.v(56[14:36])
    defparam i49087_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_15_add_2_12 (.CI(n48293), .I0(setpoint[10]), .I1(\motor_state[10] ), 
            .CO(n48294));
    SB_CARRY sub_15_add_2_5 (.CI(n48286), .I0(setpoint[3]), .I1(\motor_state[3] ), 
            .CO(n48287));
    SB_CARRY sub_15_add_2_4 (.CI(n48285), .I0(setpoint[2]), .I1(n3), .CO(n48286));
    SB_CARRY sub_15_add_2_3 (.CI(n48284), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n48285));
    SB_CARRY sub_15_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n48284));
    SB_LUT4 mult_24_i228_2_lut (.I0(\Ki[4] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_28_i16_3_lut (.I0(n28[9]), .I1(n28[21]), .I2(n455[21]), 
            .I3(GND_net), .O(n16_adj_4508));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_24_i277_2_lut (.I0(\Ki[5] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9972_bdd_4_lut_49879 (.I0(n9972), .I1(n63140), .I2(setpoint[1]), 
            .I3(n4744), .O(n67017));
    defparam n9972_bdd_4_lut_49879.LUT_INIT = 16'he4aa;
    SB_LUT4 n67017_bdd_4_lut (.I0(n67017), .I1(n535[1]), .I2(n455[1]), 
            .I3(n4744), .O(n67020));
    defparam n67017_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i46584_4_lut (.I0(n455[21]), .I1(n455[9]), .I2(n28[21]), .I3(n28[9]), 
            .O(n63646));
    defparam i46584_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mult_24_i326_2_lut (.I0(\Ki[6] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_4509));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9972_bdd_4_lut_49870 (.I0(n9972), .I1(n63139), .I2(setpoint[0]), 
            .I3(n4744), .O(n67011));
    defparam n9972_bdd_4_lut_49870.LUT_INIT = 16'he4aa;
    SB_LUT4 mult_23_i296_2_lut (.I0(\Kp[6] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n439_adj_4510));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46892_4_lut (.I0(n43_adj_4440), .I1(n41), .I2(n39), .I3(n66086), 
            .O(n63954));
    defparam i46892_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48745_4_lut (.I0(n64372), .I1(n65480), .I2(n45), .I3(n63552), 
            .O(n65807));   // verilog/motorControl.v(63[16:31])
    defparam i48745_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 n67011_bdd_4_lut (.I0(n67011), .I1(n535[0]), .I2(n455[0]), 
            .I3(n4744), .O(n67014));
    defparam n67011_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_28_i8_3_lut (.I0(n28[4]), .I1(n28[8]), .I2(n455[8]), 
            .I3(GND_net), .O(n8_adj_4511));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i8_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_28_i24_3_lut (.I0(n16_adj_4508), .I1(n28[22]), .I2(n455[22]), 
            .I3(GND_net), .O(n24_adj_4512));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46654_4_lut (.I0(n455[3]), .I1(n455[2]), .I2(n28[3]), .I3(n28[2]), 
            .O(n63716));
    defparam i46654_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_28_i9_rep_82_2_lut (.I0(n455[4]), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n67228));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i9_rep_82_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46651_4_lut (.I0(n455[5]), .I1(n67228), .I2(n28[5]), .I3(n63716), 
            .O(n63713));
    defparam i46651_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_28_i13_rep_110_2_lut (.I0(n455[6]), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n67256));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i13_rep_110_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48959_4_lut (.I0(n64332), .I1(n65472), .I2(n45_adj_4438), 
            .I3(n63941), .O(n66021));   // verilog/motorControl.v(56[14:36])
    defparam i48959_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47278_3_lut (.I0(n66149), .I1(n233[20]), .I2(n41), .I3(GND_net), 
            .O(n64340));   // verilog/motorControl.v(56[14:36])
    defparam i47278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48961_4_lut (.I0(n64340), .I1(n66021), .I2(n45_adj_4438), 
            .I3(n63954), .O(n66023));   // verilog/motorControl.v(56[14:36])
    defparam i48961_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_24_i565_2_lut (.I0(\Ki[11] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48962_3_lut (.I0(n66023), .I1(IntegralLimit[23]), .I2(n233[23]), 
            .I3(GND_net), .O(n258));   // verilog/motorControl.v(56[14:36])
    defparam i48962_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_24_i541_2_lut (.I0(\Ki[11] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i83_2_lut (.I0(\Kp[1] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n122));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i41_2_lut (.I0(n233[20]), .I1(n285[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4513));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i36_2_lut (.I0(\Kp[0] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n53));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i39_2_lut (.I0(n233[19]), .I1(n285[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4514));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i132_2_lut (.I0(\Kp[2] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n195));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i45_2_lut (.I0(n233[22]), .I1(n285[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4515));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i590_2_lut (.I0(\Ki[12] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i181_2_lut (.I0(\Kp[3] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n268));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i639_2_lut (.I0(\Ki[13] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i43_2_lut (.I0(n233[21]), .I1(n285[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4516));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i230_2_lut (.I0(\Kp[4] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n341));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i688_2_lut (.I0(\Ki[14] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i279_2_lut (.I0(\Kp[5] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n414));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n66741_bdd_4_lut (.I0(n66741), .I1(n535[22]), .I2(n455[22]), 
            .I3(n4744), .O(n66744));
    defparam n66741_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_19_i37_2_lut (.I0(n233[18]), .I1(n285[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4517));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i29_2_lut (.I0(n233[14]), .I1(n285[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4518));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i328_2_lut (.I0(\Kp[6] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n487));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i31_2_lut (.I0(n233[15]), .I1(n285[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4519));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_21_i1_3_lut (.I0(n233[0]), .I1(n285[0]), .I2(n284), .I3(GND_net), 
            .O(n310[0]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i1_3_lut (.I0(n310[0]), .I1(IntegralLimit[0]), .I2(n258), 
            .I3(GND_net), .O(n335[0]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i737_2_lut (.I0(\Ki[15] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i23_2_lut (.I0(n233[11]), .I1(n285[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4520));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_23_i377_2_lut (.I0(\Kp[7] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n560));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i13_3_lut (.I0(n233[12]), .I1(n285[12]), .I2(n284), 
            .I3(GND_net), .O(n310[12]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i13_3_lut (.I0(n310[12]), .I1(IntegralLimit[12]), .I2(n258), 
            .I3(GND_net), .O(n335[12]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i25_2_lut (.I0(n233[12]), .I1(n285[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4521));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i73_2_lut (.I0(\Ki[1] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i26_2_lut (.I0(\Ki[0] ), .I1(n335[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i35_2_lut (.I0(n233[17]), .I1(n285[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4522));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i122_2_lut (.I0(\Ki[2] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i171_2_lut (.I0(\Ki[3] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_4483));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i33_2_lut (.I0(n233[16]), .I1(n285[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4523));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i220_2_lut (.I0(\Ki[4] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i11_2_lut (.I0(n233[5]), .I1(n285[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4524));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i13_2_lut (.I0(n233[6]), .I1(n285[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4525));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i269_2_lut (.I0(\Ki[5] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i15_2_lut (.I0(n233[7]), .I1(n285[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4526));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i318_2_lut (.I0(\Ki[6] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_4481));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i367_2_lut (.I0(\Ki[7] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i27_2_lut (.I0(n233[13]), .I1(n285[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4527));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i416_2_lut (.I0(\Ki[8] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i24_3_lut (.I0(n233[23]), .I1(n285[23]), .I2(n284), 
            .I3(GND_net), .O(n310[23]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i24_3_lut (.I0(n310[23]), .I1(IntegralLimit[23]), .I2(n258), 
            .I3(GND_net), .O(n335[23]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i9_2_lut (.I0(n233[4]), .I1(n285[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4529));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i17_2_lut (.I0(n233[8]), .I1(n285[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4530));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i19_2_lut (.I0(n233[9]), .I1(n285[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4531));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_19_i21_2_lut (.I0(n233[10]), .I1(n285[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4532));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48185_4_lut (.I0(n455[7]), .I1(n67256), .I2(n28[7]), .I3(n63713), 
            .O(n65247));
    defparam i48185_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i46838_4_lut (.I0(n21_adj_4532), .I1(n19_adj_4531), .I2(n17_adj_4530), 
            .I3(n9_adj_4529), .O(n63900));
    defparam i46838_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46824_4_lut (.I0(n27_adj_4527), .I1(n15_adj_4526), .I2(n13_adj_4525), 
            .I3(n11_adj_4524), .O(n63886));
    defparam i46824_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_19_i12_3_lut (.I0(n285[7]), .I1(n285[16]), .I2(n33_adj_4523), 
            .I3(GND_net), .O(n12_adj_4533));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i10_3_lut (.I0(n285[5]), .I1(n285[6]), .I2(n13_adj_4525), 
            .I3(GND_net), .O(n10_adj_4534));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_19_i30_3_lut (.I0(n12_adj_4533), .I1(n285[17]), .I2(n35_adj_4522), 
            .I3(GND_net), .O(n30_adj_4535));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i465_2_lut (.I0(\Ki[9] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47801_4_lut (.I0(n13_adj_4525), .I1(n11_adj_4524), .I2(n9_adj_4529), 
            .I3(n63931), .O(n64863));
    defparam i47801_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_24_i514_2_lut (.I0(\Ki[10] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47793_4_lut (.I0(n19_adj_4531), .I1(n17_adj_4530), .I2(n15_adj_4526), 
            .I3(n64863), .O(n64855));
    defparam i47793_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_24_i375_2_lut (.I0(\Ki[7] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_4536));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48869_4_lut (.I0(n25_adj_4521), .I1(n23_adj_4520), .I2(n21_adj_4532), 
            .I3(n64855), .O(n65931));
    defparam i48869_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47318_3_lut (.I0(n66065), .I1(n455[20]), .I2(n41_adj_4507), 
            .I3(GND_net), .O(n64380));   // verilog/motorControl.v(63[16:31])
    defparam i47318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48975_4_lut (.I0(n64380), .I1(n65807), .I2(n45), .I3(n63555), 
            .O(n66037));   // verilog/motorControl.v(63[16:31])
    defparam i48975_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_11_i45_2_lut (.I0(setpoint[22]), .I1(n535[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4537));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i37_2_lut (.I0(setpoint[18]), .I1(n535[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4538));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i41_2_lut (.I0(setpoint[20]), .I1(n535[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4540));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i43_2_lut (.I0(setpoint[21]), .I1(n535[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4541));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5014_11_lut (.I0(GND_net), .I1(n19973[8]), .I2(n770), 
            .I3(n48611), .O(n19756[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5014_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i29_2_lut (.I0(setpoint[14]), .I1(n535[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4543));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_28_i17_rep_107_2_lut (.I0(n455[8]), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n67253));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i17_rep_107_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i31_2_lut (.I0(setpoint[15]), .I1(n535[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4544));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i33_2_lut (.I0(setpoint[16]), .I1(n535[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4545));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5014_10_lut (.I0(GND_net), .I1(n19973[7]), .I2(n697), 
            .I3(n48610), .O(n19756[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5014_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_11_i39_2_lut (.I0(setpoint[19]), .I1(n535[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4546));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i35_2_lut (.I0(setpoint[17]), .I1(n535[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4548));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5014_10 (.CI(n48610), .I0(n19973[7]), .I1(n697), .CO(n48611));
    SB_LUT4 i48257_4_lut (.I0(n31_adj_4519), .I1(n29_adj_4518), .I2(n27_adj_4527), 
            .I3(n65931), .O(n65319));
    defparam i48257_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut (.I0(control_mode[2]), .I1(control_update), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4549));
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i49018_4_lut (.I0(n37_adj_4517), .I1(n35_adj_4522), .I2(n33_adj_4523), 
            .I3(n65319), .O(n66080));
    defparam i49018_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i47612_4_lut (.I0(n455[9]), .I1(n67253), .I2(n28[9]), .I3(n65247), 
            .O(n64674));
    defparam i47612_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 mult_24_i424_2_lut (.I0(\Ki[8] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_19_i16_3_lut (.I0(n285[9]), .I1(n285[21]), .I2(n43_adj_4516), 
            .I3(GND_net), .O(n16_adj_4550));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5014_9_lut (.I0(GND_net), .I1(n19973[6]), .I2(n624), .I3(n48609), 
            .O(n19756[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5014_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut (.I0(n55181), .I1(control_mode[3]), .I2(n105), .I3(n6_adj_4549), 
            .O(n25015));
    defparam i4_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i47065_4_lut (.I0(n21_adj_4551), .I1(n19_adj_4552), .I2(n17_adj_4553), 
            .I3(n9_adj_4554), .O(n64127));
    defparam i47065_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48581_3_lut (.I0(n6_adj_4555), .I1(n285[10]), .I2(n21_adj_4532), 
            .I3(GND_net), .O(n65643));   // verilog/motorControl.v(58[23:46])
    defparam i48581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47046_4_lut (.I0(n27_adj_4556), .I1(n15_adj_4557), .I2(n13_adj_4558), 
            .I3(n11_adj_4559), .O(n64108));
    defparam i47046_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_11_i12_3_lut (.I0(n535[7]), .I1(n535[16]), .I2(n33_adj_4545), 
            .I3(GND_net), .O(n12_adj_4560));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i10_3_lut (.I0(n535[5]), .I1(n535[6]), .I2(n13_adj_4558), 
            .I3(GND_net), .O(n10_adj_4561));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i563_2_lut (.I0(\Ki[11] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i30_3_lut (.I0(n12_adj_4560), .I1(n535[17]), .I2(n35_adj_4548), 
            .I3(GND_net), .O(n30_adj_4562));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i612_2_lut (.I0(\Ki[12] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i5_3_lut (.I0(n233[4]), .I1(n285[4]), .I2(n284), .I3(GND_net), 
            .O(n310[4]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48582_3_lut (.I0(n65643), .I1(n285[11]), .I2(n23_adj_4520), 
            .I3(GND_net), .O(n65644));   // verilog/motorControl.v(58[23:46])
    defparam i48582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i5_3_lut (.I0(n310[4]), .I1(IntegralLimit[4]), .I2(n258), 
            .I3(GND_net), .O(n335[4]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4527_23_lut (.I0(GND_net), .I1(n12488[20]), .I2(GND_net), 
            .I3(n48883), .O(n10958[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i57_2_lut (.I0(\Ki[1] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4527_22_lut (.I0(GND_net), .I1(n12488[19]), .I2(GND_net), 
            .I3(n48882), .O(n10958[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47981_4_lut (.I0(n13_adj_4558), .I1(n11_adj_4559), .I2(n9_adj_4554), 
            .I3(n64177), .O(n65043));
    defparam i47981_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i47965_4_lut (.I0(n19_adj_4552), .I1(n17_adj_4553), .I2(n15_adj_4557), 
            .I3(n65043), .O(n65027));
    defparam i47965_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_19_i8_3_lut (.I0(n285[4]), .I1(n285[8]), .I2(n17_adj_4530), 
            .I3(GND_net), .O(n8_adj_4563));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48895_4_lut (.I0(n25_adj_4564), .I1(n23_adj_4565), .I2(n21_adj_4551), 
            .I3(n65027), .O(n65957));
    defparam i48895_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_19_i24_3_lut (.I0(n16_adj_4550), .I1(n285[22]), .I2(n45_adj_4515), 
            .I3(GND_net), .O(n24_adj_4566));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4980_13_lut (.I0(GND_net), .I1(n19612[10]), .I2(n910_adj_4567), 
            .I3(n49108), .O(n19326[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4980_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5014_9 (.CI(n48609), .I0(n19973[6]), .I1(n624), .CO(n48610));
    SB_LUT4 add_5014_8_lut (.I0(GND_net), .I1(n19973[5]), .I2(n551_adj_4568), 
            .I3(n48608), .O(n19756[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5014_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4980_12_lut (.I0(GND_net), .I1(n19612[9]), .I2(n837_adj_4569), 
            .I3(n49107), .O(n19326[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4980_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_22 (.CI(n48882), .I0(n12488[19]), .I1(GND_net), 
            .CO(n48883));
    SB_CARRY add_5014_8 (.CI(n48608), .I0(n19973[5]), .I1(n551_adj_4568), 
            .CO(n48609));
    SB_LUT4 add_4527_21_lut (.I0(GND_net), .I1(n12488[18]), .I2(GND_net), 
            .I3(n48881), .O(n10958[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5014_7_lut (.I0(GND_net), .I1(n19973[4]), .I2(n478_adj_4570), 
            .I3(n48607), .O(n19756[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5014_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5014_7 (.CI(n48607), .I0(n19973[4]), .I1(n478_adj_4570), 
            .CO(n48608));
    SB_CARRY add_4980_12 (.CI(n49107), .I0(n19612[9]), .I1(n837_adj_4569), 
            .CO(n49108));
    SB_LUT4 add_4980_11_lut (.I0(GND_net), .I1(n19612[8]), .I2(n764_adj_4571), 
            .I3(n49106), .O(n19326[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4980_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4980_11 (.CI(n49106), .I0(n19612[8]), .I1(n764_adj_4571), 
            .CO(n49107));
    SB_LUT4 add_4980_10_lut (.I0(GND_net), .I1(n19612[7]), .I2(n691_adj_4572), 
            .I3(n49105), .O(n19326[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4980_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4980_10 (.CI(n49105), .I0(n19612[7]), .I1(n691_adj_4572), 
            .CO(n49106));
    SB_LUT4 i48351_4_lut (.I0(n31_adj_4544), .I1(n29_adj_4543), .I2(n27_adj_4556), 
            .I3(n65957), .O(n65413));
    defparam i48351_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 add_4980_9_lut (.I0(GND_net), .I1(n19612[6]), .I2(n618_adj_4573), 
            .I3(n49104), .O(n19326[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4980_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4980_9 (.CI(n49104), .I0(n19612[6]), .I1(n618_adj_4573), 
            .CO(n49105));
    SB_LUT4 add_4980_8_lut (.I0(GND_net), .I1(n19612[5]), .I2(n545_adj_4574), 
            .I3(n49103), .O(n19326[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4980_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4980_8 (.CI(n49103), .I0(n19612[5]), .I1(n545_adj_4574), 
            .CO(n49104));
    SB_LUT4 add_4980_7_lut (.I0(GND_net), .I1(n19612[4]), .I2(n472_adj_4575), 
            .I3(n49102), .O(n19326[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4980_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4980_7 (.CI(n49102), .I0(n19612[4]), .I1(n472_adj_4575), 
            .CO(n49103));
    SB_LUT4 add_4980_6_lut (.I0(GND_net), .I1(n19612[3]), .I2(n399_adj_4576), 
            .I3(n49101), .O(n19326[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4980_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49026_4_lut (.I0(n37_adj_4538), .I1(n35_adj_4548), .I2(n33_adj_4545), 
            .I3(n65413), .O(n66088));
    defparam i49026_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_11_i16_3_lut (.I0(n535[9]), .I1(n535[21]), .I2(n43_adj_4541), 
            .I3(GND_net), .O(n16_adj_4577));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i10_2_lut (.I0(\Ki[0] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i345_2_lut (.I0(\Kp[7] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n512_adj_4578));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48611_4_lut (.I0(n455[11]), .I1(n67235), .I2(n28[11]), .I3(n64674), 
            .O(n65673));
    defparam i48611_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_4980_6 (.CI(n49101), .I0(n19612[3]), .I1(n399_adj_4576), 
            .CO(n49102));
    SB_LUT4 mult_23_i57_2_lut (.I0(\Kp[1] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4579));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i10_2_lut (.I0(\Kp[0] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4580));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4980_5_lut (.I0(GND_net), .I1(n19612[2]), .I2(n326_adj_4581), 
            .I3(n49100), .O(n19326[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4980_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5014_6_lut (.I0(GND_net), .I1(n19973[3]), .I2(n405), .I3(n48606), 
            .O(n19756[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5014_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_21 (.CI(n48881), .I0(n12488[18]), .I1(GND_net), 
            .CO(n48882));
    SB_CARRY add_4980_5 (.CI(n49100), .I0(n19612[2]), .I1(n326_adj_4581), 
            .CO(n49101));
    SB_CARRY add_5014_6 (.CI(n48606), .I0(n19973[3]), .I1(n405), .CO(n48607));
    SB_LUT4 add_5014_5_lut (.I0(GND_net), .I1(n19973[2]), .I2(n332), .I3(n48605), 
            .O(n19756[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5014_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4527_20_lut (.I0(GND_net), .I1(n12488[17]), .I2(GND_net), 
            .I3(n48880), .O(n10958[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4980_4_lut (.I0(GND_net), .I1(n19612[1]), .I2(n253_adj_4582), 
            .I3(n49099), .O(n19326[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4980_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4980_4 (.CI(n49099), .I0(n19612[1]), .I1(n253_adj_4582), 
            .CO(n49100));
    SB_LUT4 add_4980_3_lut (.I0(GND_net), .I1(n19612[0]), .I2(n180_adj_4583), 
            .I3(n49098), .O(n19326[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4980_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5014_5 (.CI(n48605), .I0(n19973[2]), .I1(n332), .CO(n48606));
    SB_LUT4 add_5014_4_lut (.I0(GND_net), .I1(n19973[1]), .I2(n259), .I3(n48604), 
            .O(n19756[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5014_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4980_3 (.CI(n49098), .I0(n19612[0]), .I1(n180_adj_4583), 
            .CO(n49099));
    SB_LUT4 add_4980_2_lut (.I0(GND_net), .I1(n38_adj_4584), .I2(n107_adj_4585), 
            .I3(GND_net), .O(n19326[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4980_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4980_2 (.CI(GND_net), .I0(n38_adj_4584), .I1(n107_adj_4585), 
            .CO(n49098));
    SB_LUT4 i48597_3_lut (.I0(n6_adj_4586), .I1(n535[10]), .I2(n21_adj_4551), 
            .I3(GND_net), .O(n65659));   // verilog/motorControl.v(47[25:43])
    defparam i48597_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4527_20 (.CI(n48880), .I0(n12488[17]), .I1(GND_net), 
            .CO(n48881));
    SB_CARRY add_5014_4 (.CI(n48604), .I0(n19973[1]), .I1(n259), .CO(n48605));
    SB_LUT4 add_4527_19_lut (.I0(GND_net), .I1(n12488[16]), .I2(GND_net), 
            .I3(n48879), .O(n10958[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46760_4_lut (.I0(n43_adj_4516), .I1(n25_adj_4521), .I2(n23_adj_4520), 
            .I3(n63900), .O(n63822));
    defparam i46760_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_5014_3_lut (.I0(GND_net), .I1(n19973[0]), .I2(n186), .I3(n48603), 
            .O(n19756[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5014_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_19 (.CI(n48879), .I0(n12488[16]), .I1(GND_net), 
            .CO(n48880));
    SB_CARRY add_5014_3 (.CI(n48603), .I0(n19973[0]), .I1(n186), .CO(n48604));
    SB_LUT4 add_4527_18_lut (.I0(GND_net), .I1(n12488[15]), .I2(GND_net), 
            .I3(n48878), .O(n10958[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5014_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n19756[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5014_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48412_4_lut (.I0(n24_adj_4566), .I1(n8_adj_4563), .I2(n45_adj_4515), 
            .I3(n63818), .O(n65474));   // verilog/motorControl.v(58[23:46])
    defparam i48412_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_5014_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n48603));
    SB_CARRY add_4527_18 (.CI(n48878), .I0(n12488[15]), .I1(GND_net), 
            .CO(n48879));
    SB_LUT4 i47280_3_lut (.I0(n65644), .I1(n285[12]), .I2(n25_adj_4521), 
            .I3(GND_net), .O(n64342));   // verilog/motorControl.v(58[23:46])
    defparam i47280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i106_2_lut (.I0(\Ki[2] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i155_2_lut (.I0(\Ki[3] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46625_4_lut (.I0(n455[13]), .I1(n67230), .I2(n28[13]), .I3(n65673), 
            .O(n63687));
    defparam i46625_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 LessThan_28_i29_rep_72_2_lut (.I0(n455[14]), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n67218));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i29_rep_72_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48171_4_lut (.I0(n455[15]), .I1(n67218), .I2(n28[15]), .I3(n63687), 
            .O(n65233));
    defparam i48171_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 LessThan_28_i33_rep_101_2_lut (.I0(n455[16]), .I1(n28[16]), 
            .I2(GND_net), .I3(GND_net), .O(n67247));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i33_rep_101_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4527_17_lut (.I0(GND_net), .I1(n12488[14]), .I2(GND_net), 
            .I3(n48877), .O(n10958[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_17 (.CI(n48877), .I0(n12488[14]), .I1(GND_net), 
            .CO(n48878));
    SB_LUT4 LessThan_19_i4_4_lut (.I0(n233[0]), .I1(n285[1]), .I2(n233[1]), 
            .I3(n285[0]), .O(n4_adj_4587));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 add_4527_16_lut (.I0(GND_net), .I1(n12488[13]), .I2(n1099_adj_4588), 
            .I3(n48876), .O(n10958[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48827_4_lut (.I0(n455[17]), .I1(n67247), .I2(n28[17]), .I3(n65233), 
            .O(n65889));
    defparam i48827_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i48598_3_lut (.I0(n65659), .I1(n535[11]), .I2(n23_adj_4565), 
            .I3(GND_net), .O(n65660));   // verilog/motorControl.v(47[25:43])
    defparam i48598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_28_i37_rep_63_2_lut (.I0(n455[18]), .I1(n28[18]), .I2(GND_net), 
            .I3(GND_net), .O(n67209));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i37_rep_63_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4527_16 (.CI(n48876), .I0(n12488[13]), .I1(n1099_adj_4588), 
            .CO(n48877));
    SB_LUT4 i48579_3_lut (.I0(n4_adj_4587), .I1(n285[13]), .I2(n27_adj_4527), 
            .I3(GND_net), .O(n65641));   // verilog/motorControl.v(58[23:46])
    defparam i48579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49092_4_lut (.I0(n455[19]), .I1(n67209), .I2(n28[19]), .I3(n65889), 
            .O(n66154));
    defparam i49092_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 add_4527_15_lut (.I0(GND_net), .I1(n12488[12]), .I2(n1026_adj_4591), 
            .I3(n48875), .O(n10958[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i106_2_lut (.I0(\Kp[2] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4592));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i106_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4527_15 (.CI(n48875), .I0(n12488[12]), .I1(n1026_adj_4591), 
            .CO(n48876));
    SB_LUT4 add_4527_14_lut (.I0(GND_net), .I1(n12488[11]), .I2(n953_adj_4593), 
            .I3(n48874), .O(n10958[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48580_3_lut (.I0(n65641), .I1(n285[14]), .I2(n29_adj_4518), 
            .I3(GND_net), .O(n65642));   // verilog/motorControl.v(58[23:46])
    defparam i48580_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4527_14 (.CI(n48874), .I0(n12488[11]), .I1(n953_adj_4593), 
            .CO(n48875));
    SB_LUT4 add_4527_13_lut (.I0(GND_net), .I1(n12488[10]), .I2(n880_adj_4594), 
            .I3(n48873), .O(n10958[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5082_7_lut (.I0(GND_net), .I1(n57914), .I2(n490_adj_4595), 
            .I3(n48596), .O(n20432[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5082_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46814_4_lut (.I0(n33_adj_4523), .I1(n31_adj_4519), .I2(n29_adj_4518), 
            .I3(n63886), .O(n63876));
    defparam i46814_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48905_4_lut (.I0(n30_adj_4535), .I1(n10_adj_4534), .I2(n35_adj_4522), 
            .I3(n63872), .O(n65967));   // verilog/motorControl.v(58[23:46])
    defparam i48905_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_24_i204_2_lut (.I0(\Ki[4] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4596));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i204_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4527_13 (.CI(n48873), .I0(n12488[10]), .I1(n880_adj_4594), 
            .CO(n48874));
    SB_LUT4 add_5082_6_lut (.I0(GND_net), .I1(n20502[3]), .I2(n417), .I3(n48595), 
            .O(n20432[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5082_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_28_i41_rep_60_2_lut (.I0(n455[20]), .I1(n28[20]), .I2(GND_net), 
            .I3(GND_net), .O(n67206));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i41_rep_60_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n9972_bdd_4_lut_49641 (.I0(n9972), .I1(n63117), .I2(setpoint[21]), 
            .I3(n4744), .O(n66735));
    defparam n9972_bdd_4_lut_49641.LUT_INIT = 16'he4aa;
    SB_CARRY add_5082_6 (.CI(n48595), .I0(n20502[3]), .I1(n417), .CO(n48596));
    SB_LUT4 LessThan_11_i8_3_lut (.I0(n535[4]), .I1(n535[8]), .I2(n17_adj_4553), 
            .I3(GND_net), .O(n8_adj_4597));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46721_4_lut (.I0(n27_adj_4598), .I1(n15_adj_4599), .I2(n13_adj_4600), 
            .I3(n11_adj_4601), .O(n63783));
    defparam i46721_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_i155_2_lut (.I0(\Kp[3] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4602));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4527_12_lut (.I0(GND_net), .I1(n12488[9]), .I2(n807_adj_4603), 
            .I3(n48872), .O(n10958[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_12 (.CI(n48872), .I0(n12488[9]), .I1(n807_adj_4603), 
            .CO(n48873));
    SB_LUT4 i47282_3_lut (.I0(n65642), .I1(n285[15]), .I2(n31_adj_4519), 
            .I3(GND_net), .O(n64344));   // verilog/motorControl.v(58[23:46])
    defparam i47282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i394_2_lut (.I0(\Kp[8] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n585_adj_4604));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5082_5_lut (.I0(GND_net), .I1(n20502[2]), .I2(n344_adj_4605), 
            .I3(n48594), .O(n20432[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5082_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i253_2_lut (.I0(\Ki[5] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i253_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5082_5 (.CI(n48594), .I0(n20502[2]), .I1(n344_adj_4605), 
            .CO(n48595));
    SB_LUT4 i49116_4_lut (.I0(n64344), .I1(n65967), .I2(n35_adj_4522), 
            .I3(n63876), .O(n66178));   // verilog/motorControl.v(58[23:46])
    defparam i49116_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_5082_4_lut (.I0(GND_net), .I1(n20502[1]), .I2(n271), .I3(n48593), 
            .O(n20432[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5082_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49117_3_lut (.I0(n66178), .I1(n285[18]), .I2(n37_adj_4517), 
            .I3(GND_net), .O(n66179));   // verilog/motorControl.v(58[23:46])
    defparam i49117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_i443_2_lut (.I0(\Kp[9] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_4606));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i492_2_lut (.I0(\Kp[10] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4607));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4527_11_lut (.I0(GND_net), .I1(n12488[8]), .I2(n734_adj_4608), 
            .I3(n48871), .O(n10958[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_11 (.CI(n48871), .I0(n12488[8]), .I1(n734_adj_4608), 
            .CO(n48872));
    SB_CARRY add_5082_4 (.CI(n48593), .I0(n20502[1]), .I1(n271), .CO(n48594));
    SB_LUT4 add_5082_3_lut (.I0(GND_net), .I1(n20502[0]), .I2(n198), .I3(n48592), 
            .O(n20432[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5082_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4527_10_lut (.I0(GND_net), .I1(n12488[7]), .I2(n661_adj_4609), 
            .I3(n48870), .O(n10958[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5082_3 (.CI(n48592), .I0(n20502[0]), .I1(n198), .CO(n48593));
    SB_LUT4 n66735_bdd_4_lut (.I0(n66735), .I1(n535[21]), .I2(n455[21]), 
            .I3(n4744), .O(n66738));
    defparam n66735_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i49085_3_lut (.I0(n66179), .I1(n285[19]), .I2(n39_adj_4514), 
            .I3(GND_net), .O(n66147));   // verilog/motorControl.v(58[23:46])
    defparam i49085_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46764_4_lut (.I0(n43_adj_4516), .I1(n41_adj_4513), .I2(n39_adj_4514), 
            .I3(n66080), .O(n63826));
    defparam i46764_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_26_i12_3_lut (.I0(n455[7]), .I1(n455[16]), .I2(n33), 
            .I3(GND_net), .O(n12_adj_4610));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i302_2_lut (.I0(\Ki[6] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4611));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_11_i24_3_lut (.I0(n16_adj_4577), .I1(n535[22]), .I2(n45_adj_4537), 
            .I3(GND_net), .O(n24_adj_4612));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n9972_bdd_4_lut_49636 (.I0(n9972), .I1(n63116), .I2(setpoint[20]), 
            .I3(n4744), .O(n66729));
    defparam n9972_bdd_4_lut_49636.LUT_INIT = 16'he4aa;
    SB_LUT4 n66729_bdd_4_lut (.I0(n66729), .I1(n535[20]), .I2(n455[20]), 
            .I3(n4744), .O(n66732));
    defparam n66729_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n9972_bdd_4_lut_49631 (.I0(n9972), .I1(n63115), .I2(setpoint[19]), 
            .I3(n4744), .O(n66723));
    defparam n9972_bdd_4_lut_49631.LUT_INIT = 16'he4aa;
    SB_LUT4 n66723_bdd_4_lut (.I0(n66723), .I1(n535[19]), .I2(n455[19]), 
            .I3(n4744), .O(n66726));
    defparam n66723_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_26_i10_3_lut (.I0(n455[5]), .I1(n455[6]), .I2(n13_adj_4600), 
            .I3(GND_net), .O(n10_adj_4613));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_add_1221_24_lut (.I0(n207[23]), .I1(n11500[21]), .I2(GND_net), 
            .I3(n49492), .O(n11041[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_23_add_1221_23_lut (.I0(GND_net), .I1(n11500[20]), .I2(GND_net), 
            .I3(n49491), .O(n360[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_23 (.CI(n49491), .I0(n11500[20]), .I1(GND_net), 
            .CO(n49492));
    SB_LUT4 LessThan_26_i30_3_lut (.I0(n12_adj_4610), .I1(n455[17]), .I2(n35), 
            .I3(GND_net), .O(n30_adj_4614));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_add_1221_22_lut (.I0(GND_net), .I1(n11500[19]), .I2(GND_net), 
            .I3(n49490), .O(n360[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_22 (.CI(n49490), .I0(n11500[19]), .I1(GND_net), 
            .CO(n49491));
    SB_LUT4 mult_23_add_1221_21_lut (.I0(GND_net), .I1(n11500[18]), .I2(GND_net), 
            .I3(n49489), .O(n360[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_21 (.CI(n49489), .I0(n11500[18]), .I1(GND_net), 
            .CO(n49490));
    SB_CARRY add_4527_10 (.CI(n48870), .I0(n12488[7]), .I1(n661_adj_4609), 
            .CO(n48871));
    SB_LUT4 mult_23_add_1221_20_lut (.I0(GND_net), .I1(n11500[17]), .I2(GND_net), 
            .I3(n49488), .O(n360[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_20 (.CI(n49488), .I0(n11500[17]), .I1(GND_net), 
            .CO(n49489));
    SB_LUT4 mult_23_add_1221_19_lut (.I0(GND_net), .I1(n11500[16]), .I2(GND_net), 
            .I3(n49487), .O(n360[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_19 (.CI(n49487), .I0(n11500[16]), .I1(GND_net), 
            .CO(n49488));
    SB_LUT4 mult_23_add_1221_18_lut (.I0(GND_net), .I1(n11500[15]), .I2(GND_net), 
            .I3(n49486), .O(n360[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_18 (.CI(n49486), .I0(n11500[15]), .I1(GND_net), 
            .CO(n49487));
    SB_LUT4 i46990_4_lut (.I0(n43_adj_4541), .I1(n25_adj_4564), .I2(n23_adj_4565), 
            .I3(n64127), .O(n64052));
    defparam i46990_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_add_1221_17_lut (.I0(GND_net), .I1(n11500[14]), .I2(GND_net), 
            .I3(n49485), .O(n360[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i204_2_lut (.I0(\Kp[4] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4615));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i204_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_23_add_1221_17 (.CI(n49485), .I0(n11500[14]), .I1(GND_net), 
            .CO(n49486));
    SB_LUT4 mult_23_add_1221_16_lut (.I0(GND_net), .I1(n11500[13]), .I2(n1096_adj_4616), 
            .I3(n49484), .O(n360[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_16 (.CI(n49484), .I0(n11500[13]), .I1(n1096_adj_4616), 
            .CO(n49485));
    SB_LUT4 mult_23_add_1221_15_lut (.I0(GND_net), .I1(n11500[12]), .I2(n1023_adj_4617), 
            .I3(n49483), .O(n360[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_15 (.CI(n49483), .I0(n11500[12]), .I1(n1023_adj_4617), 
            .CO(n49484));
    SB_LUT4 mult_23_add_1221_14_lut (.I0(GND_net), .I1(n11500[11]), .I2(n950_adj_4618), 
            .I3(n49482), .O(n360[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_14 (.CI(n49482), .I0(n11500[11]), .I1(n950_adj_4618), 
            .CO(n49483));
    SB_LUT4 mult_23_add_1221_13_lut (.I0(GND_net), .I1(n11500[10]), .I2(n877_adj_4619), 
            .I3(n49481), .O(n360[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48963_4_lut (.I0(n64342), .I1(n65474), .I2(n45_adj_4515), 
            .I3(n63822), .O(n66025));   // verilog/motorControl.v(58[23:46])
    defparam i48963_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY mult_23_add_1221_13 (.CI(n49481), .I0(n11500[10]), .I1(n877_adj_4619), 
            .CO(n49482));
    SB_LUT4 add_5082_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n20432[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5082_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_add_1221_12_lut (.I0(GND_net), .I1(n11500[9]), .I2(n804_adj_4621), 
            .I3(n49480), .O(n360[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_12 (.CI(n49480), .I0(n11500[9]), .I1(n804_adj_4621), 
            .CO(n49481));
    SB_LUT4 mult_23_add_1221_11_lut (.I0(GND_net), .I1(n11500[8]), .I2(n731_adj_4607), 
            .I3(n49479), .O(n360[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5082_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n48592));
    SB_CARRY mult_23_add_1221_11 (.CI(n49479), .I0(n11500[8]), .I1(n731_adj_4607), 
            .CO(n49480));
    SB_LUT4 mult_23_add_1221_10_lut (.I0(GND_net), .I1(n11500[7]), .I2(n658_adj_4606), 
            .I3(n49478), .O(n360[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_10 (.CI(n49478), .I0(n11500[7]), .I1(n658_adj_4606), 
            .CO(n49479));
    SB_LUT4 mult_23_add_1221_9_lut (.I0(GND_net), .I1(n11500[6]), .I2(n585_adj_4604), 
            .I3(n49477), .O(n360[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_9 (.CI(n49477), .I0(n11500[6]), .I1(n585_adj_4604), 
            .CO(n49478));
    SB_LUT4 mult_23_add_1221_8_lut (.I0(GND_net), .I1(n11500[5]), .I2(n512_adj_4578), 
            .I3(n49476), .O(n360[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_8 (.CI(n49476), .I0(n11500[5]), .I1(n512_adj_4578), 
            .CO(n49477));
    SB_LUT4 i47288_3_lut (.I0(n66147), .I1(n285[20]), .I2(n41_adj_4513), 
            .I3(GND_net), .O(n64350));   // verilog/motorControl.v(58[23:46])
    defparam i47288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_23_add_1221_7_lut (.I0(GND_net), .I1(n11500[4]), .I2(n439_adj_4510), 
            .I3(n49475), .O(n360[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47708_4_lut (.I0(n13_adj_4600), .I1(n11_adj_4601), .I2(n9_adj_4623), 
            .I3(n63814), .O(n64770));
    defparam i47708_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY mult_23_add_1221_7 (.CI(n49475), .I0(n11500[4]), .I1(n439_adj_4510), 
            .CO(n49476));
    SB_LUT4 i47702_4_lut (.I0(n19_adj_4624), .I1(n17_adj_4625), .I2(n15_adj_4599), 
            .I3(n64770), .O(n64764));
    defparam i47702_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 n9972_bdd_4_lut_49626 (.I0(n9972), .I1(n63114), .I2(setpoint[18]), 
            .I3(n4744), .O(n66705));
    defparam n9972_bdd_4_lut_49626.LUT_INIT = 16'he4aa;
    SB_LUT4 n66705_bdd_4_lut (.I0(n66705), .I1(n535[18]), .I2(n455[18]), 
            .I3(n4744), .O(n66708));
    defparam n66705_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i48851_4_lut (.I0(n25_adj_4626), .I1(n23_adj_4627), .I2(n21_adj_4628), 
            .I3(n64764), .O(n65913));
    defparam i48851_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48215_4_lut (.I0(n31), .I1(n29), .I2(n27_adj_4598), .I3(n65913), 
            .O(n65277));
    defparam i48215_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_23_add_1221_6_lut (.I0(GND_net), .I1(n11500[3]), .I2(n366), 
            .I3(n49474), .O(n360[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_6 (.CI(n49474), .I0(n11500[3]), .I1(n366), 
            .CO(n49475));
    SB_LUT4 mult_23_add_1221_5_lut (.I0(GND_net), .I1(n11500[2]), .I2(n293_adj_4477), 
            .I3(n49473), .O(n360[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_5 (.CI(n49473), .I0(n11500[2]), .I1(n293_adj_4477), 
            .CO(n49474));
    SB_LUT4 i48408_4_lut (.I0(n24_adj_4612), .I1(n8_adj_4597), .I2(n45_adj_4537), 
            .I3(n64046), .O(n65470));   // verilog/motorControl.v(47[25:43])
    defparam i48408_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_23_add_1221_4_lut (.I0(GND_net), .I1(n11500[1]), .I2(n220_adj_4476), 
            .I3(n49472), .O(n360[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_4 (.CI(n49472), .I0(n11500[1]), .I1(n220_adj_4476), 
            .CO(n49473));
    SB_LUT4 mult_23_add_1221_3_lut (.I0(GND_net), .I1(n11500[0]), .I2(n147_adj_4475), 
            .I3(n49471), .O(n360[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_3 (.CI(n49471), .I0(n11500[0]), .I1(n147_adj_4475), 
            .CO(n49472));
    SB_LUT4 mult_23_add_1221_2_lut (.I0(GND_net), .I1(n5_adj_4465), .I2(n74_adj_4464), 
            .I3(GND_net), .O(n360[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_23_add_1221_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_23_add_1221_2 (.CI(GND_net), .I0(n5_adj_4465), .I1(n74_adj_4464), 
            .CO(n49471));
    SB_LUT4 add_4527_9_lut (.I0(GND_net), .I1(n12488[6]), .I2(n588_adj_4463), 
            .I3(n48869), .O(n10958[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_9 (.CI(n48869), .I0(n12488[6]), .I1(n588_adj_4463), 
            .CO(n48870));
    SB_LUT4 i48965_4_lut (.I0(n64350), .I1(n66025), .I2(n45_adj_4515), 
            .I3(n63826), .O(n66027));   // verilog/motorControl.v(58[23:46])
    defparam i48965_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i46484_3_lut_4_lut (.I0(n455[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(n455[2]), .O(n63546));   // verilog/motorControl.v(65[25:41])
    defparam i46484_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_5033_10_lut (.I0(GND_net), .I1(n20150[7]), .I2(n700), 
            .I3(n48591), .O(n19973[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5033_9_lut (.I0(GND_net), .I1(n20150[6]), .I2(n627), .I3(n48590), 
            .O(n19973[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i49012_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n65277), 
            .O(n66074));
    defparam i49012_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_23_i541_2_lut (.I0(\Kp[11] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_4621));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4552_23_lut (.I0(GND_net), .I1(n12999[20]), .I2(GND_net), 
            .I3(n49470), .O(n11500[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48966_3_lut (.I0(n66027), .I1(n233[23]), .I2(n285[23]), .I3(GND_net), 
            .O(n284));   // verilog/motorControl.v(58[23:46])
    defparam i48966_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_21_i11_3_lut (.I0(n233[10]), .I1(n285[10]), .I2(n284), 
            .I3(GND_net), .O(n310[10]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i11_3_lut (.I0(n310[10]), .I1(IntegralLimit[10]), .I2(n258), 
            .I3(GND_net), .O(n335[10]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4552_22_lut (.I0(GND_net), .I1(n12999[19]), .I2(GND_net), 
            .I3(n49469), .O(n11500[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4527_8_lut (.I0(GND_net), .I1(n12488[5]), .I2(n515_adj_4462), 
            .I3(n48868), .O(n10958[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47260_3_lut (.I0(n65660), .I1(n535[12]), .I2(n25_adj_4564), 
            .I3(GND_net), .O(n64322));   // verilog/motorControl.v(47[25:43])
    defparam i47260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i4_4_lut (.I0(setpoint[0]), .I1(n535[1]), .I2(setpoint[1]), 
            .I3(n535[0]), .O(n4_adj_4631));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i48595_3_lut (.I0(n4_adj_4631), .I1(n535[13]), .I2(n27_adj_4556), 
            .I3(GND_net), .O(n65657));   // verilog/motorControl.v(47[25:43])
    defparam i48595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48596_3_lut (.I0(n65657), .I1(n535[14]), .I2(n29_adj_4543), 
            .I3(GND_net), .O(n65658));   // verilog/motorControl.v(47[25:43])
    defparam i48596_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5033_9 (.CI(n48590), .I0(n20150[6]), .I1(n627), .CO(n48591));
    SB_LUT4 i47027_4_lut (.I0(n33_adj_4545), .I1(n31_adj_4544), .I2(n29_adj_4543), 
            .I3(n64108), .O(n64089));
    defparam i47027_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_i85_2_lut (.I0(\Kp[1] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n125));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5033_8_lut (.I0(GND_net), .I1(n20150[5]), .I2(n554_adj_4461), 
            .I3(n48589), .O(n19973[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48901_4_lut (.I0(n30_adj_4562), .I1(n10_adj_4561), .I2(n35_adj_4548), 
            .I3(n64076), .O(n65963));   // verilog/motorControl.v(47[25:43])
    defparam i48901_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_23_i38_2_lut (.I0(\Kp[0] ), .I1(n207[22]), .I2(GND_net), 
            .I3(GND_net), .O(n56));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_32_i6_3_lut_3_lut (.I0(n455[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(GND_net), .O(n6_adj_4632));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_CARRY add_4552_22 (.CI(n49469), .I0(n12999[19]), .I1(GND_net), 
            .CO(n49470));
    SB_LUT4 add_4552_21_lut (.I0(GND_net), .I1(n12999[18]), .I2(GND_net), 
            .I3(n49468), .O(n11500[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47262_3_lut (.I0(n65658), .I1(n535[15]), .I2(n31_adj_4544), 
            .I3(GND_net), .O(n64324));   // verilog/motorControl.v(47[25:43])
    defparam i47262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49112_4_lut (.I0(n64324), .I1(n65963), .I2(n35_adj_4548), 
            .I3(n64089), .O(n66174));   // verilog/motorControl.v(47[25:43])
    defparam i49112_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49113_3_lut (.I0(n66174), .I1(n535[18]), .I2(n37_adj_4538), 
            .I3(GND_net), .O(n66175));   // verilog/motorControl.v(47[25:43])
    defparam i49113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49091_3_lut (.I0(n66175), .I1(n535[19]), .I2(n39_adj_4546), 
            .I3(GND_net), .O(n66153));   // verilog/motorControl.v(47[25:43])
    defparam i49091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46994_4_lut (.I0(n43_adj_4541), .I1(n41_adj_4540), .I2(n39_adj_4546), 
            .I3(n66088), .O(n64056));
    defparam i46994_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48955_4_lut (.I0(n64322), .I1(n65470), .I2(n45_adj_4537), 
            .I3(n64052), .O(n66017));   // verilog/motorControl.v(47[25:43])
    defparam i48955_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_4552_21 (.CI(n49468), .I0(n12999[18]), .I1(GND_net), 
            .CO(n49469));
    SB_LUT4 add_4552_20_lut (.I0(GND_net), .I1(n12999[17]), .I2(GND_net), 
            .I3(n49467), .O(n11500[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i47268_3_lut (.I0(n66153), .I1(n535[20]), .I2(n41_adj_4540), 
            .I3(GND_net), .O(n64330));   // verilog/motorControl.v(47[25:43])
    defparam i47268_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4527_8 (.CI(n48868), .I0(n12488[5]), .I1(n515_adj_4462), 
            .CO(n48869));
    SB_LUT4 i48957_4_lut (.I0(n64330), .I1(n66017), .I2(n45_adj_4537), 
            .I3(n64056), .O(n66019));   // verilog/motorControl.v(47[25:43])
    defparam i48957_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_32_i37_2_lut (.I0(n455[18]), .I1(n535[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4633));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5033_8 (.CI(n48589), .I0(n20150[5]), .I1(n554_adj_4461), 
            .CO(n48590));
    SB_LUT4 LessThan_32_i45_2_lut (.I0(n455[22]), .I1(n535[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4634));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i41_2_lut (.I0(n455[20]), .I1(n535[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4635));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47115_3_lut_4_lut (.I0(setpoint[3]), .I1(n535[3]), .I2(n535[2]), 
            .I3(setpoint[2]), .O(n64177));   // verilog/motorControl.v(47[25:43])
    defparam i47115_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_4552_20 (.CI(n49467), .I0(n12999[17]), .I1(GND_net), 
            .CO(n49468));
    SB_LUT4 add_4552_19_lut (.I0(GND_net), .I1(n12999[16]), .I2(GND_net), 
            .I3(n49466), .O(n11500[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_32_i43_2_lut (.I0(n455[21]), .I1(n535[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4636));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i35_2_lut (.I0(n455[17]), .I1(n535[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4637));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i16_3_lut (.I0(n455[9]), .I1(n455[21]), .I2(n43), 
            .I3(GND_net), .O(n16_adj_4638));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_11_i6_3_lut_3_lut (.I0(setpoint[3]), .I1(n535[3]), 
            .I2(n535[2]), .I3(GND_net), .O(n6_adj_4586));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_CARRY add_4552_19 (.CI(n49466), .I0(n12999[16]), .I1(GND_net), 
            .CO(n49467));
    SB_LUT4 add_4552_18_lut (.I0(GND_net), .I1(n12999[15]), .I2(GND_net), 
            .I3(n49465), .O(n11500[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5033_7_lut (.I0(GND_net), .I1(n20150[4]), .I2(n481), .I3(n48588), 
            .O(n19973[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5033_7 (.CI(n48588), .I0(n20150[4]), .I1(n481), .CO(n48589));
    SB_LUT4 mult_24_i365_2_lut (.I0(\Ki[7] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i590_2_lut (.I0(\Kp[12] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_4619));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46582_3_lut_4_lut (.I0(PWMLimit[3]), .I1(n455[3]), .I2(n455[2]), 
            .I3(PWMLimit[2]), .O(n63644));   // verilog/motorControl.v(63[16:31])
    defparam i46582_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 n9972_bdd_4_lut_49611 (.I0(n9972), .I1(n63111), .I2(setpoint[17]), 
            .I3(n4744), .O(n66687));
    defparam n9972_bdd_4_lut_49611.LUT_INIT = 16'he4aa;
    SB_CARRY add_4552_18 (.CI(n49465), .I0(n12999[15]), .I1(GND_net), 
            .CO(n49466));
    SB_LUT4 mult_23_i608_2_lut (.I0(\Kp[12] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4552_17_lut (.I0(GND_net), .I1(n12999[14]), .I2(GND_net), 
            .I3(n49464), .O(n11500[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_32_i39_2_lut (.I0(n455[19]), .I1(n535[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4639));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4552_17 (.CI(n49464), .I0(n12999[14]), .I1(GND_net), 
            .CO(n49465));
    SB_LUT4 LessThan_32_i31_2_lut (.I0(n455[15]), .I1(n535[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4640));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_24_i351_2_lut (.I0(\Ki[7] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_30_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(n455[3]), 
            .I2(n455[2]), .I3(GND_net), .O(n6));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 LessThan_32_i33_2_lut (.I0(n455[16]), .I1(n535[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4641));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i27_2_lut (.I0(n455[13]), .I1(n535[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4642));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i29_2_lut (.I0(n455[14]), .I1(n535[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4643));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(n7062), .I1(n7064), .I2(n24983), .I3(n38638), 
            .O(n4744));
    defparam i3_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 add_4552_16_lut (.I0(GND_net), .I1(n12999[13]), .I2(n1099), 
            .I3(n49463), .O(n11500[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4552_16 (.CI(n49463), .I0(n12999[13]), .I1(n1099), .CO(n49464));
    SB_LUT4 add_4527_7_lut (.I0(GND_net), .I1(n12488[4]), .I2(n442_adj_4443), 
            .I3(n48867), .O(n10958[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_24_i400_2_lut (.I0(\Ki[8] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5033_6_lut (.I0(GND_net), .I1(n20150[3]), .I2(n408), .I3(n48587), 
            .O(n19973[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5033_6 (.CI(n48587), .I0(n20150[3]), .I1(n408), .CO(n48588));
    SB_LUT4 i46752_3_lut_4_lut (.I0(deadband[3]), .I1(n455[3]), .I2(n455[2]), 
            .I3(deadband[2]), .O(n63814));   // verilog/motorControl.v(62[14:31])
    defparam i46752_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_4552_15_lut (.I0(GND_net), .I1(n12999[12]), .I2(n1026), 
            .I3(n49462), .O(n11500[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4552_15 (.CI(n49462), .I0(n12999[12]), .I1(n1026), .CO(n49463));
    SB_LUT4 add_4552_14_lut (.I0(GND_net), .I1(n12999[11]), .I2(n953), 
            .I3(n49461), .O(n11500[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4552_14 (.CI(n49461), .I0(n12999[11]), .I1(n953), .CO(n49462));
    SB_LUT4 add_4552_13_lut (.I0(GND_net), .I1(n12999[10]), .I2(n880), 
            .I3(n49460), .O(n11500[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4552_13 (.CI(n49460), .I0(n12999[10]), .I1(n880), .CO(n49461));
    SB_LUT4 LessThan_26_i6_3_lut_3_lut (.I0(deadband[3]), .I1(n455[3]), 
            .I2(n455[2]), .I3(GND_net), .O(n6_adj_4644));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 add_4552_12_lut (.I0(GND_net), .I1(n12999[9]), .I2(n807), 
            .I3(n49459), .O(n11500[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4552_12 (.CI(n49459), .I0(n12999[9]), .I1(n807), .CO(n49460));
    SB_LUT4 add_4552_11_lut (.I0(GND_net), .I1(n12999[8]), .I2(n734), 
            .I3(n49458), .O(n11500[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4552_11 (.CI(n49458), .I0(n12999[8]), .I1(n734), .CO(n49459));
    SB_LUT4 add_4552_10_lut (.I0(GND_net), .I1(n12999[7]), .I2(n661), 
            .I3(n49457), .O(n11500[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4552_10 (.CI(n49457), .I0(n12999[7]), .I1(n661), .CO(n49458));
    SB_LUT4 add_4552_9_lut (.I0(GND_net), .I1(n12999[6]), .I2(n588), .I3(n49456), 
            .O(n11500[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4552_9 (.CI(n49456), .I0(n12999[6]), .I1(n588), .CO(n49457));
    SB_LUT4 add_4552_8_lut (.I0(GND_net), .I1(n12999[5]), .I2(n515), .I3(n49455), 
            .O(n11500[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4552_8 (.CI(n49455), .I0(n12999[5]), .I1(n515), .CO(n49456));
    SB_LUT4 add_4552_7_lut (.I0(GND_net), .I1(n12999[4]), .I2(n442), .I3(n49454), 
            .O(n11500[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4552_7 (.CI(n49454), .I0(n12999[4]), .I1(n442), .CO(n49455));
    SB_LUT4 add_4552_6_lut (.I0(GND_net), .I1(n12999[3]), .I2(n369_adj_4439), 
            .I3(n49453), .O(n11500[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4552_6 (.CI(n49453), .I0(n12999[3]), .I1(n369_adj_4439), 
            .CO(n49454));
    SB_LUT4 add_4552_5_lut (.I0(GND_net), .I1(n12999[2]), .I2(n296_adj_4437), 
            .I3(n49452), .O(n11500[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4552_5 (.CI(n49452), .I0(n12999[2]), .I1(n296_adj_4437), 
            .CO(n49453));
    SB_LUT4 mult_23_i253_2_lut (.I0(\Kp[5] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4645));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i253_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4527_7 (.CI(n48867), .I0(n12488[4]), .I1(n442_adj_4443), 
            .CO(n48868));
    SB_LUT4 add_4552_4_lut (.I0(GND_net), .I1(n12999[1]), .I2(n223_adj_4436), 
            .I3(n49451), .O(n11500[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4552_4 (.CI(n49451), .I0(n12999[1]), .I1(n223_adj_4436), 
            .CO(n49452));
    SB_LUT4 mult_24_i449_2_lut (.I0(\Ki[9] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4552_3_lut (.I0(GND_net), .I1(n12999[0]), .I2(n150_adj_4435), 
            .I3(n49450), .O(n11500[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4527_6_lut (.I0(GND_net), .I1(n12488[3]), .I2(n369), .I3(n48866), 
            .O(n10958[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_6 (.CI(n48866), .I0(n12488[3]), .I1(n369), .CO(n48867));
    SB_CARRY add_4552_3 (.CI(n49450), .I0(n12999[0]), .I1(n150_adj_4435), 
            .CO(n49451));
    SB_LUT4 add_4527_5_lut (.I0(GND_net), .I1(n12488[2]), .I2(n296), .I3(n48865), 
            .O(n10958[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5033_5_lut (.I0(GND_net), .I1(n20150[2]), .I2(n335_c), 
            .I3(n48586), .O(n19973[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_5 (.CI(n48865), .I0(n12488[2]), .I1(n296), .CO(n48866));
    SB_CARRY add_5033_5 (.CI(n48586), .I0(n20150[2]), .I1(n335_c), .CO(n48587));
    SB_LUT4 mult_23_i302_2_lut (.I0(\Kp[6] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4646));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4552_2_lut (.I0(GND_net), .I1(n8_adj_4434), .I2(n77), 
            .I3(GND_net), .O(n11500[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4552_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4527_4_lut (.I0(GND_net), .I1(n12488[1]), .I2(n223_adj_4433), 
            .I3(n48864), .O(n10958[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_4 (.CI(n48864), .I0(n12488[1]), .I1(n223_adj_4433), 
            .CO(n48865));
    SB_CARRY add_4552_2 (.CI(GND_net), .I0(n8_adj_4434), .I1(n77), .CO(n49450));
    SB_LUT4 add_4527_3_lut (.I0(GND_net), .I1(n12488[0]), .I2(n150), .I3(n48863), 
            .O(n10958[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5033_4_lut (.I0(GND_net), .I1(n20150[1]), .I2(n262), .I3(n48585), 
            .O(n19973[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_3 (.CI(n48863), .I0(n12488[0]), .I1(n150), .CO(n48864));
    SB_CARRY add_5033_4 (.CI(n48585), .I0(n20150[1]), .I1(n262), .CO(n48586));
    SB_LUT4 mult_23_i639_2_lut (.I0(\Kp[13] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n950_adj_4618));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4639_22_lut (.I0(GND_net), .I1(n14310[19]), .I2(GND_net), 
            .I3(n49449), .O(n12999[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4527_2_lut (.I0(GND_net), .I1(n8_adj_4647), .I2(n77_adj_4648), 
            .I3(GND_net), .O(n10958[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4527_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4639_21_lut (.I0(GND_net), .I1(n14310[18]), .I2(GND_net), 
            .I3(n49448), .O(n12999[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4639_21 (.CI(n49448), .I0(n14310[18]), .I1(GND_net), 
            .CO(n49449));
    SB_LUT4 add_5033_3_lut (.I0(GND_net), .I1(n20150[0]), .I2(n189), .I3(n48584), 
            .O(n19973[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4527_2 (.CI(GND_net), .I0(n8_adj_4647), .I1(n77_adj_4648), 
            .CO(n48863));
    SB_CARRY add_5033_3 (.CI(n48584), .I0(n20150[0]), .I1(n189), .CO(n48585));
    SB_LUT4 add_4616_22_lut (.I0(GND_net), .I1(n13844[19]), .I2(GND_net), 
            .I3(n48862), .O(n12488[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4639_20_lut (.I0(GND_net), .I1(n14310[17]), .I2(GND_net), 
            .I3(n49447), .O(n12999[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5033_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n19973[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5033_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4639_20 (.CI(n49447), .I0(n14310[17]), .I1(GND_net), 
            .CO(n49448));
    SB_LUT4 i46448_4_lut (.I0(n27_adj_4642), .I1(n15_adj_4649), .I2(n13_adj_4650), 
            .I3(n11_adj_4651), .O(n63510));
    defparam i46448_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_26_i8_3_lut (.I0(n455[4]), .I1(n455[8]), .I2(n17_adj_4625), 
            .I3(GND_net), .O(n8_adj_4652));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i12_3_lut (.I0(n535[7]), .I1(n535[16]), .I2(n33_adj_4641), 
            .I3(GND_net), .O(n12_adj_4653));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4639_19_lut (.I0(GND_net), .I1(n14310[16]), .I2(GND_net), 
            .I3(n49446), .O(n12999[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4616_21_lut (.I0(GND_net), .I1(n13844[18]), .I2(GND_net), 
            .I3(n48861), .O(n12488[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5033_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n48584));
    SB_CARRY add_4616_21 (.CI(n48861), .I0(n13844[18]), .I1(GND_net), 
            .CO(n48862));
    SB_CARRY add_4639_19 (.CI(n49446), .I0(n14310[16]), .I1(GND_net), 
            .CO(n49447));
    SB_LUT4 add_4616_20_lut (.I0(GND_net), .I1(n13844[17]), .I2(GND_net), 
            .I3(n48860), .O(n12488[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i657_2_lut (.I0(\Kp[13] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i657_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4616_20 (.CI(n48860), .I0(n13844[17]), .I1(GND_net), 
            .CO(n48861));
    SB_LUT4 add_4616_19_lut (.I0(GND_net), .I1(n13844[16]), .I2(GND_net), 
            .I3(n48859), .O(n12488[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4639_18_lut (.I0(GND_net), .I1(n14310[15]), .I2(GND_net), 
            .I3(n49445), .O(n12999[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4616_19 (.CI(n48859), .I0(n13844[16]), .I1(GND_net), 
            .CO(n48860));
    SB_LUT4 add_4616_18_lut (.I0(GND_net), .I1(n13844[15]), .I2(GND_net), 
            .I3(n48858), .O(n12488[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4639_18 (.CI(n49445), .I0(n14310[15]), .I1(GND_net), 
            .CO(n49446));
    SB_CARRY add_4616_18 (.CI(n48858), .I0(n13844[15]), .I1(GND_net), 
            .CO(n48859));
    SB_LUT4 add_4639_17_lut (.I0(GND_net), .I1(n14310[14]), .I2(GND_net), 
            .I3(n49444), .O(n12999[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4616_17_lut (.I0(GND_net), .I1(n13844[14]), .I2(GND_net), 
            .I3(n48857), .O(n12488[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_26_i24_3_lut (.I0(n16_adj_4638), .I1(n455[22]), .I2(n45_adj_4654), 
            .I3(GND_net), .O(n24_adj_4655));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4616_17 (.CI(n48857), .I0(n13844[14]), .I1(GND_net), 
            .CO(n48858));
    SB_LUT4 n66687_bdd_4_lut (.I0(n66687), .I1(n535[17]), .I2(n455[17]), 
            .I3(n4744), .O(n66690));
    defparam n66687_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_4639_17 (.CI(n49444), .I0(n14310[14]), .I1(GND_net), 
            .CO(n49445));
    SB_LUT4 add_4616_16_lut (.I0(GND_net), .I1(n13844[13]), .I2(n1102), 
            .I3(n48856), .O(n12488[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4639_16_lut (.I0(GND_net), .I1(n14310[13]), .I2(n1102_adj_4656), 
            .I3(n49443), .O(n12999[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4616_16 (.CI(n48856), .I0(n13844[13]), .I1(n1102), .CO(n48857));
    SB_LUT4 mult_23_i688_2_lut (.I0(\Kp[14] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1023_adj_4617));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_32_i10_3_lut (.I0(n535[5]), .I1(n535[6]), .I2(n13_adj_4650), 
            .I3(GND_net), .O(n10_adj_4657));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i30_3_lut (.I0(n12_adj_4653), .I1(n535[17]), .I2(n35_adj_4637), 
            .I3(GND_net), .O(n30_adj_4658));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47486_4_lut (.I0(n13_adj_4650), .I1(n11_adj_4651), .I2(n9_adj_4659), 
            .I3(n63546), .O(n64548));
    defparam i47486_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i47480_4_lut (.I0(n19_adj_4660), .I1(n17_adj_4661), .I2(n15_adj_4649), 
            .I3(n64548), .O(n64542));
    defparam i47480_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i48785_4_lut (.I0(n25_adj_4662), .I1(n23_adj_4663), .I2(n21_adj_4664), 
            .I3(n64542), .O(n65847));
    defparam i48785_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48087_4_lut (.I0(n31_adj_4640), .I1(n29_adj_4643), .I2(n27_adj_4642), 
            .I3(n65847), .O(n65149));
    defparam i48087_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48985_4_lut (.I0(n37_adj_4633), .I1(n35_adj_4637), .I2(n33_adj_4641), 
            .I3(n65149), .O(n66047));
    defparam i48985_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48117_3_lut (.I0(n6_adj_4632), .I1(n535[10]), .I2(n21_adj_4664), 
            .I3(GND_net), .O(n65179));   // verilog/motorControl.v(65[25:41])
    defparam i48117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48118_3_lut (.I0(n65179), .I1(n535[11]), .I2(n23_adj_4663), 
            .I3(GND_net), .O(n65180));   // verilog/motorControl.v(65[25:41])
    defparam i48118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i16_3_lut (.I0(n535[9]), .I1(n535[21]), .I2(n43_adj_4636), 
            .I3(GND_net), .O(n16_adj_4665));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4639_16 (.CI(n49443), .I0(n14310[13]), .I1(n1102_adj_4656), 
            .CO(n49444));
    SB_LUT4 add_4616_15_lut (.I0(GND_net), .I1(n13844[12]), .I2(n1029), 
            .I3(n48855), .O(n12488[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_15_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR counter_2045_2046__i1 (.Q(counter[0]), .C(clk16MHz), .D(n61[0]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_LUT4 mult_23_i737_2_lut (.I0(\Kp[15] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1096_adj_4616));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4639_15_lut (.I0(GND_net), .I1(n14310[12]), .I2(n1029_adj_4666), 
            .I3(n49442), .O(n12999[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4616_15 (.CI(n48855), .I0(n13844[12]), .I1(n1029), .CO(n48856));
    SB_LUT4 add_4616_14_lut (.I0(GND_net), .I1(n13844[11]), .I2(n956), 
            .I3(n48854), .O(n12488[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_14_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result_i0_i23 (.Q(duty[23]), .C(clk16MHz), .E(control_update), 
            .D(n66852), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_4639_15 (.CI(n49442), .I0(n14310[12]), .I1(n1029_adj_4666), 
            .CO(n49443));
    SB_CARRY add_4616_14 (.CI(n48854), .I0(n13844[11]), .I1(n956), .CO(n48855));
    SB_LUT4 add_4616_13_lut (.I0(GND_net), .I1(n13844[10]), .I2(n883), 
            .I3(n48853), .O(n12488[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4639_14_lut (.I0(GND_net), .I1(n14310[11]), .I2(n956_adj_4667), 
            .I3(n49441), .O(n12999[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4616_13 (.CI(n48853), .I0(n13844[10]), .I1(n883), .CO(n48854));
    SB_LUT4 add_4616_12_lut (.I0(GND_net), .I1(n13844[9]), .I2(n810), 
            .I3(n48852), .O(n12488[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4616_12 (.CI(n48852), .I0(n13844[9]), .I1(n810), .CO(n48853));
    SB_CARRY add_4639_14 (.CI(n49441), .I0(n14310[11]), .I1(n956_adj_4667), 
            .CO(n49442));
    SB_LUT4 add_4639_13_lut (.I0(GND_net), .I1(n14310[10]), .I2(n883_adj_4668), 
            .I3(n49440), .O(n12999[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4616_11_lut (.I0(GND_net), .I1(n13844[8]), .I2(n737), 
            .I3(n48851), .O(n12488[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4616_11 (.CI(n48851), .I0(n13844[8]), .I1(n737), .CO(n48852));
    SB_LUT4 add_4616_10_lut (.I0(GND_net), .I1(n13844[7]), .I2(n664), 
            .I3(n48850), .O(n12488[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4639_13 (.CI(n49440), .I0(n14310[10]), .I1(n883_adj_4668), 
            .CO(n49441));
    SB_LUT4 add_4639_12_lut (.I0(GND_net), .I1(n14310[9]), .I2(n810_adj_4669), 
            .I3(n49439), .O(n12999[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4616_10 (.CI(n48850), .I0(n13844[7]), .I1(n664), .CO(n48851));
    SB_LUT4 add_4616_9_lut (.I0(GND_net), .I1(n13844[6]), .I2(n591), .I3(n48849), 
            .O(n12488[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4639_12 (.CI(n49439), .I0(n14310[9]), .I1(n810_adj_4669), 
            .CO(n49440));
    SB_LUT4 add_4639_11_lut (.I0(GND_net), .I1(n14310[8]), .I2(n737_adj_4670), 
            .I3(n49438), .O(n12999[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4616_9 (.CI(n48849), .I0(n13844[6]), .I1(n591), .CO(n48850));
    SB_CARRY add_4639_11 (.CI(n49438), .I0(n14310[8]), .I1(n737_adj_4670), 
            .CO(n49439));
    SB_LUT4 add_4639_10_lut (.I0(GND_net), .I1(n14310[7]), .I2(n664_adj_4671), 
            .I3(n49437), .O(n12999[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48575_3_lut (.I0(n6_adj_4644), .I1(n455[10]), .I2(n21_adj_4628), 
            .I3(GND_net), .O(n65637));   // verilog/motorControl.v(62[14:31])
    defparam i48575_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4616_8_lut (.I0(GND_net), .I1(n13844[5]), .I2(n518), .I3(n48848), 
            .O(n12488[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4639_10 (.CI(n49437), .I0(n14310[7]), .I1(n664_adj_4671), 
            .CO(n49438));
    SB_CARRY add_4616_8 (.CI(n48848), .I0(n13844[5]), .I1(n518), .CO(n48849));
    SB_LUT4 add_4616_7_lut (.I0(GND_net), .I1(n13844[4]), .I2(n445_adj_4672), 
            .I3(n48847), .O(n12488[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4616_7 (.CI(n48847), .I0(n13844[4]), .I1(n445_adj_4672), 
            .CO(n48848));
    SB_LUT4 add_4616_6_lut (.I0(GND_net), .I1(n13844[3]), .I2(n372), .I3(n48846), 
            .O(n12488[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4639_9_lut (.I0(GND_net), .I1(n14310[6]), .I2(n591_adj_4673), 
            .I3(n49436), .O(n12999[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4639_9 (.CI(n49436), .I0(n14310[6]), .I1(n591_adj_4673), 
            .CO(n49437));
    SB_CARRY add_4616_6 (.CI(n48846), .I0(n13844[3]), .I1(n372), .CO(n48847));
    SB_LUT4 add_4639_8_lut (.I0(GND_net), .I1(n14310[5]), .I2(n518_adj_4674), 
            .I3(n49435), .O(n12999[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4639_8 (.CI(n49435), .I0(n14310[5]), .I1(n518_adj_4674), 
            .CO(n49436));
    SB_LUT4 add_4639_7_lut (.I0(GND_net), .I1(n14310[4]), .I2(n445_adj_4675), 
            .I3(n49434), .O(n12999[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4616_5_lut (.I0(GND_net), .I1(n13844[2]), .I2(n299_adj_4676), 
            .I3(n48845), .O(n12488[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4616_5 (.CI(n48845), .I0(n13844[2]), .I1(n299_adj_4676), 
            .CO(n48846));
    SB_LUT4 add_4616_4_lut (.I0(GND_net), .I1(n13844[1]), .I2(n226_adj_4677), 
            .I3(n48844), .O(n12488[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4639_7 (.CI(n49434), .I0(n14310[4]), .I1(n445_adj_4675), 
            .CO(n49435));
    SB_LUT4 add_4639_6_lut (.I0(GND_net), .I1(n14310[3]), .I2(n372_adj_4678), 
            .I3(n49433), .O(n12999[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4639_6 (.CI(n49433), .I0(n14310[3]), .I1(n372_adj_4678), 
            .CO(n49434));
    SB_LUT4 add_4639_5_lut (.I0(GND_net), .I1(n14310[2]), .I2(n299_adj_4679), 
            .I3(n49432), .O(n12999[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4639_5 (.CI(n49432), .I0(n14310[2]), .I1(n299_adj_4679), 
            .CO(n49433));
    SB_LUT4 add_4639_4_lut (.I0(GND_net), .I1(n14310[1]), .I2(n226_adj_4680), 
            .I3(n49431), .O(n12999[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4616_4 (.CI(n48844), .I0(n13844[1]), .I1(n226_adj_4677), 
            .CO(n48845));
    SB_CARRY add_4639_4 (.CI(n49431), .I0(n14310[1]), .I1(n226_adj_4680), 
            .CO(n49432));
    SB_LUT4 add_4616_3_lut (.I0(GND_net), .I1(n13844[0]), .I2(n153), .I3(n48843), 
            .O(n12488[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4639_3_lut (.I0(GND_net), .I1(n14310[0]), .I2(n153_adj_4681), 
            .I3(n49430), .O(n12999[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4639_3 (.CI(n49430), .I0(n14310[0]), .I1(n153_adj_4681), 
            .CO(n49431));
    SB_CARRY add_4616_3 (.CI(n48843), .I0(n13844[0]), .I1(n153), .CO(n48844));
    SB_LUT4 add_4616_2_lut (.I0(GND_net), .I1(n11_adj_4682), .I2(n80), 
            .I3(GND_net), .O(n12488[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4616_2 (.CI(GND_net), .I0(n11_adj_4682), .I1(n80), .CO(n48843));
    SB_LUT4 add_4639_2_lut (.I0(GND_net), .I1(n11_adj_4683), .I2(n80_adj_4684), 
            .I3(GND_net), .O(n12999[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4639_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5022_11_lut (.I0(GND_net), .I1(n20050[8]), .I2(n770_adj_4685), 
            .I3(n48842), .O(n19852[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5022_10_lut (.I0(GND_net), .I1(n20050[7]), .I2(n697_adj_4686), 
            .I3(n48841), .O(n19852[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4639_2 (.CI(GND_net), .I0(n11_adj_4683), .I1(n80_adj_4684), 
            .CO(n49430));
    SB_LUT4 add_4699_21_lut (.I0(GND_net), .I1(n15476[18]), .I2(GND_net), 
            .I3(n49429), .O(n14310[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_10 (.CI(n48841), .I0(n20050[7]), .I1(n697_adj_4686), 
            .CO(n48842));
    SB_LUT4 add_5022_9_lut (.I0(GND_net), .I1(n20050[6]), .I2(n624_adj_4687), 
            .I3(n48840), .O(n19852[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4699_20_lut (.I0(GND_net), .I1(n15476[17]), .I2(GND_net), 
            .I3(n49428), .O(n14310[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_9 (.CI(n48840), .I0(n20050[6]), .I1(n624_adj_4687), 
            .CO(n48841));
    SB_LUT4 add_5022_8_lut (.I0(GND_net), .I1(n20050[5]), .I2(n551_adj_4688), 
            .I3(n48839), .O(n19852[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4699_20 (.CI(n49428), .I0(n15476[17]), .I1(GND_net), 
            .CO(n49429));
    SB_LUT4 add_4699_19_lut (.I0(GND_net), .I1(n15476[16]), .I2(GND_net), 
            .I3(n49427), .O(n14310[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_8 (.CI(n48839), .I0(n20050[5]), .I1(n551_adj_4688), 
            .CO(n48840));
    SB_LUT4 add_5022_7_lut (.I0(GND_net), .I1(n20050[4]), .I2(n478_adj_4689), 
            .I3(n48838), .O(n19852[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4699_19 (.CI(n49427), .I0(n15476[16]), .I1(GND_net), 
            .CO(n49428));
    SB_CARRY add_5022_7 (.CI(n48838), .I0(n20050[4]), .I1(n478_adj_4689), 
            .CO(n48839));
    SB_LUT4 add_4699_18_lut (.I0(GND_net), .I1(n15476[15]), .I2(GND_net), 
            .I3(n49426), .O(n14310[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5022_6_lut (.I0(GND_net), .I1(n20050[3]), .I2(n405_adj_4690), 
            .I3(n48837), .O(n19852[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4699_18 (.CI(n49426), .I0(n15476[15]), .I1(GND_net), 
            .CO(n49427));
    SB_CARRY add_5022_6 (.CI(n48837), .I0(n20050[3]), .I1(n405_adj_4690), 
            .CO(n48838));
    SB_LUT4 add_5022_5_lut (.I0(GND_net), .I1(n20050[2]), .I2(n332_adj_4691), 
            .I3(n48836), .O(n19852[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9972_bdd_4_lut_49597 (.I0(n9972), .I1(n63055), .I2(setpoint[16]), 
            .I3(n4744), .O(n66681));
    defparam n9972_bdd_4_lut_49597.LUT_INIT = 16'he4aa;
    SB_LUT4 n66681_bdd_4_lut (.I0(n66681), .I1(n535[16]), .I2(n455[16]), 
            .I3(n4744), .O(n66684));
    defparam n66681_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_4699_17_lut (.I0(GND_net), .I1(n15476[14]), .I2(GND_net), 
            .I3(n49425), .O(n14310[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_5 (.CI(n48836), .I0(n20050[2]), .I1(n332_adj_4691), 
            .CO(n48837));
    SB_LUT4 add_5022_4_lut (.I0(GND_net), .I1(n20050[1]), .I2(n259_adj_4692), 
            .I3(n48835), .O(n19852[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_4 (.CI(n48835), .I0(n20050[1]), .I1(n259_adj_4692), 
            .CO(n48836));
    SB_CARRY add_4699_17 (.CI(n49425), .I0(n15476[14]), .I1(GND_net), 
            .CO(n49426));
    SB_LUT4 add_5022_3_lut (.I0(GND_net), .I1(n20050[0]), .I2(n186_adj_4693), 
            .I3(n48834), .O(n19852[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_3 (.CI(n48834), .I0(n20050[0]), .I1(n186_adj_4693), 
            .CO(n48835));
    SB_LUT4 add_5022_2_lut (.I0(GND_net), .I1(n44_adj_4694), .I2(n113_adj_4695), 
            .I3(GND_net), .O(n19852[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5022_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4699_16_lut (.I0(GND_net), .I1(n15476[13]), .I2(n1105), 
            .I3(n49424), .O(n14310[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5022_2 (.CI(GND_net), .I0(n44_adj_4694), .I1(n113_adj_4695), 
            .CO(n48834));
    SB_LUT4 add_4677_21_lut (.I0(GND_net), .I1(n15053[18]), .I2(GND_net), 
            .I3(n48833), .O(n13844[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4699_16 (.CI(n49424), .I0(n15476[13]), .I1(n1105), .CO(n49425));
    SB_LUT4 add_4677_20_lut (.I0(GND_net), .I1(n15053[17]), .I2(GND_net), 
            .I3(n48832), .O(n13844[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4699_15_lut (.I0(GND_net), .I1(n15476[12]), .I2(n1032), 
            .I3(n49423), .O(n14310[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_20 (.CI(n48832), .I0(n15053[17]), .I1(GND_net), 
            .CO(n48833));
    SB_LUT4 add_4677_19_lut (.I0(GND_net), .I1(n15053[16]), .I2(GND_net), 
            .I3(n48831), .O(n13844[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4699_15 (.CI(n49423), .I0(n15476[12]), .I1(n1032), .CO(n49424));
    SB_CARRY add_4677_19 (.CI(n48831), .I0(n15053[16]), .I1(GND_net), 
            .CO(n48832));
    SB_LUT4 add_4699_14_lut (.I0(GND_net), .I1(n15476[11]), .I2(n959), 
            .I3(n49422), .O(n14310[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4677_18_lut (.I0(GND_net), .I1(n15053[15]), .I2(GND_net), 
            .I3(n48830), .O(n13844[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4699_14 (.CI(n49422), .I0(n15476[11]), .I1(n959), .CO(n49423));
    SB_CARRY add_4677_18 (.CI(n48830), .I0(n15053[15]), .I1(GND_net), 
            .CO(n48831));
    SB_LUT4 add_4699_13_lut (.I0(GND_net), .I1(n15476[10]), .I2(n886), 
            .I3(n49421), .O(n14310[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4677_17_lut (.I0(GND_net), .I1(n15053[14]), .I2(GND_net), 
            .I3(n48829), .O(n13844[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_17 (.CI(n48829), .I0(n15053[14]), .I1(GND_net), 
            .CO(n48830));
    SB_CARRY add_4699_13 (.CI(n49421), .I0(n15476[10]), .I1(n886), .CO(n49422));
    SB_LUT4 add_4677_16_lut (.I0(GND_net), .I1(n15053[13]), .I2(n1105_adj_4696), 
            .I3(n48828), .O(n13844[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_16 (.CI(n48828), .I0(n15053[13]), .I1(n1105_adj_4696), 
            .CO(n48829));
    SB_LUT4 add_4699_12_lut (.I0(GND_net), .I1(n15476[9]), .I2(n813), 
            .I3(n49420), .O(n14310[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4699_12 (.CI(n49420), .I0(n15476[9]), .I1(n813), .CO(n49421));
    SB_LUT4 add_4699_11_lut (.I0(GND_net), .I1(n15476[8]), .I2(n740), 
            .I3(n49419), .O(n14310[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4677_15_lut (.I0(GND_net), .I1(n15053[12]), .I2(n1032_adj_4697), 
            .I3(n48827), .O(n13844[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4699_11 (.CI(n49419), .I0(n15476[8]), .I1(n740), .CO(n49420));
    SB_LUT4 add_4699_10_lut (.I0(GND_net), .I1(n15476[7]), .I2(n667_adj_4698), 
            .I3(n49418), .O(n14310[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_15 (.CI(n48827), .I0(n15053[12]), .I1(n1032_adj_4697), 
            .CO(n48828));
    SB_CARRY add_4699_10 (.CI(n49418), .I0(n15476[7]), .I1(n667_adj_4698), 
            .CO(n49419));
    SB_LUT4 add_4677_14_lut (.I0(GND_net), .I1(n15053[11]), .I2(n959_adj_4699), 
            .I3(n48826), .O(n13844[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_14 (.CI(n48826), .I0(n15053[11]), .I1(n959_adj_4699), 
            .CO(n48827));
    SB_LUT4 add_4677_13_lut (.I0(GND_net), .I1(n15053[10]), .I2(n886_adj_4700), 
            .I3(n48825), .O(n13844[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_13 (.CI(n48825), .I0(n15053[10]), .I1(n886_adj_4700), 
            .CO(n48826));
    SB_LUT4 add_4677_12_lut (.I0(GND_net), .I1(n15053[9]), .I2(n813_adj_4701), 
            .I3(n48824), .O(n13844[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4699_9_lut (.I0(GND_net), .I1(n15476[6]), .I2(n594_adj_4702), 
            .I3(n49417), .O(n14310[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4699_9 (.CI(n49417), .I0(n15476[6]), .I1(n594_adj_4702), 
            .CO(n49418));
    SB_LUT4 add_4699_8_lut (.I0(GND_net), .I1(n15476[5]), .I2(n521_adj_4703), 
            .I3(n49416), .O(n14310[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_12 (.CI(n48824), .I0(n15053[9]), .I1(n813_adj_4701), 
            .CO(n48825));
    SB_LUT4 add_4677_11_lut (.I0(GND_net), .I1(n15053[8]), .I2(n740_adj_4704), 
            .I3(n48823), .O(n13844[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_11 (.CI(n48823), .I0(n15053[8]), .I1(n740_adj_4704), 
            .CO(n48824));
    SB_CARRY add_4699_8 (.CI(n49416), .I0(n15476[5]), .I1(n521_adj_4703), 
            .CO(n49417));
    SB_LUT4 add_4699_7_lut (.I0(GND_net), .I1(n15476[4]), .I2(n448_adj_4646), 
            .I3(n49415), .O(n14310[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4677_10_lut (.I0(GND_net), .I1(n15053[7]), .I2(n667), 
            .I3(n48822), .O(n13844[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4699_7 (.CI(n49415), .I0(n15476[4]), .I1(n448_adj_4646), 
            .CO(n49416));
    SB_LUT4 add_4699_6_lut (.I0(GND_net), .I1(n15476[3]), .I2(n375_adj_4645), 
            .I3(n49414), .O(n14310[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_10 (.CI(n48822), .I0(n15053[7]), .I1(n667), .CO(n48823));
    SB_LUT4 add_4677_9_lut (.I0(GND_net), .I1(n15053[6]), .I2(n594), .I3(n48821), 
            .O(n13844[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4699_6 (.CI(n49414), .I0(n15476[3]), .I1(n375_adj_4645), 
            .CO(n49415));
    SB_CARRY add_4677_9 (.CI(n48821), .I0(n15053[6]), .I1(n594), .CO(n48822));
    SB_LUT4 add_4677_8_lut (.I0(GND_net), .I1(n15053[5]), .I2(n521), .I3(n48820), 
            .O(n13844[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4699_5_lut (.I0(GND_net), .I1(n15476[2]), .I2(n302_adj_4615), 
            .I3(n49413), .O(n14310[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_8 (.CI(n48820), .I0(n15053[5]), .I1(n521), .CO(n48821));
    SB_LUT4 add_4677_7_lut (.I0(GND_net), .I1(n15053[4]), .I2(n448_adj_4611), 
            .I3(n48819), .O(n13844[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_7 (.CI(n48819), .I0(n15053[4]), .I1(n448_adj_4611), 
            .CO(n48820));
    SB_CARRY add_4699_5 (.CI(n49413), .I0(n15476[2]), .I1(n302_adj_4615), 
            .CO(n49414));
    SB_LUT4 add_4677_6_lut (.I0(GND_net), .I1(n15053[3]), .I2(n375), .I3(n48818), 
            .O(n13844[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result_i0_i22 (.Q(duty[22]), .C(clk16MHz), .E(control_update), 
            .D(n66744), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_4677_6 (.CI(n48818), .I0(n15053[3]), .I1(n375), .CO(n48819));
    SB_LUT4 add_4699_4_lut (.I0(GND_net), .I1(n15476[1]), .I2(n229_adj_4602), 
            .I3(n49412), .O(n14310[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4677_5_lut (.I0(GND_net), .I1(n15053[2]), .I2(n302_adj_4596), 
            .I3(n48817), .O(n13844[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4699_4 (.CI(n49412), .I0(n15476[1]), .I1(n229_adj_4602), 
            .CO(n49413));
    SB_LUT4 add_4699_3_lut (.I0(GND_net), .I1(n15476[0]), .I2(n156_adj_4592), 
            .I3(n49411), .O(n14310[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_3_lut.LUT_INIT = 16'hC33C;
    SB_DFFER result_i0_i21 (.Q(duty[21]), .C(clk16MHz), .E(control_update), 
            .D(n66738), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i20 (.Q(duty[20]), .C(clk16MHz), .E(control_update), 
            .D(n66732), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_4677_5 (.CI(n48817), .I0(n15053[2]), .I1(n302_adj_4596), 
            .CO(n48818));
    SB_DFFER result_i0_i19 (.Q(duty[19]), .C(clk16MHz), .E(control_update), 
            .D(n66726), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i18 (.Q(duty[18]), .C(clk16MHz), .E(control_update), 
            .D(n66708), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i17 (.Q(duty[17]), .C(clk16MHz), .E(control_update), 
            .D(n66690), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i16 (.Q(duty[16]), .C(clk16MHz), .E(control_update), 
            .D(n66684), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i15 (.Q(duty[15]), .C(clk16MHz), .E(control_update), 
            .D(n66666), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i14 (.Q(duty[14]), .C(clk16MHz), .E(control_update), 
            .D(n66660), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i13 (.Q(duty[13]), .C(clk16MHz), .E(control_update), 
            .D(n66570), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i12 (.Q(duty[12]), .C(clk16MHz), .E(control_update), 
            .D(n67098), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i11 (.Q(duty[11]), .C(clk16MHz), .E(control_update), 
            .D(n67092), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i10 (.Q(duty[10]), .C(clk16MHz), .E(control_update), 
            .D(n67086), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i9 (.Q(duty[9]), .C(clk16MHz), .E(control_update), 
            .D(n67080), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i8 (.Q(duty[8]), .C(clk16MHz), .E(control_update), 
            .D(n67074), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i7 (.Q(duty[7]), .C(clk16MHz), .E(control_update), 
            .D(n67068), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i6 (.Q(duty[6]), .C(clk16MHz), .E(control_update), 
            .D(n67062), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i5 (.Q(duty[5]), .C(clk16MHz), .E(control_update), 
            .D(n67056), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i4 (.Q(duty[4]), .C(clk16MHz), .E(control_update), 
            .D(n67050), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i3 (.Q(duty[3]), .C(clk16MHz), .E(control_update), 
            .D(n67044), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i2 (.Q(duty[2]), .C(clk16MHz), .E(control_update), 
            .D(n67032), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFER result_i0_i1 (.Q(duty[1]), .C(clk16MHz), .E(control_update), 
            .D(n67020), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_CARRY add_4699_3 (.CI(n49411), .I0(n15476[0]), .I1(n156_adj_4592), 
            .CO(n49412));
    SB_LUT4 add_4677_4_lut (.I0(GND_net), .I1(n15053[1]), .I2(n229), .I3(n48816), 
            .O(n13844[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_4 (.CI(n48816), .I0(n15053[1]), .I1(n229), .CO(n48817));
    SB_LUT4 add_4677_3_lut (.I0(GND_net), .I1(n15053[0]), .I2(n156), .I3(n48815), 
            .O(n13844[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4677_3 (.CI(n48815), .I0(n15053[0]), .I1(n156), .CO(n48816));
    SB_LUT4 add_4699_2_lut (.I0(GND_net), .I1(n14_adj_4580), .I2(n83_adj_4579), 
            .I3(GND_net), .O(n14310[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4699_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4677_2_lut (.I0(GND_net), .I1(n14), .I2(n83), .I3(GND_net), 
            .O(n13844[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4677_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4699_2 (.CI(GND_net), .I0(n14_adj_4580), .I1(n83_adj_4579), 
            .CO(n49411));
    SB_CARRY add_4677_2 (.CI(GND_net), .I0(n14), .I1(n83), .CO(n48815));
    SB_LUT4 add_5050_9_lut (.I0(GND_net), .I1(n20291[6]), .I2(n630), .I3(n49410), 
            .O(n20150[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5050_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5050_8_lut (.I0(GND_net), .I1(n20291[5]), .I2(n557_adj_4536), 
            .I3(n49409), .O(n20150[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5050_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5050_8 (.CI(n49409), .I0(n20291[5]), .I1(n557_adj_4536), 
            .CO(n49410));
    SB_LUT4 i48576_3_lut (.I0(n65637), .I1(n455[11]), .I2(n23_adj_4627), 
            .I3(GND_net), .O(n65638));   // verilog/motorControl.v(62[14:31])
    defparam i48576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5050_7_lut (.I0(GND_net), .I1(n20291[4]), .I2(n484_adj_4509), 
            .I3(n49408), .O(n20150[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5050_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5050_7 (.CI(n49408), .I0(n20291[4]), .I1(n484_adj_4509), 
            .CO(n49409));
    SB_LUT4 add_5050_6_lut (.I0(GND_net), .I1(n20291[3]), .I2(n411), .I3(n49407), 
            .O(n20150[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5050_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46731_4_lut (.I0(n21_adj_4628), .I1(n19_adj_4624), .I2(n17_adj_4625), 
            .I3(n9_adj_4623), .O(n63793));
    defparam i46731_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_5050_6 (.CI(n49407), .I0(n20291[3]), .I1(n411), .CO(n49408));
    SB_LUT4 add_5050_5_lut (.I0(GND_net), .I1(n20291[2]), .I2(n338), .I3(n49406), 
            .O(n20150[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5050_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5050_5 (.CI(n49406), .I0(n20291[2]), .I1(n338), .CO(n49407));
    SB_LUT4 mult_24_i498_2_lut (.I0(\Ki[10] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_4704));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_25_25_lut (.I0(GND_net), .I1(n11041[0]), .I2(n10361[0]), 
            .I3(n48352), .O(n455[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5050_4_lut (.I0(GND_net), .I1(n20291[1]), .I2(n265), .I3(n49405), 
            .O(n20150[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5050_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_24_lut (.I0(GND_net), .I1(n360[22]), .I2(n34[22]), 
            .I3(n48351), .O(n455[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_24 (.CI(n48351), .I0(n360[22]), .I1(n34[22]), .CO(n48352));
    SB_LUT4 add_25_23_lut (.I0(GND_net), .I1(n360[21]), .I2(n34[21]), 
            .I3(n48350), .O(n455[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_23 (.CI(n48350), .I0(n360[21]), .I1(n34[21]), .CO(n48351));
    SB_LUT4 i46662_4_lut (.I0(n43), .I1(n25_adj_4626), .I2(n23_adj_4627), 
            .I3(n63793), .O(n63724));
    defparam i46662_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48414_4_lut (.I0(n24_adj_4655), .I1(n8_adj_4652), .I2(n45_adj_4654), 
            .I3(n63718), .O(n65476));   // verilog/motorControl.v(62[14:31])
    defparam i48414_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i47290_3_lut (.I0(n65638), .I1(n455[12]), .I2(n25_adj_4626), 
            .I3(GND_net), .O(n64352));   // verilog/motorControl.v(62[14:31])
    defparam i47290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_28_i4_3_lut (.I0(n62983), .I1(n28[1]), .I2(n455[1]), 
            .I3(GND_net), .O(n4_adj_4705));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48567_3_lut (.I0(n4_adj_4705), .I1(n28[13]), .I2(n455[13]), 
            .I3(GND_net), .O(n65629));   // verilog/motorControl.v(62[35:55])
    defparam i48567_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5050_4 (.CI(n49405), .I0(n20291[1]), .I1(n265), .CO(n49406));
    SB_LUT4 add_5050_3_lut (.I0(GND_net), .I1(n20291[0]), .I2(n192), .I3(n49404), 
            .O(n20150[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5050_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_22_lut (.I0(GND_net), .I1(n360[20]), .I2(n34[20]), 
            .I3(n48349), .O(n455[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_22 (.CI(n48349), .I0(n360[20]), .I1(n34[20]), .CO(n48350));
    SB_CARRY add_5050_3 (.CI(n49404), .I0(n20291[0]), .I1(n192), .CO(n49405));
    SB_LUT4 add_5050_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n20150[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5050_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_21_lut (.I0(GND_net), .I1(n360[19]), .I2(n34[19]), 
            .I3(n48348), .O(n455[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_21 (.CI(n48348), .I0(n360[19]), .I1(n34[19]), .CO(n48349));
    SB_CARRY add_5050_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n49404));
    SB_LUT4 add_25_20_lut (.I0(GND_net), .I1(n360[18]), .I2(n34[18]), 
            .I3(n48347), .O(n455[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_20 (.CI(n48347), .I0(n360[18]), .I1(n34[18]), .CO(n48348));
    SB_LUT4 add_4754_20_lut (.I0(GND_net), .I1(n16401[17]), .I2(GND_net), 
            .I3(n49403), .O(n15476[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_19_lut (.I0(GND_net), .I1(n360[17]), .I2(n34[17]), 
            .I3(n48346), .O(n455[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_19 (.CI(n48346), .I0(n360[17]), .I1(n34[17]), .CO(n48347));
    SB_LUT4 mult_24_i445_2_lut (.I0(\Ki[9] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_4609));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4754_19_lut (.I0(GND_net), .I1(n16401[16]), .I2(GND_net), 
            .I3(n49402), .O(n15476[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_18_lut (.I0(GND_net), .I1(n360[16]), .I2(n34[16]), 
            .I3(n48345), .O(n455[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_18 (.CI(n48345), .I0(n360[16]), .I1(n34[16]), .CO(n48346));
    SB_LUT4 add_25_17_lut (.I0(GND_net), .I1(n360[15]), .I2(n34[15]), 
            .I3(n48344), .O(n455[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4733_20_lut (.I0(GND_net), .I1(n16054[17]), .I2(GND_net), 
            .I3(n48802), .O(n15053[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i134_2_lut (.I0(\Kp[2] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n198));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i134_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4754_19 (.CI(n49402), .I0(n16401[16]), .I1(GND_net), 
            .CO(n49403));
    SB_LUT4 add_4733_19_lut (.I0(GND_net), .I1(n16054[16]), .I2(GND_net), 
            .I3(n48801), .O(n15053[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4754_18_lut (.I0(GND_net), .I1(n16401[15]), .I2(GND_net), 
            .I3(n49401), .O(n15476[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4733_19 (.CI(n48801), .I0(n16054[16]), .I1(GND_net), 
            .CO(n48802));
    SB_CARRY add_4754_18 (.CI(n49401), .I0(n16401[15]), .I1(GND_net), 
            .CO(n49402));
    SB_LUT4 add_4754_17_lut (.I0(GND_net), .I1(n16401[14]), .I2(GND_net), 
            .I3(n49400), .O(n15476[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4733_18_lut (.I0(GND_net), .I1(n16054[15]), .I2(GND_net), 
            .I3(n48800), .O(n15053[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4754_17 (.CI(n49400), .I0(n16401[14]), .I1(GND_net), 
            .CO(n49401));
    SB_CARRY add_4733_18 (.CI(n48800), .I0(n16054[15]), .I1(GND_net), 
            .CO(n48801));
    SB_CARRY add_25_17 (.CI(n48344), .I0(n360[15]), .I1(n34[15]), .CO(n48345));
    SB_LUT4 add_4733_17_lut (.I0(GND_net), .I1(n16054[14]), .I2(GND_net), 
            .I3(n48799), .O(n15053[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_16_lut (.I0(GND_net), .I1(n360[14]), .I2(n34[14]), 
            .I3(n48343), .O(n455[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_16 (.CI(n48343), .I0(n360[14]), .I1(n34[14]), .CO(n48344));
    SB_LUT4 add_4754_16_lut (.I0(GND_net), .I1(n16401[13]), .I2(n1108_adj_4502), 
            .I3(n49399), .O(n15476[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4733_17 (.CI(n48799), .I0(n16054[14]), .I1(GND_net), 
            .CO(n48800));
    SB_LUT4 add_25_15_lut (.I0(GND_net), .I1(n360[13]), .I2(n34[13]), 
            .I3(n48342), .O(n455[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4733_16_lut (.I0(GND_net), .I1(n16054[13]), .I2(n1108), 
            .I3(n48798), .O(n15053[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4733_16 (.CI(n48798), .I0(n16054[13]), .I1(n1108), .CO(n48799));
    SB_CARRY add_4754_16 (.CI(n49399), .I0(n16401[13]), .I1(n1108_adj_4502), 
            .CO(n49400));
    SB_LUT4 add_4733_15_lut (.I0(GND_net), .I1(n16054[12]), .I2(n1035_adj_4499), 
            .I3(n48797), .O(n15053[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4733_15 (.CI(n48797), .I0(n16054[12]), .I1(n1035_adj_4499), 
            .CO(n48798));
    SB_CARRY add_25_15 (.CI(n48342), .I0(n360[13]), .I1(n34[13]), .CO(n48343));
    SB_LUT4 add_4754_15_lut (.I0(GND_net), .I1(n16401[12]), .I2(n1035), 
            .I3(n49398), .O(n15476[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4733_14_lut (.I0(GND_net), .I1(n16054[11]), .I2(n962_adj_4497), 
            .I3(n48796), .O(n15053[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i48568_3_lut (.I0(n65629), .I1(n28[14]), .I2(n455[14]), .I3(GND_net), 
            .O(n65630));   // verilog/motorControl.v(62[35:55])
    defparam i48568_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_4754_15 (.CI(n49398), .I0(n16401[12]), .I1(n1035), .CO(n49399));
    SB_LUT4 add_25_14_lut (.I0(GND_net), .I1(n360[12]), .I2(n34[12]), 
            .I3(n48341), .O(n455[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4733_14 (.CI(n48796), .I0(n16054[11]), .I1(n962_adj_4497), 
            .CO(n48797));
    SB_LUT4 add_4733_13_lut (.I0(GND_net), .I1(n16054[10]), .I2(n889_adj_4496), 
            .I3(n48795), .O(n15053[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4733_13 (.CI(n48795), .I0(n16054[10]), .I1(n889_adj_4496), 
            .CO(n48796));
    SB_LUT4 add_4733_12_lut (.I0(GND_net), .I1(n16054[9]), .I2(n816_adj_4493), 
            .I3(n48794), .O(n15053[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_14 (.CI(n48341), .I0(n360[12]), .I1(n34[12]), .CO(n48342));
    SB_LUT4 add_4754_14_lut (.I0(GND_net), .I1(n16401[11]), .I2(n962), 
            .I3(n49397), .O(n15476[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4733_12 (.CI(n48794), .I0(n16054[9]), .I1(n816_adj_4493), 
            .CO(n48795));
    SB_LUT4 add_25_13_lut (.I0(GND_net), .I1(n360[11]), .I2(n34[11]), 
            .I3(n48340), .O(n455[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4733_11_lut (.I0(GND_net), .I1(n16054[8]), .I2(n743_adj_4492), 
            .I3(n48793), .O(n15053[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_13 (.CI(n48340), .I0(n360[11]), .I1(n34[11]), .CO(n48341));
    SB_LUT4 add_25_12_lut (.I0(GND_net), .I1(n360[10]), .I2(n34[10]), 
            .I3(n48339), .O(n455[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_32_i8_3_lut (.I0(n535[4]), .I1(n535[8]), .I2(n17_adj_4661), 
            .I3(GND_net), .O(n8_adj_4706));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_32_i24_3_lut (.I0(n16_adj_4665), .I1(n535[22]), .I2(n45_adj_4634), 
            .I3(GND_net), .O(n24_adj_4707));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4754_14 (.CI(n49397), .I0(n16401[11]), .I1(n962), .CO(n49398));
    SB_LUT4 mult_24_i494_2_lut (.I0(\Ki[10] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_4608));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i494_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4733_11 (.CI(n48793), .I0(n16054[8]), .I1(n743_adj_4492), 
            .CO(n48794));
    SB_CARRY add_25_12 (.CI(n48339), .I0(n360[10]), .I1(n34[10]), .CO(n48340));
    SB_LUT4 add_4733_10_lut (.I0(GND_net), .I1(n16054[7]), .I2(n670_adj_4491), 
            .I3(n48792), .O(n15053[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_11_lut (.I0(GND_net), .I1(n360[9]), .I2(n34[9]), .I3(n48338), 
            .O(n455[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_11 (.CI(n48338), .I0(n360[9]), .I1(n34[9]), .CO(n48339));
    SB_LUT4 add_4754_13_lut (.I0(GND_net), .I1(n16401[10]), .I2(n889), 
            .I3(n49396), .O(n15476[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4733_10 (.CI(n48792), .I0(n16054[7]), .I1(n670_adj_4491), 
            .CO(n48793));
    SB_LUT4 add_25_10_lut (.I0(GND_net), .I1(n360[8]), .I2(n34[8]), .I3(n48337), 
            .O(n455[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_10 (.CI(n48337), .I0(n360[8]), .I1(n34[8]), .CO(n48338));
    SB_CARRY add_4754_13 (.CI(n49396), .I0(n16401[10]), .I1(n889), .CO(n49397));
    SB_LUT4 add_4733_9_lut (.I0(GND_net), .I1(n16054[6]), .I2(n597_adj_4482), 
            .I3(n48791), .O(n15053[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4733_9 (.CI(n48791), .I0(n16054[6]), .I1(n597_adj_4482), 
            .CO(n48792));
    SB_LUT4 add_4754_12_lut (.I0(GND_net), .I1(n16401[9]), .I2(n816), 
            .I3(n49395), .O(n15476[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4733_8_lut (.I0(GND_net), .I1(n16054[5]), .I2(n524_adj_4479), 
            .I3(n48790), .O(n15053[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4733_8 (.CI(n48790), .I0(n16054[5]), .I1(n524_adj_4479), 
            .CO(n48791));
    SB_LUT4 add_4733_7_lut (.I0(GND_net), .I1(n16054[4]), .I2(n451), .I3(n48789), 
            .O(n15053[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_9_lut (.I0(GND_net), .I1(n360[7]), .I2(n34[7]), .I3(n48336), 
            .O(n455[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_9 (.CI(n48336), .I0(n360[7]), .I1(n34[7]), .CO(n48337));
    SB_CARRY add_4754_12 (.CI(n49395), .I0(n16401[9]), .I1(n816), .CO(n49396));
    SB_LUT4 i46459_4_lut (.I0(n21_adj_4664), .I1(n19_adj_4660), .I2(n17_adj_4661), 
            .I3(n9_adj_4659), .O(n63521));
    defparam i46459_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46412_4_lut (.I0(n43_adj_4636), .I1(n25_adj_4662), .I2(n23_adj_4663), 
            .I3(n63521), .O(n63474));
    defparam i46412_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48420_4_lut (.I0(n24_adj_4707), .I1(n8_adj_4706), .I2(n45_adj_4634), 
            .I3(n63464), .O(n65482));   // verilog/motorControl.v(65[25:41])
    defparam i48420_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_4733_7 (.CI(n48789), .I0(n16054[4]), .I1(n451), .CO(n48790));
    SB_LUT4 i47320_3_lut (.I0(n65180), .I1(n535[12]), .I2(n25_adj_4662), 
            .I3(GND_net), .O(n64382));   // verilog/motorControl.v(65[25:41])
    defparam i47320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_25_8_lut (.I0(GND_net), .I1(n360[6]), .I2(n34[6]), .I3(n48335), 
            .O(n455[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_8 (.CI(n48335), .I0(n360[6]), .I1(n34[6]), .CO(n48336));
    SB_LUT4 add_4754_11_lut (.I0(GND_net), .I1(n16401[8]), .I2(n743), 
            .I3(n49394), .O(n15476[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4754_11 (.CI(n49394), .I0(n16401[8]), .I1(n743), .CO(n49395));
    SB_LUT4 add_4733_6_lut (.I0(GND_net), .I1(n16054[3]), .I2(n378), .I3(n48788), 
            .O(n15053[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4733_6 (.CI(n48788), .I0(n16054[3]), .I1(n378), .CO(n48789));
    SB_LUT4 mult_23_i351_2_lut (.I0(\Kp[7] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_4703));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i183_2_lut (.I0(\Kp[3] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n271));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(n207[23]), .I1(\Kp[2] ), .I2(n48015), .I3(n207[22]), 
            .O(n59388));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_4733_5_lut (.I0(GND_net), .I1(n16054[2]), .I2(n305), .I3(n48787), 
            .O(n15053[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_7_lut (.I0(GND_net), .I1(n360[5]), .I2(n34[5]), .I3(n48334), 
            .O(n455[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_7 (.CI(n48334), .I0(n360[5]), .I1(n34[5]), .CO(n48335));
    SB_LUT4 add_4754_10_lut (.I0(GND_net), .I1(n16401[7]), .I2(n670), 
            .I3(n49393), .O(n15476[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4754_10 (.CI(n49393), .I0(n16401[7]), .I1(n670), .CO(n49394));
    SB_CARRY add_4733_5 (.CI(n48787), .I0(n16054[2]), .I1(n305), .CO(n48788));
    SB_LUT4 add_25_6_lut (.I0(GND_net), .I1(n360[4]), .I2(n34[4]), .I3(n48333), 
            .O(n455[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_6 (.CI(n48333), .I0(n360[4]), .I1(n34[4]), .CO(n48334));
    SB_LUT4 LessThan_26_i45_2_lut (.I0(deadband[22]), .I1(n455[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4654));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4754_9_lut (.I0(GND_net), .I1(n16401[6]), .I2(n597), .I3(n49392), 
            .O(n15476[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4754_9 (.CI(n49392), .I0(n16401[6]), .I1(n597), .CO(n49393));
    SB_LUT4 LessThan_26_i39_2_lut (.I0(deadband[19]), .I1(n455[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4708));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4754_8_lut (.I0(GND_net), .I1(n16401[5]), .I2(n524), .I3(n49391), 
            .O(n15476[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4733_4_lut (.I0(GND_net), .I1(n16054[1]), .I2(n232), .I3(n48786), 
            .O(n15053[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9972_bdd_4_lut (.I0(n9972), .I1(n63178), .I2(setpoint[12]), 
            .I3(n4744), .O(n67095));
    defparam n9972_bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_CARRY add_4733_4 (.CI(n48786), .I0(n16054[1]), .I1(n232), .CO(n48787));
    SB_LUT4 add_4733_3_lut (.I0(GND_net), .I1(n16054[0]), .I2(n159), .I3(n48785), 
            .O(n15053[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_3_lut.LUT_INIT = 16'hC33C;
    SB_DFFR \PID_CONTROLLER.integral_i0_i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk16MHz), .D(n29778), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk16MHz), .D(n29777), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk16MHz), .D(n29776), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk16MHz), .D(n29775), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk16MHz), .D(n29774), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk16MHz), .D(n29773), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk16MHz), .D(n29772), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk16MHz), .D(n29771), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk16MHz), .D(n29770), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk16MHz), .D(n29769), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk16MHz), .D(n29768), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk16MHz), .D(n29767), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk16MHz), .D(n29766), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk16MHz), .D(n29765), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk16MHz), .D(n29764), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk16MHz), .D(n29763), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk16MHz), .D(n29762), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk16MHz), .D(n29761), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk16MHz), .D(n29760), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk16MHz), .D(n29759), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk16MHz), .D(n29758), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk16MHz), .D(n29757), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_DFFR \PID_CONTROLLER.integral_i0_i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk16MHz), .D(n29754), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_25_5_lut (.I0(GND_net), .I1(n360[3]), .I2(n34[3]), .I3(n48332), 
            .O(n455[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_5 (.CI(n48332), .I0(n360[3]), .I1(n34[3]), .CO(n48333));
    SB_LUT4 LessThan_28_i12_3_lut (.I0(n28[7]), .I1(n28[16]), .I2(n455[16]), 
            .I3(GND_net), .O(n12_adj_4709));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_4754_8 (.CI(n49391), .I0(n16401[5]), .I1(n524), .CO(n49392));
    SB_CARRY add_4733_3 (.CI(n48785), .I0(n16054[0]), .I1(n159), .CO(n48786));
    SB_LUT4 add_25_4_lut (.I0(GND_net), .I1(n360[2]), .I2(n34[2]), .I3(n48331), 
            .O(n455[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_4 (.CI(n48331), .I0(n360[2]), .I1(n34[2]), .CO(n48332));
    SB_LUT4 add_4733_2_lut (.I0(GND_net), .I1(n17_adj_4710), .I2(n86), 
            .I3(GND_net), .O(n15053[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4733_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[23]), 
            .I3(n48498), .O(n535[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_25_3_lut (.I0(GND_net), .I1(n360[1]), .I2(n34[1]), .I3(n48330), 
            .O(n455[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_3 (.CI(n48330), .I0(n360[1]), .I1(n34[1]), .CO(n48331));
    SB_LUT4 add_4754_7_lut (.I0(GND_net), .I1(n16401[4]), .I2(n451_adj_4711), 
            .I3(n49390), .O(n15476[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4733_2 (.CI(GND_net), .I0(n17_adj_4710), .I1(n86), .CO(n48785));
    SB_LUT4 unary_minus_33_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[22]), 
            .I3(n48497), .O(n535[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_24 (.CI(n48497), .I0(GND_net), .I1(n1_adj_4992[22]), 
            .CO(n48498));
    SB_LUT4 add_25_2_lut (.I0(GND_net), .I1(n360[0]), .I2(n34[0]), .I3(GND_net), 
            .O(n455[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_25_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_25_2 (.CI(GND_net), .I0(n360[0]), .I1(n34[0]), .CO(n48330));
    SB_LUT4 unary_minus_33_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[21]), 
            .I3(n48496), .O(n535[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_23 (.CI(n48496), .I0(GND_net), .I1(n1_adj_4992[21]), 
            .CO(n48497));
    SB_LUT4 add_16_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n207[23]), .I3(n48329), .O(n233[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n207[23]), .I3(n48328), .O(n233[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4754_7 (.CI(n49390), .I0(n16401[4]), .I1(n451_adj_4711), 
            .CO(n49391));
    SB_LUT4 add_4754_6_lut (.I0(GND_net), .I1(n16401[3]), .I2(n378_adj_4714), 
            .I3(n49389), .O(n15476[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[20]), 
            .I3(n48495), .O(n535[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_22 (.CI(n48495), .I0(GND_net), .I1(n1_adj_4992[20]), 
            .CO(n48496));
    SB_CARRY add_16_24 (.CI(n48328), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n207[23]), .CO(n48329));
    SB_LUT4 add_16_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n207[23]), .I3(n48327), .O(n233[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4754_6 (.CI(n49389), .I0(n16401[3]), .I1(n378_adj_4714), 
            .CO(n49390));
    SB_LUT4 add_4754_5_lut (.I0(GND_net), .I1(n16401[2]), .I2(n305_adj_4716), 
            .I3(n49388), .O(n15476[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[19]), 
            .I3(n48494), .O(n535[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4754_5 (.CI(n49388), .I0(n16401[2]), .I1(n305_adj_4716), 
            .CO(n49389));
    SB_CARRY unary_minus_33_add_3_21 (.CI(n48494), .I0(GND_net), .I1(n1_adj_4992[19]), 
            .CO(n48495));
    SB_CARRY add_16_23 (.CI(n48327), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n207[23]), .CO(n48328));
    SB_LUT4 unary_minus_33_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[18]), 
            .I3(n48493), .O(n535[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4754_4_lut (.I0(GND_net), .I1(n16401[1]), .I2(n232_adj_4718), 
            .I3(n49387), .O(n15476[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n207[23]), .I3(n48326), .O(n233[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4754_4 (.CI(n49387), .I0(n16401[1]), .I1(n232_adj_4718), 
            .CO(n49388));
    SB_LUT4 add_4754_3_lut (.I0(GND_net), .I1(n16401[0]), .I2(n159_adj_4719), 
            .I3(n49386), .O(n15476[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4754_3 (.CI(n49386), .I0(n16401[0]), .I1(n159_adj_4719), 
            .CO(n49387));
    SB_CARRY unary_minus_33_add_3_20 (.CI(n48493), .I0(GND_net), .I1(n1_adj_4992[18]), 
            .CO(n48494));
    SB_LUT4 unary_minus_33_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[17]), 
            .I3(n48492), .O(n535[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4754_2_lut (.I0(GND_net), .I1(n17_adj_4721), .I2(n86_adj_4722), 
            .I3(GND_net), .O(n15476[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4754_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4754_2 (.CI(GND_net), .I0(n17_adj_4721), .I1(n86_adj_4722), 
            .CO(n49386));
    SB_LUT4 add_4805_19_lut (.I0(GND_net), .I1(n17048[16]), .I2(GND_net), 
            .I3(n49385), .O(n16401[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4805_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_19 (.CI(n48492), .I0(GND_net), .I1(n1_adj_4992[17]), 
            .CO(n48493));
    SB_LUT4 unary_minus_33_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[16]), 
            .I3(n48491), .O(n535[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i232_2_lut (.I0(\Kp[4] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4605));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_944 (.I0(n207[22]), .I1(n20550[1]), .I2(n4_adj_4724), 
            .I3(\Kp[3] ), .O(n20502[2]));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_944.LUT_INIT = 16'hc66c;
    SB_LUT4 add_4805_18_lut (.I0(GND_net), .I1(n17048[15]), .I2(GND_net), 
            .I3(n49384), .O(n16401[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4805_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i46607_4_lut (.I0(n455[16]), .I1(n455[7]), .I2(n28[16]), .I3(n28[7]), 
            .O(n63669));
    defparam i46607_4_lut.LUT_INIT = 16'h7bde;
    SB_CARRY add_4805_18 (.CI(n49384), .I0(n17048[15]), .I1(GND_net), 
            .CO(n49385));
    SB_LUT4 add_4805_17_lut (.I0(GND_net), .I1(n17048[14]), .I2(GND_net), 
            .I3(n49383), .O(n16401[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4805_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4805_17 (.CI(n49383), .I0(n17048[14]), .I1(GND_net), 
            .CO(n49384));
    SB_LUT4 add_4805_16_lut (.I0(GND_net), .I1(n17048[13]), .I2(n1111), 
            .I3(n49382), .O(n16401[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4805_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4805_16 (.CI(n49382), .I0(n17048[13]), .I1(n1111), .CO(n49383));
    SB_LUT4 add_4786_19_lut (.I0(GND_net), .I1(n16763[16]), .I2(GND_net), 
            .I3(n48773), .O(n16054[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4786_18_lut (.I0(GND_net), .I1(n16763[15]), .I2(GND_net), 
            .I3(n48772), .O(n16054[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n67095_bdd_4_lut (.I0(n67095), .I1(n535[12]), .I2(n455[12]), 
            .I3(n4744), .O(n67098));
    defparam n67095_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_4786_18 (.CI(n48772), .I0(n16763[15]), .I1(GND_net), 
            .CO(n48773));
    SB_LUT4 add_4805_15_lut (.I0(GND_net), .I1(n17048[12]), .I2(n1038), 
            .I3(n49381), .O(n16401[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4805_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4786_17_lut (.I0(GND_net), .I1(n16763[14]), .I2(GND_net), 
            .I3(n48771), .O(n16054[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_17 (.CI(n48771), .I0(n16763[14]), .I1(GND_net), 
            .CO(n48772));
    SB_CARRY add_16_22 (.CI(n48326), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n207[23]), .CO(n48327));
    SB_LUT4 add_4786_16_lut (.I0(GND_net), .I1(n16763[13]), .I2(n1111_adj_4725), 
            .I3(n48770), .O(n16054[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_16 (.CI(n48770), .I0(n16763[13]), .I1(n1111_adj_4725), 
            .CO(n48771));
    SB_DFFSR counter_2045_2046__i2 (.Q(counter[1]), .C(clk16MHz), .D(n61[1]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_CARRY add_4805_15 (.CI(n49381), .I0(n17048[12]), .I1(n1038), .CO(n49382));
    SB_LUT4 LessThan_28_i35_rep_95_2_lut (.I0(n455[17]), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n67241));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i35_rep_95_2_lut.LUT_INIT = 16'h6666;
    SB_DFFSR counter_2045_2046__i3 (.Q(counter[2]), .C(clk16MHz), .D(n61[2]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i4 (.Q(counter[3]), .C(clk16MHz), .D(n61[3]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i5 (.Q(counter[4]), .C(clk16MHz), .D(n61[4]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i6 (.Q(counter[5]), .C(clk16MHz), .D(n61[5]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i7 (.Q(counter[6]), .C(clk16MHz), .D(n61[6]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i8 (.Q(counter[7]), .C(clk16MHz), .D(n61[7]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i9 (.Q(counter[8]), .C(clk16MHz), .D(n61[8]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i10 (.Q(counter[9]), .C(clk16MHz), .D(n61[9]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i11 (.Q(counter[10]), .C(clk16MHz), .D(n61[10]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i12 (.Q(counter[11]), .C(clk16MHz), .D(n61[11]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i13 (.Q(counter[12]), .C(clk16MHz), .D(n61[12]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_DFFSR counter_2045_2046__i14 (.Q(counter[13]), .C(clk16MHz), .D(n61[13]), 
            .R(counter_31__N_3714));   // verilog/motorControl.v(25[16:25])
    SB_LUT4 add_4786_15_lut (.I0(GND_net), .I1(n16763[12]), .I2(n1038_adj_4726), 
            .I3(n48769), .O(n16054[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4805_14_lut (.I0(GND_net), .I1(n17048[11]), .I2(n965), 
            .I3(n49380), .O(n16401[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4805_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_15 (.CI(n48769), .I0(n16763[12]), .I1(n1038_adj_4726), 
            .CO(n48770));
    SB_LUT4 mult_24_i543_2_lut (.I0(\Ki[11] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807_adj_4603));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4786_14_lut (.I0(GND_net), .I1(n16763[11]), .I2(n965_adj_4727), 
            .I3(n48768), .O(n16054[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_18 (.CI(n48491), .I0(GND_net), .I1(n1_adj_4992[16]), 
            .CO(n48492));
    SB_CARRY add_4786_14 (.CI(n48768), .I0(n16763[11]), .I1(n965_adj_4727), 
            .CO(n48769));
    SB_CARRY add_4805_14 (.CI(n49380), .I0(n17048[11]), .I1(n965), .CO(n49381));
    SB_DFFR \PID_CONTROLLER.integral_i0_i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk16MHz), .D(n28910), .R(reset));   // verilog/motorControl.v(42[14] 73[8])
    SB_LUT4 add_4786_13_lut (.I0(GND_net), .I1(n16763[10]), .I2(n892), 
            .I3(n48767), .O(n16054[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[15]), 
            .I3(n48490), .O(n535[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4805_13_lut (.I0(GND_net), .I1(n17048[10]), .I2(n892_adj_4729), 
            .I3(n49379), .O(n16401[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4805_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_13 (.CI(n48767), .I0(n16763[10]), .I1(n892), .CO(n48768));
    SB_LUT4 add_4786_12_lut (.I0(GND_net), .I1(n16763[9]), .I2(n819), 
            .I3(n48766), .O(n16054[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4805_13 (.CI(n49379), .I0(n17048[10]), .I1(n892_adj_4729), 
            .CO(n49380));
    SB_CARRY add_4786_12 (.CI(n48766), .I0(n16763[9]), .I1(n819), .CO(n48767));
    SB_CARRY unary_minus_33_add_3_17 (.CI(n48490), .I0(GND_net), .I1(n1_adj_4992[15]), 
            .CO(n48491));
    SB_LUT4 add_4786_11_lut (.I0(GND_net), .I1(n16763[8]), .I2(n746), 
            .I3(n48765), .O(n16054[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[14]), 
            .I3(n48489), .O(n535[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_16 (.CI(n48489), .I0(GND_net), .I1(n1_adj_4992[14]), 
            .CO(n48490));
    SB_LUT4 add_4805_12_lut (.I0(GND_net), .I1(n17048[9]), .I2(n819_adj_4731), 
            .I3(n49378), .O(n16401[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4805_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_11 (.CI(n48765), .I0(n16763[8]), .I1(n746), .CO(n48766));
    SB_LUT4 add_4786_10_lut (.I0(GND_net), .I1(n16763[7]), .I2(n673), 
            .I3(n48764), .O(n16054[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[13]), 
            .I3(n48488), .O(n535[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4805_12 (.CI(n49378), .I0(n17048[9]), .I1(n819_adj_4731), 
            .CO(n49379));
    SB_CARRY add_4786_10 (.CI(n48764), .I0(n16763[7]), .I1(n673), .CO(n48765));
    SB_LUT4 add_4805_11_lut (.I0(GND_net), .I1(n17048[8]), .I2(n746_adj_4733), 
            .I3(n49377), .O(n16401[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4805_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_15 (.CI(n48488), .I0(GND_net), .I1(n1_adj_4992[13]), 
            .CO(n48489));
    SB_LUT4 add_4786_9_lut (.I0(GND_net), .I1(n16763[6]), .I2(n600), .I3(n48763), 
            .O(n16054[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4805_11 (.CI(n49377), .I0(n17048[8]), .I1(n746_adj_4733), 
            .CO(n49378));
    SB_CARRY add_4786_9 (.CI(n48763), .I0(n16763[6]), .I1(n600), .CO(n48764));
    SB_LUT4 add_4805_10_lut (.I0(GND_net), .I1(n17048[7]), .I2(n673_adj_4734), 
            .I3(n49376), .O(n16401[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4805_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4805_10 (.CI(n49376), .I0(n17048[7]), .I1(n673_adj_4734), 
            .CO(n49377));
    SB_LUT4 add_4805_9_lut (.I0(GND_net), .I1(n17048[6]), .I2(n600_adj_4735), 
            .I3(n49375), .O(n16401[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4805_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4805_9 (.CI(n49375), .I0(n17048[6]), .I1(n600_adj_4735), 
            .CO(n49376));
    SB_LUT4 n9972_bdd_4_lut_49934 (.I0(n9972), .I1(n63177), .I2(setpoint[11]), 
            .I3(n4744), .O(n67089));
    defparam n9972_bdd_4_lut_49934.LUT_INIT = 16'he4aa;
    SB_LUT4 add_4786_8_lut (.I0(GND_net), .I1(n16763[5]), .I2(n527), .I3(n48762), 
            .O(n16054[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4805_8_lut (.I0(GND_net), .I1(n17048[5]), .I2(n527_adj_4736), 
            .I3(n49374), .O(n16401[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4805_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[12]), 
            .I3(n48487), .O(n535[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4805_8 (.CI(n49374), .I0(n17048[5]), .I1(n527_adj_4736), 
            .CO(n49375));
    SB_LUT4 add_4805_7_lut (.I0(GND_net), .I1(n17048[4]), .I2(n454), .I3(n49373), 
            .O(n16401[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4805_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_8 (.CI(n48762), .I0(n16763[5]), .I1(n527), .CO(n48763));
    SB_LUT4 add_4786_7_lut (.I0(GND_net), .I1(n16763[4]), .I2(n454_adj_4738), 
            .I3(n48761), .O(n16054[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4805_7 (.CI(n49373), .I0(n17048[4]), .I1(n454), .CO(n49374));
    SB_CARRY add_4786_7 (.CI(n48761), .I0(n16763[4]), .I1(n454_adj_4738), 
            .CO(n48762));
    SB_LUT4 add_4786_6_lut (.I0(GND_net), .I1(n16763[3]), .I2(n381), .I3(n48760), 
            .O(n16054[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n67089_bdd_4_lut (.I0(n67089), .I1(n535[11]), .I2(n455[11]), 
            .I3(n4744), .O(n67092));
    defparam n67089_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_4805_6_lut (.I0(GND_net), .I1(n17048[3]), .I2(n381_adj_4739), 
            .I3(n49372), .O(n16401[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4805_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_6 (.CI(n48760), .I0(n16763[3]), .I1(n381), .CO(n48761));
    SB_LUT4 add_4786_5_lut (.I0(GND_net), .I1(n16763[2]), .I2(n308_adj_4740), 
            .I3(n48759), .O(n16054[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_5 (.CI(n48759), .I0(n16763[2]), .I1(n308_adj_4740), 
            .CO(n48760));
    SB_CARRY add_4805_6 (.CI(n49372), .I0(n17048[3]), .I1(n381_adj_4739), 
            .CO(n49373));
    SB_LUT4 add_4805_5_lut (.I0(GND_net), .I1(n17048[2]), .I2(n308_adj_4741), 
            .I3(n49371), .O(n16401[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4805_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4786_4_lut (.I0(GND_net), .I1(n16763[1]), .I2(n235_adj_4742), 
            .I3(n48758), .O(n16054[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_4 (.CI(n48758), .I0(n16763[1]), .I1(n235_adj_4742), 
            .CO(n48759));
    SB_CARRY add_4805_5 (.CI(n49371), .I0(n17048[2]), .I1(n308_adj_4741), 
            .CO(n49372));
    SB_LUT4 add_4786_3_lut (.I0(GND_net), .I1(n16763[0]), .I2(n162), .I3(n48757), 
            .O(n16054[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_3 (.CI(n48757), .I0(n16763[0]), .I1(n162), .CO(n48758));
    SB_LUT4 add_4786_2_lut (.I0(GND_net), .I1(n20), .I2(n89), .I3(GND_net), 
            .O(n16054[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4786_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4805_4_lut (.I0(GND_net), .I1(n17048[1]), .I2(n235_adj_4743), 
            .I3(n49370), .O(n16401[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4805_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4786_2 (.CI(GND_net), .I0(n20), .I1(n89), .CO(n48757));
    SB_CARRY unary_minus_33_add_3_14 (.CI(n48487), .I0(GND_net), .I1(n1_adj_4992[12]), 
            .CO(n48488));
    SB_CARRY add_4805_4 (.CI(n49370), .I0(n17048[1]), .I1(n235_adj_4743), 
            .CO(n49371));
    SB_LUT4 add_4824_18_lut (.I0(GND_net), .I1(n17373[15]), .I2(GND_net), 
            .I3(n48756), .O(n16763[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4824_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4824_17_lut (.I0(GND_net), .I1(n17373[14]), .I2(GND_net), 
            .I3(n48755), .O(n16763[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4824_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[11]), 
            .I3(n48486), .O(n535[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4805_3_lut (.I0(GND_net), .I1(n17048[0]), .I2(n162_adj_4745), 
            .I3(n49369), .O(n16401[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4805_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4824_17 (.CI(n48755), .I0(n17373[14]), .I1(GND_net), 
            .CO(n48756));
    SB_LUT4 add_4824_16_lut (.I0(GND_net), .I1(n17373[13]), .I2(n1114), 
            .I3(n48754), .O(n16763[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4824_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4805_3 (.CI(n49369), .I0(n17048[0]), .I1(n162_adj_4745), 
            .CO(n49370));
    SB_CARRY add_4824_16 (.CI(n48754), .I0(n17373[13]), .I1(n1114), .CO(n48755));
    SB_LUT4 add_4824_15_lut (.I0(GND_net), .I1(n17373[12]), .I2(n1041), 
            .I3(n48753), .O(n16763[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4824_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4805_2_lut (.I0(GND_net), .I1(n20_adj_4746), .I2(n89_adj_4747), 
            .I3(GND_net), .O(n16401[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4805_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4824_15 (.CI(n48753), .I0(n17373[12]), .I1(n1041), .CO(n48754));
    SB_CARRY add_4805_2 (.CI(GND_net), .I0(n20_adj_4746), .I1(n89_adj_4747), 
            .CO(n49369));
    SB_LUT4 add_4824_14_lut (.I0(GND_net), .I1(n17373[11]), .I2(n968), 
            .I3(n48752), .O(n16763[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4824_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4824_14 (.CI(n48752), .I0(n17373[11]), .I1(n968), .CO(n48753));
    SB_LUT4 add_4839_18_lut (.I0(GND_net), .I1(n17625[15]), .I2(GND_net), 
            .I3(n49368), .O(n17048[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4839_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4824_13_lut (.I0(GND_net), .I1(n17373[10]), .I2(n895), 
            .I3(n48751), .O(n16763[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4824_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4824_13 (.CI(n48751), .I0(n17373[10]), .I1(n895), .CO(n48752));
    SB_LUT4 add_4839_17_lut (.I0(GND_net), .I1(n17625[14]), .I2(GND_net), 
            .I3(n49367), .O(n17048[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4839_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4824_12_lut (.I0(GND_net), .I1(n17373[9]), .I2(n822), 
            .I3(n48750), .O(n16763[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4824_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4824_12 (.CI(n48750), .I0(n17373[9]), .I1(n822), .CO(n48751));
    SB_CARRY add_4839_17 (.CI(n49367), .I0(n17625[14]), .I1(GND_net), 
            .CO(n49368));
    SB_LUT4 add_4824_11_lut (.I0(GND_net), .I1(n17373[8]), .I2(n749), 
            .I3(n48749), .O(n16763[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4824_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4824_11 (.CI(n48749), .I0(n17373[8]), .I1(n749), .CO(n48750));
    SB_LUT4 add_4839_16_lut (.I0(GND_net), .I1(n17625[13]), .I2(n1114_adj_4748), 
            .I3(n49366), .O(n17048[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4839_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4824_10_lut (.I0(GND_net), .I1(n17373[7]), .I2(n676), 
            .I3(n48748), .O(n16763[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4824_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4824_10 (.CI(n48748), .I0(n17373[7]), .I1(n676), .CO(n48749));
    SB_CARRY add_4839_16 (.CI(n49366), .I0(n17625[13]), .I1(n1114_adj_4748), 
            .CO(n49367));
    SB_LUT4 add_4824_9_lut (.I0(GND_net), .I1(n17373[6]), .I2(n603), .I3(n48747), 
            .O(n16763[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4824_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4824_9 (.CI(n48747), .I0(n17373[6]), .I1(n603), .CO(n48748));
    SB_LUT4 add_4824_8_lut (.I0(GND_net), .I1(n17373[5]), .I2(n530), .I3(n48746), 
            .O(n16763[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4824_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4839_15_lut (.I0(GND_net), .I1(n17625[12]), .I2(n1041_adj_4749), 
            .I3(n49365), .O(n17048[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4839_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4824_8 (.CI(n48746), .I0(n17373[5]), .I1(n530), .CO(n48747));
    SB_LUT4 add_4824_7_lut (.I0(GND_net), .I1(n17373[4]), .I2(n457_adj_4750), 
            .I3(n48745), .O(n16763[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4824_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4839_15 (.CI(n49365), .I0(n17625[12]), .I1(n1041_adj_4749), 
            .CO(n49366));
    SB_CARRY add_4824_7 (.CI(n48745), .I0(n17373[4]), .I1(n457_adj_4750), 
            .CO(n48746));
    SB_LUT4 add_4824_6_lut (.I0(GND_net), .I1(n17373[3]), .I2(n384_adj_4751), 
            .I3(n48744), .O(n16763[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4824_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4839_14_lut (.I0(GND_net), .I1(n17625[11]), .I2(n968_adj_4752), 
            .I3(n49364), .O(n17048[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4839_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4824_6 (.CI(n48744), .I0(n17373[3]), .I1(n384_adj_4751), 
            .CO(n48745));
    SB_LUT4 add_4824_5_lut (.I0(GND_net), .I1(n17373[2]), .I2(n311_adj_4753), 
            .I3(n48743), .O(n16763[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4824_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_28_i10_3_lut (.I0(n28[5]), .I1(n28[6]), .I2(n455[6]), 
            .I3(GND_net), .O(n10_adj_4754));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_4839_14 (.CI(n49364), .I0(n17625[11]), .I1(n968_adj_4752), 
            .CO(n49365));
    SB_CARRY add_4824_5 (.CI(n48743), .I0(n17373[2]), .I1(n311_adj_4753), 
            .CO(n48744));
    SB_LUT4 add_4824_4_lut (.I0(GND_net), .I1(n17373[1]), .I2(n238_adj_4755), 
            .I3(n48742), .O(n16763[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4824_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_13 (.CI(n48486), .I0(GND_net), .I1(n1_adj_4992[11]), 
            .CO(n48487));
    SB_LUT4 add_4839_13_lut (.I0(GND_net), .I1(n17625[10]), .I2(n895_adj_4756), 
            .I3(n49363), .O(n17048[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4839_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4824_4 (.CI(n48742), .I0(n17373[1]), .I1(n238_adj_4755), 
            .CO(n48743));
    SB_LUT4 add_4824_3_lut (.I0(GND_net), .I1(n17373[0]), .I2(n165), .I3(n48741), 
            .O(n16763[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4824_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4839_13 (.CI(n49363), .I0(n17625[10]), .I1(n895_adj_4756), 
            .CO(n49364));
    SB_CARRY add_4824_3 (.CI(n48741), .I0(n17373[0]), .I1(n165), .CO(n48742));
    SB_LUT4 add_4824_2_lut (.I0(GND_net), .I1(n23_adj_4757), .I2(n92), 
            .I3(GND_net), .O(n16763[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4824_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[10]), 
            .I3(n48485), .O(n535[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4839_12_lut (.I0(GND_net), .I1(n17625[9]), .I2(n822_adj_4759), 
            .I3(n49362), .O(n17048[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4839_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4824_2 (.CI(GND_net), .I0(n23_adj_4757), .I1(n92), .CO(n48741));
    SB_LUT4 add_4858_17_lut (.I0(GND_net), .I1(n17931[14]), .I2(GND_net), 
            .I3(n48740), .O(n17373[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4858_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4839_12 (.CI(n49362), .I0(n17625[9]), .I1(n822_adj_4759), 
            .CO(n49363));
    SB_LUT4 add_4858_16_lut (.I0(GND_net), .I1(n17931[13]), .I2(n1117), 
            .I3(n48739), .O(n17373[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4858_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4858_16 (.CI(n48739), .I0(n17931[13]), .I1(n1117), .CO(n48740));
    SB_LUT4 add_4839_11_lut (.I0(GND_net), .I1(n17625[8]), .I2(n749_adj_4760), 
            .I3(n49361), .O(n17048[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4839_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4839_11 (.CI(n49361), .I0(n17625[8]), .I1(n749_adj_4760), 
            .CO(n49362));
    SB_CARRY unary_minus_33_add_3_12 (.CI(n48485), .I0(GND_net), .I1(n1_adj_4992[10]), 
            .CO(n48486));
    SB_LUT4 unary_minus_33_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[9]), 
            .I3(n48484), .O(n535[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4858_15_lut (.I0(GND_net), .I1(n17931[12]), .I2(n1044), 
            .I3(n48738), .O(n17373[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4858_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4839_10_lut (.I0(GND_net), .I1(n17625[7]), .I2(n676_adj_4762), 
            .I3(n49360), .O(n17048[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4839_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4858_15 (.CI(n48738), .I0(n17931[12]), .I1(n1044), .CO(n48739));
    SB_LUT4 add_4858_14_lut (.I0(GND_net), .I1(n17931[11]), .I2(n971), 
            .I3(n48737), .O(n17373[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4858_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4839_10 (.CI(n49360), .I0(n17625[7]), .I1(n676_adj_4762), 
            .CO(n49361));
    SB_CARRY add_4858_14 (.CI(n48737), .I0(n17931[11]), .I1(n971), .CO(n48738));
    SB_LUT4 add_4858_13_lut (.I0(GND_net), .I1(n17931[10]), .I2(n898), 
            .I3(n48736), .O(n17373[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4858_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_11 (.CI(n48484), .I0(GND_net), .I1(n1_adj_4992[9]), 
            .CO(n48485));
    SB_CARRY add_4858_13 (.CI(n48736), .I0(n17931[10]), .I1(n898), .CO(n48737));
    SB_LUT4 add_4858_12_lut (.I0(GND_net), .I1(n17931[9]), .I2(n825), 
            .I3(n48735), .O(n17373[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4858_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4839_9_lut (.I0(GND_net), .I1(n17625[6]), .I2(n603_adj_4763), 
            .I3(n49359), .O(n17048[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4839_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4858_12 (.CI(n48735), .I0(n17931[9]), .I1(n825), .CO(n48736));
    SB_LUT4 add_4858_11_lut (.I0(GND_net), .I1(n17931[8]), .I2(n752), 
            .I3(n48734), .O(n17373[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4858_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_33_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[8]), 
            .I3(n48483), .O(n535[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n9972_bdd_4_lut_49929 (.I0(n9972), .I1(n63176), .I2(setpoint[10]), 
            .I3(n4744), .O(n67083));
    defparam n9972_bdd_4_lut_49929.LUT_INIT = 16'he4aa;
    SB_LUT4 add_5002_12_lut (.I0(GND_net), .I1(n19852[9]), .I2(n840_adj_4765), 
            .I3(n48972), .O(n19612[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4839_9 (.CI(n49359), .I0(n17625[6]), .I1(n603_adj_4763), 
            .CO(n49360));
    SB_LUT4 add_16_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n207[23]), .I3(n48325), .O(n233[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_21 (.CI(n48325), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n207[23]), .CO(n48326));
    SB_LUT4 add_4839_8_lut (.I0(GND_net), .I1(n17625[5]), .I2(n530_adj_4766), 
            .I3(n49358), .O(n17048[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4839_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4839_8 (.CI(n49358), .I0(n17625[5]), .I1(n530_adj_4766), 
            .CO(n49359));
    SB_CARRY add_4858_11 (.CI(n48734), .I0(n17931[8]), .I1(n752), .CO(n48735));
    SB_CARRY unary_minus_33_add_3_10 (.CI(n48483), .I0(GND_net), .I1(n1_adj_4992[8]), 
            .CO(n48484));
    SB_LUT4 unary_minus_33_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[7]), 
            .I3(n48482), .O(n535[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n207[22]), .I3(n48324), .O(n233[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4858_10_lut (.I0(GND_net), .I1(n17931[7]), .I2(n679), 
            .I3(n48733), .O(n17373[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4858_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_9 (.CI(n48482), .I0(GND_net), .I1(n1_adj_4992[7]), 
            .CO(n48483));
    SB_LUT4 unary_minus_33_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[6]), 
            .I3(n48481), .O(n535[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_20 (.CI(n48324), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n207[22]), .CO(n48325));
    SB_LUT4 add_4839_7_lut (.I0(GND_net), .I1(n17625[4]), .I2(n457_adj_4768), 
            .I3(n49357), .O(n17048[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4839_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4858_10 (.CI(n48733), .I0(n17931[7]), .I1(n679), .CO(n48734));
    SB_CARRY unary_minus_33_add_3_8 (.CI(n48481), .I0(GND_net), .I1(n1_adj_4992[6]), 
            .CO(n48482));
    SB_LUT4 unary_minus_33_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[5]), 
            .I3(n48480), .O(n535[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4858_9_lut (.I0(GND_net), .I1(n17931[6]), .I2(n606), .I3(n48732), 
            .O(n17373[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4858_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_7 (.CI(n48480), .I0(GND_net), .I1(n1_adj_4992[5]), 
            .CO(n48481));
    SB_LUT4 unary_minus_33_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[4]), 
            .I3(n48479), .O(n535[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4839_7 (.CI(n49357), .I0(n17625[4]), .I1(n457_adj_4768), 
            .CO(n49358));
    SB_CARRY add_4858_9 (.CI(n48732), .I0(n17931[6]), .I1(n606), .CO(n48733));
    SB_CARRY unary_minus_33_add_3_6 (.CI(n48479), .I0(GND_net), .I1(n1_adj_4992[4]), 
            .CO(n48480));
    SB_LUT4 unary_minus_33_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[3]), 
            .I3(n48478), .O(n535[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n207[21]), .I3(n48323), .O(n233[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n67083_bdd_4_lut (.I0(n67083), .I1(n535[10]), .I2(n455[10]), 
            .I3(n4744), .O(n67086));
    defparam n67083_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_4858_8_lut (.I0(GND_net), .I1(n17931[5]), .I2(n533), .I3(n48731), 
            .O(n17373[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4858_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_5 (.CI(n48478), .I0(GND_net), .I1(n1_adj_4992[3]), 
            .CO(n48479));
    SB_LUT4 unary_minus_33_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[2]), 
            .I3(n48477), .O(n535[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_19 (.CI(n48323), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n207[21]), .CO(n48324));
    SB_LUT4 add_16_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n207[20]), .I3(n48322), .O(n233[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4839_6_lut (.I0(GND_net), .I1(n17625[3]), .I2(n384_adj_4772), 
            .I3(n49356), .O(n17048[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4839_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5002_11_lut (.I0(GND_net), .I1(n19852[8]), .I2(n767_adj_4773), 
            .I3(n48971), .O(n19612[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4858_8 (.CI(n48731), .I0(n17931[5]), .I1(n533), .CO(n48732));
    SB_CARRY add_4839_6 (.CI(n49356), .I0(n17625[3]), .I1(n384_adj_4772), 
            .CO(n49357));
    SB_LUT4 add_4839_5_lut (.I0(GND_net), .I1(n17625[2]), .I2(n311_adj_4774), 
            .I3(n49355), .O(n17048[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4839_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4858_7_lut (.I0(GND_net), .I1(n17931[4]), .I2(n460_adj_4775), 
            .I3(n48730), .O(n17373[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4858_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5002_11 (.CI(n48971), .I0(n19852[8]), .I1(n767_adj_4773), 
            .CO(n48972));
    SB_LUT4 LessThan_28_i30_3_lut (.I0(n12_adj_4709), .I1(n28[17]), .I2(n455[17]), 
            .I3(GND_net), .O(n30_adj_4776));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY unary_minus_33_add_3_4 (.CI(n48477), .I0(GND_net), .I1(n1_adj_4992[2]), 
            .CO(n48478));
    SB_CARRY add_4858_7 (.CI(n48730), .I0(n17931[4]), .I1(n460_adj_4775), 
            .CO(n48731));
    SB_LUT4 unary_minus_33_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[1]), 
            .I3(n48476), .O(n535[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4839_5 (.CI(n49355), .I0(n17625[2]), .I1(n311_adj_4774), 
            .CO(n49356));
    SB_LUT4 add_4858_6_lut (.I0(GND_net), .I1(n17931[3]), .I2(n387_adj_4778), 
            .I3(n48729), .O(n17373[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4858_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_33_add_3_3 (.CI(n48476), .I0(GND_net), .I1(n1_adj_4992[1]), 
            .CO(n48477));
    SB_LUT4 unary_minus_33_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4992[0]), 
            .I3(VCC_net), .O(n535[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_33_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4858_6 (.CI(n48729), .I0(n17931[3]), .I1(n387_adj_4778), 
            .CO(n48730));
    SB_CARRY unary_minus_33_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4992[0]), 
            .CO(n48476));
    SB_LUT4 unary_minus_27_add_3_25_lut (.I0(n455[23]), .I1(GND_net), .I2(n1_adj_4993[23]), 
            .I3(n48475), .O(n47_adj_4780)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_16_18 (.CI(n48322), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n207[20]), .CO(n48323));
    SB_LUT4 add_4839_4_lut (.I0(GND_net), .I1(n17625[1]), .I2(n238_adj_4782), 
            .I3(n49354), .O(n17048[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4839_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4858_5_lut (.I0(GND_net), .I1(n17931[2]), .I2(n314), .I3(n48728), 
            .O(n17373[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4858_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[22]), 
            .I3(n48474), .O(n28[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4839_4 (.CI(n49354), .I0(n17625[1]), .I1(n238_adj_4782), 
            .CO(n49355));
    SB_CARRY add_4858_5 (.CI(n48728), .I0(n17931[2]), .I1(n314), .CO(n48729));
    SB_LUT4 add_5002_10_lut (.I0(GND_net), .I1(n19852[7]), .I2(n694_adj_4784), 
            .I3(n48970), .O(n19612[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_24 (.CI(n48474), .I0(GND_net), .I1(n1_adj_4993[22]), 
            .CO(n48475));
    SB_LUT4 add_4858_4_lut (.I0(GND_net), .I1(n17931[1]), .I2(n241_adj_4785), 
            .I3(n48727), .O(n17373[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4858_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4858_4 (.CI(n48727), .I0(n17931[1]), .I1(n241_adj_4785), 
            .CO(n48728));
    SB_LUT4 unary_minus_27_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[21]), 
            .I3(n48473), .O(n28[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4858_3_lut (.I0(GND_net), .I1(n17931[0]), .I2(n168), .I3(n48726), 
            .O(n17373[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4858_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_23 (.CI(n48473), .I0(GND_net), .I1(n1_adj_4993[21]), 
            .CO(n48474));
    SB_LUT4 unary_minus_27_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[20]), 
            .I3(n48472), .O(n28[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4839_3_lut (.I0(GND_net), .I1(n17625[0]), .I2(n165_adj_4788), 
            .I3(n49353), .O(n17048[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4839_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4858_3 (.CI(n48726), .I0(n17931[0]), .I1(n168), .CO(n48727));
    SB_CARRY unary_minus_27_add_3_22 (.CI(n48472), .I0(GND_net), .I1(n1_adj_4993[20]), 
            .CO(n48473));
    SB_LUT4 unary_minus_27_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[19]), 
            .I3(n48471), .O(n28[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4858_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n17373[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4858_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_21 (.CI(n48471), .I0(GND_net), .I1(n1_adj_4993[19]), 
            .CO(n48472));
    SB_LUT4 unary_minus_27_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[18]), 
            .I3(n48470), .O(n28[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4839_3 (.CI(n49353), .I0(n17625[0]), .I1(n165_adj_4788), 
            .CO(n49354));
    SB_CARRY add_4858_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n48726));
    SB_CARRY unary_minus_27_add_3_20 (.CI(n48470), .I0(GND_net), .I1(n1_adj_4993[18]), 
            .CO(n48471));
    SB_LUT4 unary_minus_27_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[17]), 
            .I3(n48469), .O(n28[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5040_10_lut (.I0(GND_net), .I1(n20210[7]), .I2(n700_adj_4792), 
            .I3(n48725), .O(n20050[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_19 (.CI(n48469), .I0(GND_net), .I1(n1_adj_4993[17]), 
            .CO(n48470));
    SB_LUT4 unary_minus_27_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[16]), 
            .I3(n48468), .O(n28[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n207[19]), .I3(n48321), .O(n233[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4839_2_lut (.I0(GND_net), .I1(n23_adj_4794), .I2(n92_adj_4795), 
            .I3(GND_net), .O(n17048[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4839_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5040_9_lut (.I0(GND_net), .I1(n20210[6]), .I2(n627_adj_4796), 
            .I3(n48724), .O(n20050[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_18 (.CI(n48468), .I0(GND_net), .I1(n1_adj_4993[16]), 
            .CO(n48469));
    SB_LUT4 unary_minus_27_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[15]), 
            .I3(n48467), .O(n28[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5040_9 (.CI(n48724), .I0(n20210[6]), .I1(n627_adj_4796), 
            .CO(n48725));
    SB_CARRY unary_minus_27_add_3_17 (.CI(n48467), .I0(GND_net), .I1(n1_adj_4993[15]), 
            .CO(n48468));
    SB_LUT4 unary_minus_27_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[14]), 
            .I3(n48466), .O(n28[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_17 (.CI(n48321), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n207[19]), .CO(n48322));
    SB_CARRY add_4839_2 (.CI(GND_net), .I0(n23_adj_4794), .I1(n92_adj_4795), 
            .CO(n49353));
    SB_LUT4 i46615_4_lut (.I0(n455[16]), .I1(n67215), .I2(n28[16]), .I3(n64658), 
            .O(n63677));
    defparam i46615_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 add_5040_8_lut (.I0(GND_net), .I1(n20210[5]), .I2(n554_adj_4799), 
            .I3(n48723), .O(n20050[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_16 (.CI(n48466), .I0(GND_net), .I1(n1_adj_4993[14]), 
            .CO(n48467));
    SB_LUT4 unary_minus_27_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[13]), 
            .I3(n48465), .O(n28[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n207[18]), .I3(n48320), .O(n233[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_16 (.CI(n48320), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n207[18]), .CO(n48321));
    SB_CARRY add_5040_8 (.CI(n48723), .I0(n20210[5]), .I1(n554_adj_4799), 
            .CO(n48724));
    SB_CARRY unary_minus_27_add_3_15 (.CI(n48465), .I0(GND_net), .I1(n1_adj_4993[13]), 
            .CO(n48466));
    SB_LUT4 unary_minus_27_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[12]), 
            .I3(n48464), .O(n28[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n207[17]), .I3(n48319), .O(n233[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_15 (.CI(n48319), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n207[17]), .CO(n48320));
    SB_LUT4 add_5065_8_lut (.I0(GND_net), .I1(n20400[5]), .I2(n560_adj_4802), 
            .I3(n49352), .O(n20291[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5040_7_lut (.I0(GND_net), .I1(n20210[4]), .I2(n481_adj_4803), 
            .I3(n48722), .O(n20050[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_14 (.CI(n48464), .I0(GND_net), .I1(n1_adj_4993[12]), 
            .CO(n48465));
    SB_LUT4 unary_minus_27_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[11]), 
            .I3(n48463), .O(n28[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n207[16]), .I3(n48318), .O(n233[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_14 (.CI(n48318), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n207[16]), .CO(n48319));
    SB_CARRY add_5040_7 (.CI(n48722), .I0(n20210[4]), .I1(n481_adj_4803), 
            .CO(n48723));
    SB_CARRY unary_minus_27_add_3_13 (.CI(n48463), .I0(GND_net), .I1(n1_adj_4993[11]), 
            .CO(n48464));
    SB_LUT4 unary_minus_27_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[10]), 
            .I3(n48462), .O(n28[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n207[15]), .I3(n48317), .O(n233[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_13 (.CI(n48317), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n207[15]), .CO(n48318));
    SB_LUT4 add_5065_7_lut (.I0(GND_net), .I1(n20400[4]), .I2(n487_adj_4806), 
            .I3(n49351), .O(n20291[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5065_7 (.CI(n49351), .I0(n20400[4]), .I1(n487_adj_4806), 
            .CO(n49352));
    SB_LUT4 add_5040_6_lut (.I0(GND_net), .I1(n20210[3]), .I2(n408_adj_4807), 
            .I3(n48721), .O(n20050[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_12 (.CI(n48462), .I0(GND_net), .I1(n1_adj_4993[10]), 
            .CO(n48463));
    SB_LUT4 unary_minus_27_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[9]), 
            .I3(n48461), .O(n28[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n207[14]), .I3(n48316), .O(n233[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_12 (.CI(n48316), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n207[14]), .CO(n48317));
    SB_CARRY add_5002_10 (.CI(n48970), .I0(n19852[7]), .I1(n694_adj_4784), 
            .CO(n48971));
    SB_LUT4 add_5065_6_lut (.I0(GND_net), .I1(n20400[3]), .I2(n414_adj_4809), 
            .I3(n49350), .O(n20291[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5065_6 (.CI(n49350), .I0(n20400[3]), .I1(n414_adj_4809), 
            .CO(n49351));
    SB_CARRY unary_minus_27_add_3_11 (.CI(n48461), .I0(GND_net), .I1(n1_adj_4993[9]), 
            .CO(n48462));
    SB_LUT4 unary_minus_27_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[8]), 
            .I3(n48460), .O(n28[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5040_6 (.CI(n48721), .I0(n20210[3]), .I1(n408_adj_4807), 
            .CO(n48722));
    SB_CARRY unary_minus_27_add_3_10 (.CI(n48460), .I0(GND_net), .I1(n1_adj_4993[8]), 
            .CO(n48461));
    SB_LUT4 unary_minus_27_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[7]), 
            .I3(n48459), .O(n28[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n207[13]), .I3(n48315), .O(n233[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_11 (.CI(n48315), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n207[13]), .CO(n48316));
    SB_LUT4 add_5002_9_lut (.I0(GND_net), .I1(n19852[6]), .I2(n621_adj_4812), 
            .I3(n48969), .O(n19612[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5065_5_lut (.I0(GND_net), .I1(n20400[2]), .I2(n341_adj_4813), 
            .I3(n49349), .O(n20291[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5040_5_lut (.I0(GND_net), .I1(n20210[2]), .I2(n335_adj_4814), 
            .I3(n48720), .O(n20050[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_9 (.CI(n48459), .I0(GND_net), .I1(n1_adj_4993[7]), 
            .CO(n48460));
    SB_LUT4 unary_minus_27_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[6]), 
            .I3(n48458), .O(n28[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5040_5 (.CI(n48720), .I0(n20210[2]), .I1(n335_adj_4814), 
            .CO(n48721));
    SB_CARRY add_5002_9 (.CI(n48969), .I0(n19852[6]), .I1(n621_adj_4812), 
            .CO(n48970));
    SB_CARRY unary_minus_27_add_3_8 (.CI(n48458), .I0(GND_net), .I1(n1_adj_4993[6]), 
            .CO(n48459));
    SB_CARRY add_5065_5 (.CI(n49349), .I0(n20400[2]), .I1(n341_adj_4813), 
            .CO(n49350));
    SB_LUT4 add_5040_4_lut (.I0(GND_net), .I1(n20210[1]), .I2(n262_adj_4816), 
            .I3(n48719), .O(n20050[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[5]), 
            .I3(n48457), .O(n28[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5065_4_lut (.I0(GND_net), .I1(n20400[1]), .I2(n268_adj_4818), 
            .I3(n49348), .O(n20291[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5040_4 (.CI(n48719), .I0(n20210[1]), .I1(n262_adj_4816), 
            .CO(n48720));
    SB_LUT4 add_5002_8_lut (.I0(GND_net), .I1(n19852[5]), .I2(n548_adj_4819), 
            .I3(n48968), .O(n19612[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_7 (.CI(n48457), .I0(GND_net), .I1(n1_adj_4993[5]), 
            .CO(n48458));
    SB_CARRY add_5002_8 (.CI(n48968), .I0(n19852[5]), .I1(n548_adj_4819), 
            .CO(n48969));
    SB_LUT4 add_5002_7_lut (.I0(GND_net), .I1(n19852[4]), .I2(n475_adj_4820), 
            .I3(n48967), .O(n19612[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n207[12]), .I3(n48314), .O(n233[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_10 (.CI(n48314), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n207[12]), .CO(n48315));
    SB_LUT4 add_5040_3_lut (.I0(GND_net), .I1(n20210[0]), .I2(n189_adj_4821), 
            .I3(n48718), .O(n20050[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[4]), 
            .I3(n48456), .O(n28[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_6 (.CI(n48456), .I0(GND_net), .I1(n1_adj_4993[4]), 
            .CO(n48457));
    SB_LUT4 add_16_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n207[11]), .I3(n48313), .O(n233[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_9 (.CI(n48313), .I0(\PID_CONTROLLER.integral [7]), .I1(n207[11]), 
            .CO(n48314));
    SB_CARRY add_5065_4 (.CI(n49348), .I0(n20400[1]), .I1(n268_adj_4818), 
            .CO(n49349));
    SB_CARRY add_5040_3 (.CI(n48718), .I0(n20210[0]), .I1(n189_adj_4821), 
            .CO(n48719));
    SB_LUT4 unary_minus_27_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[3]), 
            .I3(n48455), .O(n28[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_5 (.CI(n48455), .I0(GND_net), .I1(n1_adj_4993[3]), 
            .CO(n48456));
    SB_LUT4 add_16_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n207[10]), .I3(n48312), .O(n233[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_8 (.CI(n48312), .I0(\PID_CONTROLLER.integral [6]), .I1(n207[10]), 
            .CO(n48313));
    SB_CARRY add_5002_7 (.CI(n48967), .I0(n19852[4]), .I1(n475_adj_4820), 
            .CO(n48968));
    SB_LUT4 add_5065_3_lut (.I0(GND_net), .I1(n20400[0]), .I2(n195_adj_4825), 
            .I3(n49347), .O(n20291[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5040_2_lut (.I0(GND_net), .I1(n47_adj_4826), .I2(n116_adj_4827), 
            .I3(GND_net), .O(n20050[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5040_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[2]), 
            .I3(n48454), .O(n28[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_4 (.CI(n48454), .I0(GND_net), .I1(n1_adj_4993[2]), 
            .CO(n48455));
    SB_LUT4 add_5002_6_lut (.I0(GND_net), .I1(n19852[3]), .I2(n402_adj_4829), 
            .I3(n48966), .O(n19612[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5065_3 (.CI(n49347), .I0(n20400[0]), .I1(n195_adj_4825), 
            .CO(n49348));
    SB_CARRY add_5002_6 (.CI(n48966), .I0(n19852[3]), .I1(n402_adj_4829), 
            .CO(n48967));
    SB_LUT4 add_5002_5_lut (.I0(GND_net), .I1(n19852[2]), .I2(n329_adj_4830), 
            .I3(n48965), .O(n19612[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5065_2_lut (.I0(GND_net), .I1(n53_adj_4831), .I2(n122_adj_4832), 
            .I3(GND_net), .O(n20291[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5065_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5040_2 (.CI(GND_net), .I0(n47_adj_4826), .I1(n116_adj_4827), 
            .CO(n48718));
    SB_CARRY add_5065_2 (.CI(GND_net), .I0(n53_adj_4831), .I1(n122_adj_4832), 
            .CO(n49347));
    SB_CARRY add_5002_5 (.CI(n48965), .I0(n19852[2]), .I1(n329_adj_4830), 
            .CO(n48966));
    SB_LUT4 add_5002_4_lut (.I0(GND_net), .I1(n19852[1]), .I2(n256_adj_4833), 
            .I3(n48964), .O(n19612[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_27_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4993[1]), 
            .I3(n48453), .O(n28[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5002_4 (.CI(n48964), .I0(n19852[1]), .I1(n256_adj_4833), 
            .CO(n48965));
    SB_LUT4 add_16_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n207[9]), .I3(n48311), .O(n233[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_7 (.CI(n48311), .I0(\PID_CONTROLLER.integral [5]), .I1(n207[9]), 
            .CO(n48312));
    SB_LUT4 add_4872_17_lut (.I0(GND_net), .I1(n18152[14]), .I2(GND_net), 
            .I3(n49346), .O(n17625[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4872_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4872_16_lut (.I0(GND_net), .I1(n18152[13]), .I2(n1117_adj_4835), 
            .I3(n49345), .O(n17625[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4872_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_27_add_3_3 (.CI(n48453), .I0(GND_net), .I1(n1_adj_4993[1]), 
            .CO(n48454));
    SB_LUT4 add_16_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n207[8]), .I3(n48310), .O(n233[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_6 (.CI(n48310), .I0(\PID_CONTROLLER.integral [4]), .I1(n207[8]), 
            .CO(n48311));
    SB_LUT4 unary_minus_27_add_3_2_lut (.I0(n38672), .I1(GND_net), .I2(n1_adj_4993[0]), 
            .I3(VCC_net), .O(n62983)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_27_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_27_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4993[0]), 
            .CO(n48453));
    SB_LUT4 unary_minus_20_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[23]), 
            .I3(n48452), .O(n285[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[22]), 
            .I3(n48451), .O(n285[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4872_16 (.CI(n49345), .I0(n18152[13]), .I1(n1117_adj_4835), 
            .CO(n49346));
    SB_LUT4 add_5002_3_lut (.I0(GND_net), .I1(n19852[0]), .I2(n183_adj_4839), 
            .I3(n48963), .O(n19612[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4872_15_lut (.I0(GND_net), .I1(n18152[12]), .I2(n1044_adj_4840), 
            .I3(n49344), .O(n17625[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4872_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5002_3 (.CI(n48963), .I0(n19852[0]), .I1(n183_adj_4839), 
            .CO(n48964));
    SB_CARRY unary_minus_20_add_3_24 (.CI(n48451), .I0(GND_net), .I1(n1_adj_4994[22]), 
            .CO(n48452));
    SB_LUT4 add_5002_2_lut (.I0(GND_net), .I1(n41_adj_4841), .I2(n110_adj_4842), 
            .I3(GND_net), .O(n19612[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4872_15 (.CI(n49344), .I0(n18152[12]), .I1(n1044_adj_4840), 
            .CO(n49345));
    SB_LUT4 add_16_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n207[7]), .I3(n48309), .O(n233[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_5 (.CI(n48309), .I0(\PID_CONTROLLER.integral [3]), .I1(n207[7]), 
            .CO(n48310));
    SB_CARRY add_5002_2 (.CI(GND_net), .I0(n41_adj_4841), .I1(n110_adj_4842), 
            .CO(n48963));
    SB_LUT4 add_4872_14_lut (.I0(GND_net), .I1(n18152[11]), .I2(n971_adj_4843), 
            .I3(n49343), .O(n17625[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4872_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4872_14 (.CI(n49343), .I0(n18152[11]), .I1(n971_adj_4843), 
            .CO(n49344));
    SB_LUT4 unary_minus_20_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[21]), 
            .I3(n48450), .O(n285[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_23 (.CI(n48450), .I0(GND_net), .I1(n1_adj_4994[21]), 
            .CO(n48451));
    SB_LUT4 add_16_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n207[6]), .I3(n48308), .O(n233[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_16_4 (.CI(n48308), .I0(\PID_CONTROLLER.integral [2]), .I1(n207[6]), 
            .CO(n48309));
    SB_LUT4 unary_minus_20_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[20]), 
            .I3(n48449), .O(n285[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i400_2_lut (.I0(\Kp[8] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_4702));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i281_2_lut (.I0(\Kp[5] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n417));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4872_13_lut (.I0(GND_net), .I1(n18152[10]), .I2(n898_adj_4846), 
            .I3(n49342), .O(n17625[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4872_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_22 (.CI(n48449), .I0(GND_net), .I1(n1_adj_4994[20]), 
            .CO(n48450));
    SB_LUT4 unary_minus_20_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[19]), 
            .I3(n48448), .O(n285[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i234_2_lut (.I0(\Kp[4] ), .I1(n207[22]), .I2(GND_net), 
            .I3(GND_net), .O(n347_adj_4848));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i234_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_20_add_3_21 (.CI(n48448), .I0(GND_net), .I1(n1_adj_4994[19]), 
            .CO(n48449));
    SB_LUT4 unary_minus_20_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[18]), 
            .I3(n48447), .O(n285[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4872_13 (.CI(n49342), .I0(n18152[10]), .I1(n898_adj_4846), 
            .CO(n49343));
    SB_CARRY unary_minus_20_add_3_20 (.CI(n48447), .I0(GND_net), .I1(n1_adj_4994[18]), 
            .CO(n48448));
    SB_LUT4 unary_minus_20_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[17]), 
            .I3(n48446), .O(n285[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_19 (.CI(n48446), .I0(GND_net), .I1(n1_adj_4994[17]), 
            .CO(n48447));
    SB_LUT4 unary_minus_20_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[16]), 
            .I3(n48445), .O(n285[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4872_12_lut (.I0(GND_net), .I1(n18152[9]), .I2(n825_adj_4852), 
            .I3(n49341), .O(n17625[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4872_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_18 (.CI(n48445), .I0(GND_net), .I1(n1_adj_4994[16]), 
            .CO(n48446));
    SB_LUT4 unary_minus_20_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[15]), 
            .I3(n48444), .O(n285[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4872_12 (.CI(n49341), .I0(n18152[9]), .I1(n825_adj_4852), 
            .CO(n49342));
    SB_CARRY unary_minus_20_add_3_17 (.CI(n48444), .I0(GND_net), .I1(n1_adj_4994[15]), 
            .CO(n48445));
    SB_LUT4 i1_4_lut_adj_945 (.I0(n20550[1]), .I1(n6_adj_4854), .I2(n347_adj_4848), 
            .I3(n55858), .O(n20502[3]));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_945.LUT_INIT = 16'h6996;
    SB_LUT4 add_4872_11_lut (.I0(GND_net), .I1(n18152[8]), .I2(n752_adj_4855), 
            .I3(n49340), .O(n17625[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4872_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4872_11 (.CI(n49340), .I0(n18152[8]), .I1(n752_adj_4855), 
            .CO(n49341));
    SB_LUT4 unary_minus_20_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[14]), 
            .I3(n48443), .O(n285[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_16 (.CI(n48443), .I0(GND_net), .I1(n1_adj_4994[14]), 
            .CO(n48444));
    SB_LUT4 unary_minus_20_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[13]), 
            .I3(n48442), .O(n285[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_15 (.CI(n48442), .I0(GND_net), .I1(n1_adj_4994[13]), 
            .CO(n48443));
    SB_LUT4 unary_minus_20_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[12]), 
            .I3(n48441), .O(n285[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_16_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n207[5]), .I3(n48307), .O(n233[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4872_10_lut (.I0(GND_net), .I1(n18152[7]), .I2(n679_adj_4859), 
            .I3(n49339), .O(n17625[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4872_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4889_16_lut (.I0(GND_net), .I1(n18408[13]), .I2(n1120), 
            .I3(n48708), .O(n17931[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_14 (.CI(n48441), .I0(GND_net), .I1(n1_adj_4994[12]), 
            .CO(n48442));
    SB_LUT4 unary_minus_20_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[11]), 
            .I3(n48440), .O(n285[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4889_15_lut (.I0(GND_net), .I1(n18408[12]), .I2(n1047), 
            .I3(n48707), .O(n17931[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_13 (.CI(n48440), .I0(GND_net), .I1(n1_adj_4994[11]), 
            .CO(n48441));
    SB_LUT4 unary_minus_20_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[10]), 
            .I3(n48439), .O(n285[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_15 (.CI(n48707), .I0(n18408[12]), .I1(n1047), .CO(n48708));
    SB_CARRY unary_minus_20_add_3_12 (.CI(n48439), .I0(GND_net), .I1(n1_adj_4994[10]), 
            .CO(n48440));
    SB_CARRY add_4872_10 (.CI(n49339), .I0(n18152[7]), .I1(n679_adj_4859), 
            .CO(n49340));
    SB_LUT4 add_4889_14_lut (.I0(GND_net), .I1(n18408[11]), .I2(n974), 
            .I3(n48706), .O(n17931[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_14 (.CI(n48706), .I0(n18408[11]), .I1(n974), .CO(n48707));
    SB_LUT4 unary_minus_20_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[9]), 
            .I3(n48438), .O(n285[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4889_13_lut (.I0(GND_net), .I1(n18408[10]), .I2(n901), 
            .I3(n48705), .O(n17931[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4872_9_lut (.I0(GND_net), .I1(n18152[6]), .I2(n606_adj_4863), 
            .I3(n49338), .O(n17625[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4872_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_11 (.CI(n48438), .I0(GND_net), .I1(n1_adj_4994[9]), 
            .CO(n48439));
    SB_CARRY add_4889_13 (.CI(n48705), .I0(n18408[10]), .I1(n901), .CO(n48706));
    SB_CARRY add_16_3 (.CI(n48307), .I0(\PID_CONTROLLER.integral [1]), .I1(n207[5]), 
            .CO(n48308));
    SB_CARRY add_4872_9 (.CI(n49338), .I0(n18152[6]), .I1(n606_adj_4863), 
            .CO(n49339));
    SB_LUT4 add_4889_12_lut (.I0(GND_net), .I1(n18408[9]), .I2(n828), 
            .I3(n48704), .O(n17931[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[8]), 
            .I3(n48437), .O(n285[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_10 (.CI(n48437), .I0(GND_net), .I1(n1_adj_4994[8]), 
            .CO(n48438));
    SB_CARRY add_4889_12 (.CI(n48704), .I0(n18408[9]), .I1(n828), .CO(n48705));
    SB_LUT4 unary_minus_20_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[7]), 
            .I3(n48436), .O(n285[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4872_8_lut (.I0(GND_net), .I1(n18152[5]), .I2(n533_adj_4866), 
            .I3(n49337), .O(n17625[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4872_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_9 (.CI(n48436), .I0(GND_net), .I1(n1_adj_4994[7]), 
            .CO(n48437));
    SB_CARRY add_4872_8 (.CI(n49337), .I0(n18152[5]), .I1(n533_adj_4866), 
            .CO(n49338));
    SB_LUT4 add_4889_11_lut (.I0(GND_net), .I1(n18408[8]), .I2(n755), 
            .I3(n48703), .O(n17931[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[6]), 
            .I3(n48435), .O(n285[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_8 (.CI(n48435), .I0(GND_net), .I1(n1_adj_4994[6]), 
            .CO(n48436));
    SB_CARRY add_4889_11 (.CI(n48703), .I0(n18408[8]), .I1(n755), .CO(n48704));
    SB_LUT4 unary_minus_20_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[5]), 
            .I3(n48434), .O(n285[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_7 (.CI(n48434), .I0(GND_net), .I1(n1_adj_4994[5]), 
            .CO(n48435));
    SB_LUT4 add_4872_7_lut (.I0(GND_net), .I1(n18152[4]), .I2(n460_adj_4869), 
            .I3(n49336), .O(n17625[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4872_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4889_10_lut (.I0(GND_net), .I1(n18408[7]), .I2(n682), 
            .I3(n48702), .O(n17931[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[4]), 
            .I3(n48433), .O(n285[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_6 (.CI(n48433), .I0(GND_net), .I1(n1_adj_4994[4]), 
            .CO(n48434));
    SB_CARRY add_4889_10 (.CI(n48702), .I0(n18408[7]), .I1(n682), .CO(n48703));
    SB_LUT4 unary_minus_20_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[3]), 
            .I3(n48432), .O(n285[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_5 (.CI(n48432), .I0(GND_net), .I1(n1_adj_4994[3]), 
            .CO(n48433));
    SB_LUT4 add_16_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n207[4]), .I3(GND_net), .O(n233[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_16_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4872_7 (.CI(n49336), .I0(n18152[4]), .I1(n460_adj_4869), 
            .CO(n49337));
    SB_LUT4 add_4889_9_lut (.I0(GND_net), .I1(n18408[6]), .I2(n609), .I3(n48701), 
            .O(n17931[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[2]), 
            .I3(n48431), .O(n285[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4872_6_lut (.I0(GND_net), .I1(n18152[3]), .I2(n387_adj_4873), 
            .I3(n49335), .O(n17625[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4872_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_4 (.CI(n48431), .I0(GND_net), .I1(n1_adj_4994[2]), 
            .CO(n48432));
    SB_CARRY add_4889_9 (.CI(n48701), .I0(n18408[6]), .I1(n609), .CO(n48702));
    SB_LUT4 add_4889_8_lut (.I0(GND_net), .I1(n18408[5]), .I2(n536_adj_4874), 
            .I3(n48700), .O(n17931[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_20_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[1]), 
            .I3(n48430), .O(n285[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_8 (.CI(n48700), .I0(n18408[5]), .I1(n536_adj_4874), 
            .CO(n48701));
    SB_CARRY unary_minus_20_add_3_3 (.CI(n48430), .I0(GND_net), .I1(n1_adj_4994[1]), 
            .CO(n48431));
    SB_LUT4 unary_minus_20_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4994[0]), 
            .I3(VCC_net), .O(n285[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_20_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_20_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4994[0]), 
            .CO(n48430));
    SB_CARRY add_16_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n207[4]), .CO(n48307));
    SB_LUT4 i1_3_lut (.I0(\Kp[0] ), .I1(\Kp[2] ), .I2(\Kp[1] ), .I3(GND_net), 
            .O(n59384));   // verilog/motorControl.v(61[20:26])
    defparam i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY add_4872_6 (.CI(n49335), .I0(n18152[3]), .I1(n387_adj_4873), 
            .CO(n49336));
    SB_LUT4 add_4889_7_lut (.I0(GND_net), .I1(n18408[4]), .I2(n463_adj_4877), 
            .I3(n48699), .O(n17931[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4872_5_lut (.I0(GND_net), .I1(n18152[2]), .I2(n314_adj_4878), 
            .I3(n49334), .O(n17625[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4872_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(\motor_state[23] ), 
            .I3(n48306), .O(n207[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(\motor_state[22] ), 
            .I3(n48305), .O(n207[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_7 (.CI(n48699), .I0(n18408[4]), .I1(n463_adj_4877), 
            .CO(n48700));
    SB_CARRY sub_15_add_2_24 (.CI(n48305), .I0(setpoint[22]), .I1(\motor_state[22] ), 
            .CO(n48306));
    SB_LUT4 sub_15_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(\motor_state[21] ), 
            .I3(n48304), .O(n207[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4889_6_lut (.I0(GND_net), .I1(n18408[3]), .I2(n390_adj_4879), 
            .I3(n48698), .O(n17931[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4872_5 (.CI(n49334), .I0(n18152[2]), .I1(n314_adj_4878), 
            .CO(n49335));
    SB_CARRY add_4889_6 (.CI(n48698), .I0(n18408[3]), .I1(n390_adj_4879), 
            .CO(n48699));
    SB_CARRY sub_15_add_2_23 (.CI(n48304), .I0(setpoint[21]), .I1(\motor_state[21] ), 
            .CO(n48305));
    SB_LUT4 sub_15_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(\motor_state[20] ), 
            .I3(n48303), .O(n207[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4889_5_lut (.I0(GND_net), .I1(n18408[2]), .I2(n317), .I3(n48697), 
            .O(n17931[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_22 (.CI(n48303), .I0(setpoint[20]), .I1(\motor_state[20] ), 
            .CO(n48304));
    SB_LUT4 sub_15_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(\motor_state[19] ), 
            .I3(n48302), .O(n207[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_946 (.I0(n59384), .I1(n207[23]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4724));   // verilog/motorControl.v(61[20:26])
    defparam i1_2_lut_adj_946.LUT_INIT = 16'h8888;
    SB_LUT4 add_4872_4_lut (.I0(GND_net), .I1(n18152[1]), .I2(n241_adj_4880), 
            .I3(n49333), .O(n17625[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4872_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4872_4 (.CI(n49333), .I0(n18152[1]), .I1(n241_adj_4880), 
            .CO(n49334));
    SB_CARRY add_4889_5 (.CI(n48697), .I0(n18408[2]), .I1(n317), .CO(n48698));
    SB_LUT4 add_4872_3_lut (.I0(GND_net), .I1(n18152[0]), .I2(n168_adj_4881), 
            .I3(n49332), .O(n17625[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4872_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4872_3 (.CI(n49332), .I0(n18152[0]), .I1(n168_adj_4881), 
            .CO(n49333));
    SB_LUT4 add_4889_4_lut (.I0(GND_net), .I1(n18408[1]), .I2(n244_adj_4882), 
            .I3(n48696), .O(n17931[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_4 (.CI(n48696), .I0(n18408[1]), .I1(n244_adj_4882), 
            .CO(n48697));
    SB_CARRY sub_15_add_2_21 (.CI(n48302), .I0(setpoint[19]), .I1(\motor_state[19] ), 
            .CO(n48303));
    SB_LUT4 add_4872_2_lut (.I0(GND_net), .I1(n26_adj_4883), .I2(n95_adj_4884), 
            .I3(GND_net), .O(n17625[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4872_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4889_3_lut (.I0(GND_net), .I1(n18408[0]), .I2(n171), .I3(n48695), 
            .O(n17931[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_3 (.CI(n48695), .I0(n18408[0]), .I1(n171), .CO(n48696));
    SB_CARRY add_4872_2 (.CI(GND_net), .I0(n26_adj_4883), .I1(n95_adj_4884), 
            .CO(n49332));
    SB_LUT4 add_4889_2_lut (.I0(GND_net), .I1(n29_adj_4885), .I2(n98), 
            .I3(GND_net), .O(n17931[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4889_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(\motor_state[18] ), 
            .I3(n48301), .O(n207[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_20 (.CI(n48301), .I0(setpoint[18]), .I1(\motor_state[18] ), 
            .CO(n48302));
    SB_LUT4 sub_15_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(\motor_state[17] ), 
            .I3(n48300), .O(n207[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4902_16_lut (.I0(GND_net), .I1(n18600[13]), .I2(n1120_adj_4886), 
            .I3(n49331), .O(n18152[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4902_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4902_15_lut (.I0(GND_net), .I1(n18600[12]), .I2(n1047_adj_4887), 
            .I3(n49330), .O(n18152[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4902_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4889_2 (.CI(GND_net), .I0(n29_adj_4885), .I1(n98), .CO(n48695));
    SB_CARRY sub_15_add_2_19 (.CI(n48300), .I0(setpoint[17]), .I1(\motor_state[17] ), 
            .CO(n48301));
    SB_LUT4 sub_15_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(\motor_state[16] ), 
            .I3(n48299), .O(n207[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4902_15 (.CI(n49330), .I0(n18600[12]), .I1(n1047_adj_4887), 
            .CO(n49331));
    SB_LUT4 add_4902_14_lut (.I0(GND_net), .I1(n18600[11]), .I2(n974_adj_4888), 
            .I3(n49329), .O(n18152[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4902_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4918_15_lut (.I0(GND_net), .I1(n18825[12]), .I2(n1050), 
            .I3(n48694), .O(n18408[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4918_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_18 (.CI(n48299), .I0(setpoint[16]), .I1(\motor_state[16] ), 
            .CO(n48300));
    SB_LUT4 add_4918_14_lut (.I0(GND_net), .I1(n18825[11]), .I2(n977_adj_4889), 
            .I3(n48693), .O(n18408[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4918_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(\motor_state[15] ), 
            .I3(n48298), .O(n207[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4902_14 (.CI(n49329), .I0(n18600[11]), .I1(n974_adj_4888), 
            .CO(n49330));
    SB_LUT4 add_4902_13_lut (.I0(GND_net), .I1(n18600[10]), .I2(n901_adj_4890), 
            .I3(n49328), .O(n18152[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4902_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4918_14 (.CI(n48693), .I0(n18825[11]), .I1(n977_adj_4889), 
            .CO(n48694));
    SB_CARRY add_4902_13 (.CI(n49328), .I0(n18600[10]), .I1(n901_adj_4890), 
            .CO(n49329));
    SB_LUT4 add_4918_13_lut (.I0(GND_net), .I1(n18825[10]), .I2(n904_adj_4891), 
            .I3(n48692), .O(n18408[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4918_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_17 (.CI(n48298), .I0(setpoint[15]), .I1(\motor_state[15] ), 
            .CO(n48299));
    SB_LUT4 sub_15_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(n9), 
            .I3(n48297), .O(n207[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4918_13 (.CI(n48692), .I0(n18825[10]), .I1(n904_adj_4891), 
            .CO(n48693));
    SB_CARRY sub_15_add_2_16 (.CI(n48297), .I0(setpoint[14]), .I1(n9), 
            .CO(n48298));
    SB_LUT4 sub_15_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(\motor_state[13] ), 
            .I3(n48296), .O(n207[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4918_12_lut (.I0(GND_net), .I1(n18825[9]), .I2(n831_adj_4893), 
            .I3(n48691), .O(n18408[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4918_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_15 (.CI(n48296), .I0(setpoint[13]), .I1(\motor_state[13] ), 
            .CO(n48297));
    SB_CARRY add_4918_12 (.CI(n48691), .I0(n18825[9]), .I1(n831_adj_4893), 
            .CO(n48692));
    SB_LUT4 add_4902_12_lut (.I0(GND_net), .I1(n18600[9]), .I2(n828_adj_4894), 
            .I3(n49327), .O(n18152[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4902_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4902_12 (.CI(n49327), .I0(n18600[9]), .I1(n828_adj_4894), 
            .CO(n49328));
    SB_LUT4 add_4902_11_lut (.I0(GND_net), .I1(n18600[8]), .I2(n755_adj_4895), 
            .I3(n49326), .O(n18152[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4902_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4918_11_lut (.I0(GND_net), .I1(n18825[8]), .I2(n758_adj_4896), 
            .I3(n48690), .O(n18408[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4918_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_15_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(\motor_state[12] ), 
            .I3(n48295), .O(n207[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_14 (.CI(n48295), .I0(setpoint[12]), .I1(\motor_state[12] ), 
            .CO(n48296));
    SB_CARRY add_4918_11 (.CI(n48690), .I0(n18825[8]), .I1(n758_adj_4896), 
            .CO(n48691));
    SB_LUT4 sub_15_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(\motor_state[11] ), 
            .I3(n48294), .O(n207[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_15_add_2_13 (.CI(n48294), .I0(setpoint[11]), .I1(\motor_state[11] ), 
            .CO(n48295));
    SB_LUT4 i32495_4_lut (.I0(n20550[1]), .I1(\Kp[3] ), .I2(n4_adj_4724), 
            .I3(n207[22]), .O(n6_adj_4854));   // verilog/motorControl.v(61[20:26])
    defparam i32495_4_lut.LUT_INIT = 16'he800;
    SB_LUT4 add_4918_10_lut (.I0(GND_net), .I1(n18825[7]), .I2(n685_adj_4897), 
            .I3(n48689), .O(n18408[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4918_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4902_11 (.CI(n49326), .I0(n18600[8]), .I1(n755_adj_4895), 
            .CO(n49327));
    SB_LUT4 add_4902_10_lut (.I0(GND_net), .I1(n18600[7]), .I2(n682_adj_4898), 
            .I3(n49325), .O(n18152[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4902_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4918_10 (.CI(n48689), .I0(n18825[7]), .I1(n685_adj_4897), 
            .CO(n48690));
    SB_LUT4 sub_15_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(\motor_state[10] ), 
            .I3(n48293), .O(n207[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_15_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4902_10 (.CI(n49325), .I0(n18600[7]), .I1(n682_adj_4898), 
            .CO(n49326));
    SB_LUT4 add_4902_9_lut (.I0(GND_net), .I1(n18600[6]), .I2(n609_adj_4899), 
            .I3(n49324), .O(n18152[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4902_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4918_9_lut (.I0(GND_net), .I1(n18825[6]), .I2(n612_adj_4900), 
            .I3(n48688), .O(n18408[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4918_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4902_9 (.CI(n49324), .I0(n18600[6]), .I1(n609_adj_4899), 
            .CO(n49325));
    SB_LUT4 add_4902_8_lut (.I0(GND_net), .I1(n18600[5]), .I2(n536_adj_4901), 
            .I3(n49323), .O(n18152[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4902_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4902_8 (.CI(n49323), .I0(n18600[5]), .I1(n536_adj_4901), 
            .CO(n49324));
    SB_CARRY add_4918_9 (.CI(n48688), .I0(n18825[6]), .I1(n612_adj_4900), 
            .CO(n48689));
    SB_LUT4 mult_24_i547_2_lut (.I0(\Ki[11] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813_adj_4701));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4902_7_lut (.I0(GND_net), .I1(n18600[4]), .I2(n463_adj_4902), 
            .I3(n49322), .O(n18152[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4902_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_23_i46_2_lut (.I0(\Kp[0] ), .I1(n207[23]), .I2(GND_net), 
            .I3(GND_net), .O(n68_adj_4903));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n9972_bdd_4_lut_49924 (.I0(n9972), .I1(n63175), .I2(setpoint[9]), 
            .I3(n4744), .O(n67077));
    defparam n9972_bdd_4_lut_49924.LUT_INIT = 16'he4aa;
    SB_CARRY add_4902_7 (.CI(n49322), .I0(n18600[4]), .I1(n463_adj_4902), 
            .CO(n49323));
    SB_LUT4 add_4918_8_lut (.I0(GND_net), .I1(n18825[5]), .I2(n539_adj_4904), 
            .I3(n48687), .O(n18408[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4918_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4918_8 (.CI(n48687), .I0(n18825[5]), .I1(n539_adj_4904), 
            .CO(n48688));
    SB_LUT4 i32433_2_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n48015));   // verilog/motorControl.v(61[20:26])
    defparam i32433_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4902_6_lut (.I0(GND_net), .I1(n18600[3]), .I2(n390_adj_4905), 
            .I3(n49321), .O(n18152[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4902_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4918_7_lut (.I0(GND_net), .I1(n18825[4]), .I2(n466_adj_4906), 
            .I3(n48686), .O(n18408[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4918_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4918_7 (.CI(n48686), .I0(n18825[4]), .I1(n466_adj_4906), 
            .CO(n48687));
    SB_LUT4 add_4918_6_lut (.I0(GND_net), .I1(n18825[3]), .I2(n393_adj_4907), 
            .I3(n48685), .O(n18408[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4918_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4902_6 (.CI(n49321), .I0(n18600[3]), .I1(n390_adj_4905), 
            .CO(n49322));
    SB_CARRY add_4918_6 (.CI(n48685), .I0(n18825[3]), .I1(n393_adj_4907), 
            .CO(n48686));
    SB_LUT4 add_4918_5_lut (.I0(GND_net), .I1(n18825[2]), .I2(n320_adj_4908), 
            .I3(n48684), .O(n18408[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4918_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4902_5_lut (.I0(GND_net), .I1(n18600[2]), .I2(n317_adj_4909), 
            .I3(n49320), .O(n18152[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4902_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4918_5 (.CI(n48684), .I0(n18825[2]), .I1(n320_adj_4908), 
            .CO(n48685));
    SB_LUT4 add_4918_4_lut (.I0(GND_net), .I1(n18825[1]), .I2(n247_adj_4910), 
            .I3(n48683), .O(n18408[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4918_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4902_5 (.CI(n49320), .I0(n18600[2]), .I1(n317_adj_4909), 
            .CO(n49321));
    SB_LUT4 add_4902_4_lut (.I0(GND_net), .I1(n18600[1]), .I2(n244_adj_4911), 
            .I3(n49319), .O(n18152[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4902_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4918_4 (.CI(n48683), .I0(n18825[1]), .I1(n247_adj_4910), 
            .CO(n48684));
    SB_LUT4 add_4918_3_lut (.I0(GND_net), .I1(n18825[0]), .I2(n174_adj_4912), 
            .I3(n48682), .O(n18408[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4918_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4902_4 (.CI(n49319), .I0(n18600[1]), .I1(n244_adj_4911), 
            .CO(n49320));
    SB_CARRY add_4918_3 (.CI(n48682), .I0(n18825[0]), .I1(n174_adj_4912), 
            .CO(n48683));
    SB_LUT4 add_4918_2_lut (.I0(GND_net), .I1(n32_adj_4913), .I2(n101_adj_4914), 
            .I3(GND_net), .O(n18408[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4918_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4902_3_lut (.I0(GND_net), .I1(n18600[0]), .I2(n171_adj_4915), 
            .I3(n49318), .O(n18152[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4902_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4918_2 (.CI(GND_net), .I0(n32_adj_4913), .I1(n101_adj_4914), 
            .CO(n48682));
    SB_LUT4 add_5056_9_lut (.I0(GND_net), .I1(n20336[6]), .I2(n630_adj_4916), 
            .I3(n48681), .O(n20210[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5056_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4902_3 (.CI(n49318), .I0(n18600[0]), .I1(n171_adj_4915), 
            .CO(n49319));
    SB_LUT4 add_5056_8_lut (.I0(GND_net), .I1(n20336[5]), .I2(n557_adj_4917), 
            .I3(n48680), .O(n20210[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5056_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5056_8 (.CI(n48680), .I0(n20336[5]), .I1(n557_adj_4917), 
            .CO(n48681));
    SB_LUT4 add_4902_2_lut (.I0(GND_net), .I1(n29_adj_4918), .I2(n98_adj_4919), 
            .I3(GND_net), .O(n18152[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4902_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5056_7_lut (.I0(GND_net), .I1(n20336[4]), .I2(n484_adj_4920), 
            .I3(n48679), .O(n20210[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5056_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5056_7 (.CI(n48679), .I0(n20336[4]), .I1(n484_adj_4920), 
            .CO(n48680));
    SB_CARRY add_4902_2 (.CI(GND_net), .I0(n29_adj_4918), .I1(n98_adj_4919), 
            .CO(n49318));
    SB_LUT4 add_5056_6_lut (.I0(GND_net), .I1(n20336[3]), .I2(n411_adj_4921), 
            .I3(n48678), .O(n20210[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5056_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5078_7_lut (.I0(GND_net), .I1(n57863), .I2(n490_adj_4922), 
            .I3(n49317), .O(n20400[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5078_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5056_6 (.CI(n48678), .I0(n20336[3]), .I1(n411_adj_4921), 
            .CO(n48679));
    SB_LUT4 add_5078_6_lut (.I0(GND_net), .I1(n20481[3]), .I2(n417_adj_4923), 
            .I3(n49316), .O(n20400[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5078_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5056_5_lut (.I0(GND_net), .I1(n20336[2]), .I2(n338_adj_4924), 
            .I3(n48677), .O(n20210[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5056_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5056_5 (.CI(n48677), .I0(n20336[2]), .I1(n338_adj_4924), 
            .CO(n48678));
    SB_CARRY add_5078_6 (.CI(n49316), .I0(n20481[3]), .I1(n417_adj_4923), 
            .CO(n49317));
    SB_LUT4 add_5078_5_lut (.I0(GND_net), .I1(n20481[2]), .I2(n344_adj_4925), 
            .I3(n49315), .O(n20400[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5078_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5056_4_lut (.I0(GND_net), .I1(n20336[1]), .I2(n265_adj_4926), 
            .I3(n48676), .O(n20210[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5056_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5056_4 (.CI(n48676), .I0(n20336[1]), .I1(n265_adj_4926), 
            .CO(n48677));
    SB_CARRY add_5078_5 (.CI(n49315), .I0(n20481[2]), .I1(n344_adj_4925), 
            .CO(n49316));
    SB_LUT4 add_5056_3_lut (.I0(GND_net), .I1(n20336[0]), .I2(n192_adj_4927), 
            .I3(n48675), .O(n20210[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5056_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5056_3 (.CI(n48675), .I0(n20336[0]), .I1(n192_adj_4927), 
            .CO(n48676));
    SB_LUT4 add_5056_2_lut (.I0(GND_net), .I1(n50_adj_4928), .I2(n119_adj_4929), 
            .I3(GND_net), .O(n20210[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5056_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5078_4_lut (.I0(GND_net), .I1(n20481[1]), .I2(n271_adj_4930), 
            .I3(n49314), .O(n20400[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5078_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5078_4 (.CI(n49314), .I0(n20481[1]), .I1(n271_adj_4930), 
            .CO(n49315));
    SB_CARRY add_5056_2 (.CI(GND_net), .I0(n50_adj_4928), .I1(n119_adj_4929), 
            .CO(n48675));
    SB_LUT4 add_5078_3_lut (.I0(GND_net), .I1(n20481[0]), .I2(n198_adj_4931), 
            .I3(n49313), .O(n20400[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5078_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4945_14_lut (.I0(GND_net), .I1(n19186[11]), .I2(n980_adj_4932), 
            .I3(n48674), .O(n18825[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4945_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4945_13_lut (.I0(GND_net), .I1(n19186[10]), .I2(n907_adj_4933), 
            .I3(n48673), .O(n18825[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4945_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5078_3 (.CI(n49313), .I0(n20481[0]), .I1(n198_adj_4931), 
            .CO(n49314));
    SB_CARRY add_4945_13 (.CI(n48673), .I0(n19186[10]), .I1(n907_adj_4933), 
            .CO(n48674));
    SB_LUT4 add_4945_12_lut (.I0(GND_net), .I1(n19186[9]), .I2(n834_adj_4934), 
            .I3(n48672), .O(n18825[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4945_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n67077_bdd_4_lut (.I0(n67077), .I1(n535[9]), .I2(n455[9]), 
            .I3(n4744), .O(n67080));
    defparam n67077_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_5078_2_lut (.I0(GND_net), .I1(n56_adj_4935), .I2(n125_adj_4936), 
            .I3(GND_net), .O(n20400[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5078_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4945_12 (.CI(n48672), .I0(n19186[9]), .I1(n834_adj_4934), 
            .CO(n48673));
    SB_LUT4 add_4945_11_lut (.I0(GND_net), .I1(n19186[8]), .I2(n761_adj_4937), 
            .I3(n48671), .O(n18825[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4945_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5078_2 (.CI(GND_net), .I0(n56_adj_4935), .I1(n125_adj_4936), 
            .CO(n49313));
    SB_CARRY add_4945_11 (.CI(n48671), .I0(n19186[8]), .I1(n761_adj_4937), 
            .CO(n48672));
    SB_LUT4 add_4945_10_lut (.I0(GND_net), .I1(n19186[7]), .I2(n688_adj_4938), 
            .I3(n48670), .O(n18825[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4945_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4945_10 (.CI(n48670), .I0(n19186[7]), .I1(n688_adj_4938), 
            .CO(n48671));
    SB_LUT4 add_4930_15_lut (.I0(GND_net), .I1(n18990[12]), .I2(n1050_adj_4939), 
            .I3(n49312), .O(n18600[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4930_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4945_9_lut (.I0(GND_net), .I1(n19186[6]), .I2(n615_adj_4940), 
            .I3(n48669), .O(n18825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4945_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4945_9 (.CI(n48669), .I0(n19186[6]), .I1(n615_adj_4940), 
            .CO(n48670));
    SB_LUT4 i42659_3_lut (.I0(n207[23]), .I1(n59384), .I2(\Kp[3] ), .I3(GND_net), 
            .O(n55858));   // verilog/motorControl.v(61[20:26])
    defparam i42659_3_lut.LUT_INIT = 16'h2828;
    SB_LUT4 i32442_3_lut (.I0(n207[23]), .I1(n48010), .I2(n49517), .I3(GND_net), 
            .O(n20550[1]));   // verilog/motorControl.v(61[20:26])
    defparam i32442_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_23_i330_2_lut (.I0(\Kp[6] ), .I1(n207[21]), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_4595));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_947 (.I0(n207[23]), .I1(\Kp[5] ), .I2(n49517), 
            .I3(n207[22]), .O(n59374));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_947.LUT_INIT = 16'hc60a;
    SB_LUT4 i1_rep_356_2_lut (.I0(n20550[1]), .I1(n55858), .I2(GND_net), 
            .I3(GND_net), .O(n67502));   // verilog/motorControl.v(61[20:26])
    defparam i1_rep_356_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_948 (.I0(n48010), .I1(n59374), .I2(\Kp[4] ), 
            .I3(n207[23]), .O(n59378));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_948.LUT_INIT = 16'h9666;
    SB_LUT4 i48909_4_lut (.I0(n30_adj_4776), .I1(n10_adj_4754), .I2(n67241), 
            .I3(n63669), .O(n65971));   // verilog/motorControl.v(62[35:55])
    defparam i48909_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32503_4_lut (.I0(n67502), .I1(\Kp[4] ), .I2(n6_adj_4854), 
            .I3(n207[22]), .O(n8_adj_4941));   // verilog/motorControl.v(61[20:26])
    defparam i32503_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i32456_4_lut (.I0(n20550[1]), .I1(\Kp[3] ), .I2(n59384), .I3(n207[23]), 
            .O(n6_adj_4942));   // verilog/motorControl.v(61[20:26])
    defparam i32456_4_lut.LUT_INIT = 16'he800;
    SB_LUT4 i1_4_lut_adj_949 (.I0(n6_adj_4942), .I1(n8_adj_4941), .I2(n59378), 
            .I3(n55858), .O(n57914));   // verilog/motorControl.v(61[20:26])
    defparam i1_4_lut_adj_949.LUT_INIT = 16'h6996;
    SB_LUT4 mult_24_i592_2_lut (.I0(\Ki[12] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_4594));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i641_2_lut (.I0(\Ki[13] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_4593));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i596_2_lut (.I0(\Ki[12] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886_adj_4700));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i690_2_lut (.I0(\Ki[14] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_4591));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i645_2_lut (.I0(\Ki[13] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959_adj_4699));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i449_2_lut (.I0(\Kp[9] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n667_adj_4698));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i694_2_lut (.I0(\Ki[14] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032_adj_4697));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i498_2_lut (.I0(\Kp[10] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_26_i11_2_lut (.I0(deadband[5]), .I1(n455[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4601));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i13_2_lut (.I0(deadband[6]), .I1(n455[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4600));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i15_2_lut (.I0(deadband[7]), .I1(n455[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4599));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i9_2_lut (.I0(deadband[4]), .I1(n455[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4623));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i17_2_lut (.I0(deadband[8]), .I1(n455[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4625));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i19_2_lut (.I0(deadband[9]), .I1(n455[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4624));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i21_2_lut (.I0(deadband[10]), .I1(n455[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4628));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i23_2_lut (.I0(deadband[11]), .I1(n455[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4627));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i25_2_lut (.I0(deadband[12]), .I1(n455[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4626));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_26_i27_2_lut (.I0(deadband[13]), .I1(n455[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4598));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i9_2_lut (.I0(PWMLimit[4]), .I1(n455[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4943));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i11_2_lut (.I0(PWMLimit[5]), .I1(n455[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4944));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i13_2_lut (.I0(PWMLimit[6]), .I1(n455[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4945));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i15_2_lut (.I0(PWMLimit[7]), .I1(n455[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4946));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i21_2_lut (.I0(PWMLimit[10]), .I1(n455[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_c));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i19_2_lut (.I0(PWMLimit[9]), .I1(n455[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4947));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i17_2_lut (.I0(PWMLimit[8]), .I1(n455[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i23_2_lut (.I0(PWMLimit[11]), .I1(n455[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i25_2_lut (.I0(PWMLimit[12]), .I1(n455[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_c));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i27_2_lut (.I0(PWMLimit[13]), .I1(n455[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i9_2_lut (.I0(setpoint[4]), .I1(n535[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4554));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i11_2_lut (.I0(setpoint[5]), .I1(n535[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4559));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i13_2_lut (.I0(setpoint[6]), .I1(n535[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4558));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i15_2_lut (.I0(setpoint[7]), .I1(n535[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4557));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i21_2_lut (.I0(setpoint[10]), .I1(n535[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4551));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i19_2_lut (.I0(setpoint[9]), .I1(n535[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4552));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i17_2_lut (.I0(setpoint[8]), .I1(n535[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4553));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i23_2_lut (.I0(setpoint[11]), .I1(n535[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4565));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i25_2_lut (.I0(setpoint[12]), .I1(n535[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4564));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_11_i27_2_lut (.I0(setpoint[13]), .I1(n535[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4556));   // verilog/motorControl.v(47[25:43])
    defparam LessThan_11_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i11_2_lut (.I0(n455[5]), .I1(n535[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4651));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i13_2_lut (.I0(n455[6]), .I1(n535[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4650));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i15_2_lut (.I0(n455[7]), .I1(n535[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4649));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i9_2_lut (.I0(n455[4]), .I1(n535[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4659));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i17_2_lut (.I0(n455[8]), .I1(n535[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4661));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i47302_3_lut (.I0(n65630), .I1(n28[15]), .I2(n455[15]), .I3(GND_net), 
            .O(n64364));   // verilog/motorControl.v(62[35:55])
    defparam i47302_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_32_i19_2_lut (.I0(n455[9]), .I1(n535[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4660));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i21_2_lut (.I0(n455[10]), .I1(n535[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4664));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i23_2_lut (.I0(n455[11]), .I1(n535[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4663));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_32_i25_2_lut (.I0(n455[12]), .I1(n535[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4662));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32474_2_lut_3_lut (.I0(\Kp[1] ), .I1(n207[22]), .I2(n68_adj_4903), 
            .I3(GND_net), .O(n20502[0]));   // verilog/motorControl.v(61[20:26])
    defparam i32474_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 mult_24_i739_2_lut (.I0(\Ki[15] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_4588));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut (.I0(\Kp[1] ), .I1(n207[22]), .I2(n68_adj_4903), 
            .I3(n59388), .O(n20502[1]));   // verilog/motorControl.v(61[20:26])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h7f80;
    SB_LUT4 mult_24_i414_2_lut (.I0(\Ki[8] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_4940));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i706_2_lut (.I0(\Kp[14] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n1050_adj_4939));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i463_2_lut (.I0(\Ki[9] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_4938));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i512_2_lut (.I0(\Ki[10] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761_adj_4937));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i85_2_lut (.I0(\Ki[1] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_4936));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i547_2_lut (.I0(\Kp[11] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i38_2_lut (.I0(\Ki[0] ), .I1(n335[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_4935));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i561_2_lut (.I0(\Ki[11] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_4934));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i610_2_lut (.I0(\Ki[12] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_4933));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i659_2_lut (.I0(\Ki[13] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_4932));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i134_2_lut (.I0(\Ki[2] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_4931));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i183_2_lut (.I0(\Ki[3] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_4930));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i81_2_lut (.I0(\Kp[1] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_4929));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i34_2_lut (.I0(\Kp[0] ), .I1(n207[20]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_4928));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i130_2_lut (.I0(\Kp[2] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_4927));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i179_2_lut (.I0(\Kp[3] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_4926));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i232_2_lut (.I0(\Ki[4] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4925));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i228_2_lut (.I0(\Kp[4] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_4924));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i281_2_lut (.I0(\Ki[5] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_4923));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_950 (.I0(n20538[2]), .I1(n6_adj_4949), .I2(\Ki[4] ), 
            .I3(n335[18]), .O(n20481[3]));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_950.LUT_INIT = 16'h9666;
    SB_LUT4 mux_21_i15_3_lut (.I0(n233[14]), .I1(n285[14]), .I2(n284), 
            .I3(GND_net), .O(n310[14]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i15_3_lut (.I0(n310[14]), .I1(IntegralLimit[14]), .I2(n258), 
            .I3(GND_net), .O(n335[14]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i77_2_lut (.I0(\Ki[1] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i30_2_lut (.I0(\Ki[0] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i126_2_lut (.I0(\Ki[2] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49120_4_lut (.I0(n64364), .I1(n65971), .I2(n67241), .I3(n63677), 
            .O(n66182));   // verilog/motorControl.v(62[35:55])
    defparam i49120_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_32_i4_4_lut (.I0(n455[0]), .I1(n535[1]), .I2(n455[1]), 
            .I3(n535[0]), .O(n4_adj_4951));   // verilog/motorControl.v(65[25:41])
    defparam LessThan_32_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i48115_3_lut (.I0(n4_adj_4951), .I1(n535[13]), .I2(n27_adj_4642), 
            .I3(GND_net), .O(n65177));   // verilog/motorControl.v(65[25:41])
    defparam i48115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49121_3_lut (.I0(n66182), .I1(n28[18]), .I2(n455[18]), .I3(GND_net), 
            .O(n66183));   // verilog/motorControl.v(62[35:55])
    defparam i49121_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48116_3_lut (.I0(n65177), .I1(n535[14]), .I2(n29_adj_4643), 
            .I3(GND_net), .O(n65178));   // verilog/motorControl.v(65[25:41])
    defparam i48116_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_951 (.I0(n20596[0]), .I1(n47985), .I2(\Ki[2] ), 
            .I3(n335[20]), .O(n20575[1]));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_951.LUT_INIT = 16'h9666;
    SB_LUT4 i49081_3_lut (.I0(n66183), .I1(n28[19]), .I2(n455[19]), .I3(GND_net), 
            .O(n66143));   // verilog/motorControl.v(62[35:55])
    defparam i49081_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_24_i330_2_lut (.I0(\Ki[6] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_4922));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_952 (.I0(\Ki[1] ), .I1(\Ki[0] ), .I2(n335[22]), 
            .I3(n335[23]), .O(n59342));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_952.LUT_INIT = 16'h93a0;
    SB_LUT4 i1_4_lut_adj_953 (.I0(\Ki[5] ), .I1(\Ki[4] ), .I2(n335[18]), 
            .I3(n335[19]), .O(n59346));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_953.LUT_INIT = 16'h6ca0;
    SB_LUT4 i1_4_lut_adj_954 (.I0(\Ki[3] ), .I1(\Ki[2] ), .I2(n335[20]), 
            .I3(n335[21]), .O(n59344));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_954.LUT_INIT = 16'h6ca0;
    SB_LUT4 i46430_4_lut (.I0(n33_adj_4641), .I1(n31_adj_4640), .I2(n29_adj_4643), 
            .I3(n63510), .O(n63492));
    defparam i46430_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i1_4_lut_adj_955 (.I0(n59344), .I1(n47955), .I2(n59346), .I3(n59342), 
            .O(n59352));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_955.LUT_INIT = 16'h6996;
    SB_LUT4 i32285_4_lut (.I0(n20596[0]), .I1(\Ki[2] ), .I2(n47985), .I3(n335[20]), 
            .O(n4_adj_4953));   // verilog/motorControl.v(61[29:40])
    defparam i32285_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 mult_23_i73_2_lut (.I0(\Kp[1] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_4585));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32423_4_lut (.I0(n20538[2]), .I1(\Ki[4] ), .I2(n6_adj_4949), 
            .I3(n335[18]), .O(n8_adj_4954));   // verilog/motorControl.v(61[29:40])
    defparam i32423_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_956 (.I0(n6_adj_4955), .I1(n8_adj_4954), .I2(n4_adj_4953), 
            .I3(n59352), .O(n57863));   // verilog/motorControl.v(61[29:40])
    defparam i1_4_lut_adj_956.LUT_INIT = 16'h6996;
    SB_LUT4 LessThan_28_i6_3_lut (.I0(n28[2]), .I1(n28[3]), .I2(n455[3]), 
            .I3(GND_net), .O(n6_adj_4956));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_23_i26_2_lut (.I0(\Kp[0] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_4584));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i277_2_lut (.I0(\Kp[5] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_4921));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i175_2_lut (.I0(\Ki[3] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i326_2_lut (.I0(\Kp[6] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_4920));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i122_2_lut (.I0(\Kp[2] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_4583));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i67_2_lut (.I0(\Kp[1] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_4919));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i20_2_lut (.I0(\Kp[0] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4918));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i375_2_lut (.I0(\Kp[7] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_4917));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i171_2_lut (.I0(\Kp[3] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_4582));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i424_2_lut (.I0(\Kp[8] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_4916));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i116_2_lut (.I0(\Kp[2] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4915));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i224_2_lut (.I0(\Ki[4] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i273_2_lut (.I0(\Ki[5] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i69_2_lut (.I0(\Ki[1] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_4914));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i22_2_lut (.I0(\Ki[0] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_4913));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i118_2_lut (.I0(\Ki[2] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174_adj_4912));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i165_2_lut (.I0(\Kp[3] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4911));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i167_2_lut (.I0(\Ki[3] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_4910));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i214_2_lut (.I0(\Kp[4] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4909));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i220_2_lut (.I0(\Kp[4] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_4581));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i216_2_lut (.I0(\Ki[4] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_4908));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i265_2_lut (.I0(\Ki[5] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_4907));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i314_2_lut (.I0(\Ki[6] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_4906));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i263_2_lut (.I0(\Kp[5] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4905));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i363_2_lut (.I0(\Ki[7] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_4904));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i312_2_lut (.I0(\Kp[6] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_4902));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i361_2_lut (.I0(\Kp[7] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4901));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i412_2_lut (.I0(\Ki[8] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_4900));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i410_2_lut (.I0(\Kp[8] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_4899));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i459_2_lut (.I0(\Kp[9] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_4898));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i461_2_lut (.I0(\Ki[9] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_4897));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i743_2_lut (.I0(\Ki[15] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105_adj_4696));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i510_2_lut (.I0(\Ki[10] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_4896));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i508_2_lut (.I0(\Kp[10] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_4895));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46515_2_lut_4_lut (.I0(PWMLimit[16]), .I1(n455[16]), .I2(PWMLimit[7]), 
            .I3(n455[7]), .O(n63577));
    defparam i46515_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i557_2_lut (.I0(\Kp[11] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_4894));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i559_2_lut (.I0(\Ki[11] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831_adj_4893));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i596_2_lut (.I0(\Kp[12] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i608_2_lut (.I0(\Ki[12] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904_adj_4891));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i606_2_lut (.I0(\Kp[12] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_4890));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i269_2_lut (.I0(\Kp[5] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_4576));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i657_2_lut (.I0(\Ki[13] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977_adj_4889));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i706_2_lut (.I0(\Ki[14] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i655_2_lut (.I0(\Kp[13] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_4888));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i704_2_lut (.I0(\Kp[14] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_4887));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i318_2_lut (.I0(\Kp[6] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_4575));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i753_2_lut (.I0(\Kp[15] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_4886));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i367_2_lut (.I0(\Kp[7] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_4574));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i416_2_lut (.I0(\Kp[8] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_4573));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i465_2_lut (.I0(\Kp[9] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_4572));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i67_2_lut (.I0(\Ki[1] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i20_2_lut (.I0(\Ki[0] ), .I1(n335[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4885));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i514_2_lut (.I0(\Kp[10] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_4571));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i116_2_lut (.I0(\Ki[2] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i65_2_lut (.I0(\Kp[1] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_4884));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i18_2_lut (.I0(\Kp[0] ), .I1(n207[12]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4883));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i322_2_lut (.I0(\Ki[6] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4570));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i165_2_lut (.I0(\Ki[3] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4882));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i6_3_lut_3_lut (.I0(setpoint[2]), .I1(setpoint[3]), 
            .I2(PWMLimit[3]), .I3(GND_net), .O(n6_adj_4957));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_23_i114_2_lut (.I0(\Kp[2] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n168_adj_4881));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i163_2_lut (.I0(\Kp[3] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4880));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46177_2_lut_4_lut (.I0(PWMLimit[8]), .I1(setpoint[8]), .I2(PWMLimit[4]), 
            .I3(setpoint[4]), .O(n63239));
    defparam i46177_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i214_2_lut (.I0(\Ki[4] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i8_3_lut_3_lut (.I0(setpoint[4]), .I1(setpoint[8]), 
            .I2(PWMLimit[8]), .I3(GND_net), .O(n8_adj_4958));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_24_i263_2_lut (.I0(\Ki[5] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4879));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_9_i10_3_lut_3_lut (.I0(setpoint[5]), .I1(setpoint[6]), 
            .I2(PWMLimit[6]), .I3(GND_net), .O(n10_adj_4959));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48569_3_lut (.I0(n6_adj_4956), .I1(n28[10]), .I2(n455[10]), 
            .I3(GND_net), .O(n65631));   // verilog/motorControl.v(62[35:55])
    defparam i48569_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_23_i563_2_lut (.I0(\Kp[11] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_4569));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i212_2_lut (.I0(\Kp[4] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_4878));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i371_2_lut (.I0(\Ki[7] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4568));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i312_2_lut (.I0(\Ki[6] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_4877));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[0]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[1]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i361_2_lut (.I0(\Ki[7] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4874));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i261_2_lut (.I0(\Kp[5] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4873));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[2]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i410_2_lut (.I0(\Ki[8] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[3]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[4]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i48803_4_lut (.I0(n30_adj_4658), .I1(n10_adj_4657), .I2(n35_adj_4637), 
            .I3(n63488), .O(n65865));   // verilog/motorControl.v(65[25:41])
    defparam i48803_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_24_i459_2_lut (.I0(\Ki[9] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i310_2_lut (.I0(\Kp[6] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4869));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[5]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i46197_2_lut_4_lut (.I0(PWMLimit[6]), .I1(setpoint[6]), .I2(PWMLimit[5]), 
            .I3(setpoint[5]), .O(n63259));
    defparam i46197_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i612_2_lut (.I0(\Kp[12] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_4567));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[6]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i508_2_lut (.I0(\Ki[10] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i359_2_lut (.I0(\Kp[7] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n533_adj_4866));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48570_3_lut (.I0(n65631), .I1(n28[11]), .I2(n455[11]), .I3(GND_net), 
            .O(n65632));   // verilog/motorControl.v(62[35:55])
    defparam i48570_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_20_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[7]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[8]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i557_2_lut (.I0(\Ki[11] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i408_2_lut (.I0(\Kp[8] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n606_adj_4863));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i606_2_lut (.I0(\Ki[12] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[9]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i655_2_lut (.I0(\Ki[13] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[10]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i704_2_lut (.I0(\Ki[14] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[11]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i753_2_lut (.I0(\Ki[15] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i457_2_lut (.I0(\Kp[9] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_4859));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[12]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[13]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[14]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i506_2_lut (.I0(\Kp[10] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_4855));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[15]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i555_2_lut (.I0(\Kp[11] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_4852));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[16]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[17]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[18]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i47322_3_lut (.I0(n65178), .I1(n535[15]), .I2(n31_adj_4640), 
            .I3(GND_net), .O(n64384));   // verilog/motorControl.v(65[25:41])
    defparam i47322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_20_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[19]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i604_2_lut (.I0(\Kp[12] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n898_adj_4846));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[20]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[21]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i653_2_lut (.I0(\Kp[13] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n971_adj_4843));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i75_2_lut (.I0(\Kp[1] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_4842));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i28_2_lut (.I0(\Kp[0] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4841));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i702_2_lut (.I0(\Kp[14] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1044_adj_4840));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i124_2_lut (.I0(\Kp[2] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_4839));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_20_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[22]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_20_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4994[23]));   // verilog/motorControl.v(59[24:38])
    defparam unary_minus_20_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22927_1_lut (.I0(n455[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38672));   // verilog/motorControl.v(61[20:40])
    defparam i22927_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i1_1_lut (.I0(deadband[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[0]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i751_2_lut (.I0(\Kp[15] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_4835));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i2_1_lut (.I0(deadband[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[1]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i173_2_lut (.I0(\Kp[3] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4833));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i83_2_lut (.I0(\Ki[1] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_4832));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i36_2_lut (.I0(\Ki[0] ), .I1(n335[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_4831));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i222_2_lut (.I0(\Kp[4] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_4830));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i271_2_lut (.I0(\Kp[5] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_4829));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i3_1_lut (.I0(deadband[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[2]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i79_2_lut (.I0(\Kp[1] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4827));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i32_2_lut (.I0(\Kp[0] ), .I1(n207[19]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4826));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i132_2_lut (.I0(\Ki[2] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_4825));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i4_1_lut (.I0(deadband[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[3]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i5_1_lut (.I0(deadband[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[4]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i128_2_lut (.I0(\Kp[2] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4821));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i320_2_lut (.I0(\Kp[6] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4820));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i369_2_lut (.I0(\Kp[7] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_4819));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i181_2_lut (.I0(\Ki[3] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4818));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i6_1_lut (.I0(deadband[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[5]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i177_2_lut (.I0(\Kp[3] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4816));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i7_1_lut (.I0(deadband[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[6]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i226_2_lut (.I0(\Kp[4] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_4814));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i71_2_lut (.I0(\Kp[1] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_4457));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i230_2_lut (.I0(\Ki[4] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_4813));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i24_2_lut (.I0(\Kp[0] ), .I1(n207[15]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4456));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i418_2_lut (.I0(\Kp[8] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_4812));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i8_1_lut (.I0(deadband[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[7]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i645_2_lut (.I0(\Kp[13] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i9_1_lut (.I0(deadband[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[8]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i279_2_lut (.I0(\Ki[5] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_4809));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i10_1_lut (.I0(deadband[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[9]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i275_2_lut (.I0(\Kp[5] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_4807));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i328_2_lut (.I0(\Ki[6] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_4806));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i11_1_lut (.I0(deadband[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[10]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i12_1_lut (.I0(deadband[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[11]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i324_2_lut (.I0(\Kp[6] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_4803));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i377_2_lut (.I0(\Ki[7] ), .I1(n335[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_4802));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i13_1_lut (.I0(deadband[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[12]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i14_1_lut (.I0(deadband[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[13]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i373_2_lut (.I0(\Kp[7] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4799));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i15_1_lut (.I0(deadband[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[14]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_27_inv_0_i16_1_lut (.I0(deadband[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[15]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i422_2_lut (.I0(\Kp[8] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_4796));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i63_2_lut (.I0(\Kp[1] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n92_adj_4795));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i16_2_lut (.I0(\Kp[0] ), .I1(n207[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4794));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46587_4_lut (.I0(n455[21]), .I1(n67230), .I2(n28[21]), .I3(n64666), 
            .O(n63649));
    defparam i46587_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 unary_minus_27_inv_0_i17_1_lut (.I0(deadband[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[16]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i471_2_lut (.I0(\Kp[9] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_4792));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i18_1_lut (.I0(deadband[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[17]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i694_2_lut (.I0(\Kp[14] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i19_1_lut (.I0(deadband[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[18]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i65_2_lut (.I0(\Ki[1] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i18_2_lut (.I0(\Ki[0] ), .I1(n335[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i20_1_lut (.I0(deadband[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[19]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i112_2_lut (.I0(\Kp[2] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n165_adj_4788));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i21_1_lut (.I0(deadband[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[20]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i114_2_lut (.I0(\Ki[2] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i22_1_lut (.I0(deadband[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[21]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i163_2_lut (.I0(\Ki[3] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4785));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i467_2_lut (.I0(\Kp[9] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_4784));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i23_1_lut (.I0(deadband[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[22]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i49030_4_lut (.I0(n64384), .I1(n65865), .I2(n35_adj_4637), 
            .I3(n63492), .O(n66092));   // verilog/motorControl.v(65[25:41])
    defparam i49030_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_23_i743_2_lut (.I0(\Kp[15] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i212_2_lut (.I0(\Ki[4] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i77_2_lut (.I0(\Kp[1] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_4695));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i420_2_lut (.I0(\Ki[8] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i161_2_lut (.I0(\Kp[3] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4782));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_27_inv_0_i24_1_lut (.I0(deadband[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4993[23]));   // verilog/motorControl.v(62[45:54])
    defparam unary_minus_27_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[0]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i261_2_lut (.I0(\Ki[5] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4778));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[1]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i310_2_lut (.I0(\Ki[6] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4775));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i120_2_lut (.I0(\Kp[2] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_4455));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i30_2_lut (.I0(\Kp[0] ), .I1(n207[18]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_4694));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i210_2_lut (.I0(\Kp[4] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_4774));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i126_2_lut (.I0(\Kp[2] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4693));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i516_2_lut (.I0(\Kp[10] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_4773));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i259_2_lut (.I0(\Kp[5] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4772));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[2]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i359_2_lut (.I0(\Ki[7] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[3]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[4]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i49031_3_lut (.I0(n66092), .I1(n535[18]), .I2(n37_adj_4633), 
            .I3(GND_net), .O(n66093));   // verilog/motorControl.v(65[25:41])
    defparam i49031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i408_2_lut (.I0(\Ki[8] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i169_2_lut (.I0(\Kp[3] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_4454));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[5]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i308_2_lut (.I0(\Kp[6] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4768));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[6]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i457_2_lut (.I0(\Ki[9] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i175_2_lut (.I0(\Kp[3] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_4692));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[7]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i357_2_lut (.I0(\Kp[7] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n530_adj_4766));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i565_2_lut (.I0(\Kp[11] ), .I1(n207[16]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_4765));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[8]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i506_2_lut (.I0(\Ki[10] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i406_2_lut (.I0(\Kp[8] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n603_adj_4763));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i555_2_lut (.I0(\Ki[11] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i604_2_lut (.I0(\Ki[12] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i218_2_lut (.I0(\Kp[4] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_4453));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i653_2_lut (.I0(\Ki[13] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i267_2_lut (.I0(\Kp[5] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_4452));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i455_2_lut (.I0(\Kp[9] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_4762));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i702_2_lut (.I0(\Ki[14] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[9]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i504_2_lut (.I0(\Kp[10] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_4760));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i751_2_lut (.I0(\Ki[15] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i553_2_lut (.I0(\Kp[11] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_4759));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[10]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i63_2_lut (.I0(\Ki[1] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i16_2_lut (.I0(\Ki[0] ), .I1(n335[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4757));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i112_2_lut (.I0(\Ki[2] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i602_2_lut (.I0(\Kp[12] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_4756));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i161_2_lut (.I0(\Ki[3] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4755));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i224_2_lut (.I0(\Kp[4] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_4691));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i210_2_lut (.I0(\Ki[4] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_4753));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i651_2_lut (.I0(\Kp[13] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_4752));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i259_2_lut (.I0(\Ki[5] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4751));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i308_2_lut (.I0(\Ki[6] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4750));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i700_2_lut (.I0(\Kp[14] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1041_adj_4749));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i357_2_lut (.I0(\Ki[7] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i406_2_lut (.I0(\Ki[8] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i455_2_lut (.I0(\Ki[9] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i749_2_lut (.I0(\Kp[15] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n1114_adj_4748));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i504_2_lut (.I0(\Ki[10] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i553_2_lut (.I0(\Ki[11] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i602_2_lut (.I0(\Ki[12] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i651_2_lut (.I0(\Ki[13] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i61_2_lut (.I0(\Kp[1] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n89_adj_4747));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i14_2_lut (.I0(\Kp[0] ), .I1(n207[10]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4746));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i700_2_lut (.I0(\Ki[14] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i749_2_lut (.I0(\Ki[15] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i110_2_lut (.I0(\Kp[2] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n162_adj_4745));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[11]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i159_2_lut (.I0(\Kp[3] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_4743));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i61_2_lut (.I0(\Ki[1] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i14_2_lut (.I0(\Ki[0] ), .I1(n335[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i110_2_lut (.I0(\Ki[2] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i159_2_lut (.I0(\Ki[3] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_4742));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i208_2_lut (.I0(\Kp[4] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_4741));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i208_2_lut (.I0(\Ki[4] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_4740));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i257_2_lut (.I0(\Kp[5] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n381_adj_4739));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48416_4_lut (.I0(n24_adj_4512), .I1(n8_adj_4511), .I2(n67204), 
            .I3(n63646), .O(n65478));   // verilog/motorControl.v(62[35:55])
    defparam i48416_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_23_i273_2_lut (.I0(\Kp[5] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n405_adj_4690));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i257_2_lut (.I0(\Ki[5] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i322_2_lut (.I0(\Kp[6] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4689));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i306_2_lut (.I0(\Ki[6] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_4738));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i306_2_lut (.I0(\Kp[6] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[12]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i355_2_lut (.I0(\Kp[7] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n527_adj_4736));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i355_2_lut (.I0(\Ki[7] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i404_2_lut (.I0(\Kp[8] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n600_adj_4735));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i453_2_lut (.I0(\Kp[9] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n673_adj_4734));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i404_2_lut (.I0(\Ki[8] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i371_2_lut (.I0(\Kp[7] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4688));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i502_2_lut (.I0(\Kp[10] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_4733));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[13]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i453_2_lut (.I0(\Ki[9] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i551_2_lut (.I0(\Kp[11] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_4731));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i420_2_lut (.I0(\Kp[8] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_4687));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[14]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i502_2_lut (.I0(\Ki[10] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i551_2_lut (.I0(\Ki[11] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i469_2_lut (.I0(\Kp[9] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_4686));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i600_2_lut (.I0(\Kp[12] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_4729));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[15]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i600_2_lut (.I0(\Ki[12] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i649_2_lut (.I0(\Ki[13] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_4727));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i649_2_lut (.I0(\Kp[13] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i518_2_lut (.I0(\Kp[10] ), .I1(n207[17]), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_4685));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i55_2_lut (.I0(\Kp[1] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_4684));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i47300_3_lut (.I0(n65632), .I1(n28[12]), .I2(n455[12]), .I3(GND_net), 
            .O(n64362));   // verilog/motorControl.v(62[35:55])
    defparam i47300_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_23_i8_2_lut (.I0(\Kp[0] ), .I1(n207[7]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4683));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i698_2_lut (.I0(\Ki[14] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038_adj_4726));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i747_2_lut (.I0(\Ki[15] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111_adj_4725));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i4_3_lut (.I0(n233[3]), .I1(n285[3]), .I2(n284), .I3(GND_net), 
            .O(n310[3]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i4_3_lut (.I0(n310[3]), .I1(IntegralLimit[3]), .I2(n258), 
            .I3(GND_net), .O(n335[3]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i55_2_lut (.I0(\Ki[1] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i49001_3_lut (.I0(n66093), .I1(n535[19]), .I2(n39_adj_4639), 
            .I3(GND_net), .O(n66063));   // verilog/motorControl.v(65[25:41])
    defparam i49001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i8_2_lut (.I0(\Ki[0] ), .I1(n335[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4682));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i698_2_lut (.I0(\Kp[14] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i747_2_lut (.I0(\Kp[15] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[16]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i59_2_lut (.I0(\Kp[1] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_4722));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i12_2_lut (.I0(\Kp[0] ), .I1(n207[9]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4721));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[17]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i104_2_lut (.I0(\Kp[2] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4681));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i108_2_lut (.I0(\Kp[2] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n159_adj_4719));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i104_2_lut (.I0(\Ki[2] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i153_2_lut (.I0(\Kp[3] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4680));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i202_2_lut (.I0(\Kp[4] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4679));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i251_2_lut (.I0(\Kp[5] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n372_adj_4678));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i153_2_lut (.I0(\Ki[3] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4677));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i202_2_lut (.I0(\Ki[4] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299_adj_4676));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i300_2_lut (.I0(\Kp[6] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4675));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i157_2_lut (.I0(\Kp[3] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n232_adj_4718));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i349_2_lut (.I0(\Kp[7] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n518_adj_4674));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i398_2_lut (.I0(\Kp[8] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n591_adj_4673));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[18]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_33_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[19]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i251_2_lut (.I0(\Ki[5] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i206_2_lut (.I0(\Kp[4] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n305_adj_4716));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i300_2_lut (.I0(\Ki[6] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445_adj_4672));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i349_2_lut (.I0(\Ki[7] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[20]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i46414_4_lut (.I0(n43_adj_4636), .I1(n41_adj_4635), .I2(n39_adj_4639), 
            .I3(n66047), .O(n63476));
    defparam i46414_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_23_i447_2_lut (.I0(\Kp[9] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n664_adj_4671));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i496_2_lut (.I0(\Kp[10] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_4670));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i398_2_lut (.I0(\Ki[8] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i255_2_lut (.I0(\Kp[5] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n378_adj_4714));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i545_2_lut (.I0(\Kp[11] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n810_adj_4669));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46589_4_lut (.I0(n455[21]), .I1(n67206), .I2(n28[21]), .I3(n66154), 
            .O(n63651));
    defparam i46589_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_24_i469_2_lut (.I0(\Ki[9] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i447_2_lut (.I0(\Ki[9] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i496_2_lut (.I0(\Ki[10] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i518_2_lut (.I0(\Ki[10] ), .I1(n335[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i594_2_lut (.I0(\Kp[12] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n883_adj_4668));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i545_2_lut (.I0(\Ki[11] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i643_2_lut (.I0(\Kp[13] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n956_adj_4667));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i594_2_lut (.I0(\Ki[12] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[21]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i2_2_lut (.I0(\Ki[0] ), .I1(n335[0]), .I2(GND_net), 
            .I3(GND_net), .O(n34[0]));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i2_2_lut (.I0(\Kp[0] ), .I1(n207[4]), .I2(GND_net), 
            .I3(GND_net), .O(n360[0]));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[22]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_23_i304_2_lut (.I0(\Kp[6] ), .I1(n207[8]), .I2(GND_net), 
            .I3(GND_net), .O(n451_adj_4711));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_33_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4992[23]));   // verilog/motorControl.v(66[24:33])
    defparam unary_minus_33_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i59_2_lut (.I0(\Ki[1] ), .I1(n335[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i12_2_lut (.I0(\Ki[0] ), .I1(n335[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4710));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22914_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n38659));   // verilog/motorControl.v(42[14] 73[8])
    defparam i22914_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_24_i643_2_lut (.I0(\Ki[13] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i692_2_lut (.I0(\Kp[14] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1029_adj_4666));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i692_2_lut (.I0(\Ki[14] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i741_2_lut (.I0(\Kp[15] ), .I1(n207[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1102_adj_4656));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i741_2_lut (.I0(\Ki[15] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_28_i45_rep_58_2_lut (.I0(n455[22]), .I1(n28[22]), .I2(GND_net), 
            .I3(GND_net), .O(n67204));   // verilog/motorControl.v(62[35:55])
    defparam LessThan_28_i45_rep_58_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_21_i16_3_lut (.I0(n233[15]), .I1(n285[15]), .I2(n284), 
            .I3(GND_net), .O(n310[15]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i16_3_lut (.I0(n310[15]), .I1(IntegralLimit[15]), .I2(n258), 
            .I3(GND_net), .O(n335[15]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i23_3_lut (.I0(n233[22]), .I1(n285[22]), .I2(n284), 
            .I3(GND_net), .O(n310[22]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i23_3_lut (.I0(n310[22]), .I1(IntegralLimit[22]), .I2(n258), 
            .I3(GND_net), .O(n335[22]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i22_3_lut (.I0(n233[21]), .I1(n285[21]), .I2(n284), 
            .I3(GND_net), .O(n310[21]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i22_3_lut (.I0(n310[21]), .I1(IntegralLimit[21]), .I2(n258), 
            .I3(GND_net), .O(n335[21]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i79_2_lut (.I0(\Ki[1] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i21_3_lut (.I0(n233[20]), .I1(n285[20]), .I2(n284), 
            .I3(GND_net), .O(n310[20]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i21_3_lut (.I0(n310[20]), .I1(IntegralLimit[20]), .I2(n258), 
            .I3(GND_net), .O(n335[20]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i20_3_lut (.I0(n233[19]), .I1(n285[19]), .I2(n284), 
            .I3(GND_net), .O(n310[19]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i20_3_lut (.I0(n310[19]), .I1(IntegralLimit[19]), .I2(n258), 
            .I3(GND_net), .O(n335[19]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i19_3_lut (.I0(n233[18]), .I1(n285[18]), .I2(n284), 
            .I3(GND_net), .O(n310[18]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i19_3_lut (.I0(n310[18]), .I1(IntegralLimit[18]), .I2(n258), 
            .I3(GND_net), .O(n335[18]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i32_2_lut (.I0(\Ki[0] ), .I1(n335[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i18_3_lut (.I0(n233[17]), .I1(n285[17]), .I2(n284), 
            .I3(GND_net), .O(n310[17]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i18_3_lut (.I0(n310[17]), .I1(IntegralLimit[17]), .I2(n258), 
            .I3(GND_net), .O(n335[17]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i128_2_lut (.I0(\Ki[2] ), .I1(n335[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i3_3_lut (.I0(n233[2]), .I1(n285[2]), .I2(n284), .I3(GND_net), 
            .O(n310[2]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i3_3_lut (.I0(n310[2]), .I1(IntegralLimit[2]), .I2(n258), 
            .I3(GND_net), .O(n335[2]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i53_2_lut (.I0(\Ki[1] ), .I1(n335[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_4648));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i10_3_lut (.I0(n233[9]), .I1(n285[9]), .I2(n284), .I3(GND_net), 
            .O(n310[9]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i6_2_lut (.I0(\Ki[0] ), .I1(n335[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4647));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_22_i10_3_lut (.I0(n310[9]), .I1(IntegralLimit[9]), .I2(n258), 
            .I3(GND_net), .O(n335[9]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i9_3_lut (.I0(n233[8]), .I1(n285[8]), .I2(n284), .I3(GND_net), 
            .O(n310[8]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i9_3_lut (.I0(n310[8]), .I1(IntegralLimit[8]), .I2(n258), 
            .I3(GND_net), .O(n335[8]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i8_3_lut (.I0(n233[7]), .I1(n285[7]), .I2(n284), .I3(GND_net), 
            .O(n310[7]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i8_3_lut (.I0(n310[7]), .I1(IntegralLimit[7]), .I2(n258), 
            .I3(GND_net), .O(n335[7]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i7_3_lut (.I0(n233[6]), .I1(n285[6]), .I2(n284), .I3(GND_net), 
            .O(n310[6]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i7_3_lut (.I0(n310[6]), .I1(IntegralLimit[6]), .I2(n258), 
            .I3(GND_net), .O(n335[6]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_21_i6_3_lut (.I0(n233[5]), .I1(n285[5]), .I2(n284), .I3(GND_net), 
            .O(n310[5]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i6_3_lut (.I0(n310[5]), .I1(IntegralLimit[5]), .I2(n258), 
            .I3(GND_net), .O(n335[5]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n9972_bdd_4_lut_49865 (.I0(n9972), .I1(n63132), .I2(setpoint[23]), 
            .I3(n4744), .O(n66849));
    defparam n9972_bdd_4_lut_49865.LUT_INIT = 16'he4aa;
    SB_LUT4 n66849_bdd_4_lut (.I0(n66849), .I1(n535[23]), .I2(n455[23]), 
            .I3(n4744), .O(n66852));
    defparam n66849_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i48747_4_lut (.I0(n64382), .I1(n65482), .I2(n45_adj_4634), 
            .I3(n63474), .O(n65809));   // verilog/motorControl.v(65[25:41])
    defparam i48747_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48971_4_lut (.I0(n64362), .I1(n65478), .I2(n67204), .I3(n63649), 
            .O(n66033));   // verilog/motorControl.v(62[35:55])
    defparam i48971_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i47328_3_lut (.I0(n66063), .I1(n535[20]), .I2(n41_adj_4635), 
            .I3(GND_net), .O(n64390));   // verilog/motorControl.v(65[25:41])
    defparam i47328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47308_3_lut (.I0(n66143), .I1(n28[20]), .I2(n455[20]), .I3(GND_net), 
            .O(n64370));   // verilog/motorControl.v(62[35:55])
    defparam i47308_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48973_4_lut (.I0(n64370), .I1(n66033), .I2(n67204), .I3(n63651), 
            .O(n66035));   // verilog/motorControl.v(62[35:55])
    defparam i48973_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_26_i4_4_lut (.I0(deadband[0]), .I1(n455[1]), .I2(deadband[1]), 
            .I3(n455[0]), .O(n4_adj_4965));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i48573_3_lut (.I0(n4_adj_4965), .I1(n455[13]), .I2(n27_adj_4598), 
            .I3(GND_net), .O(n65635));   // verilog/motorControl.v(62[14:31])
    defparam i48573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48977_4_lut (.I0(n64390), .I1(n65809), .I2(n45_adj_4634), 
            .I3(n63476), .O(n66039));   // verilog/motorControl.v(65[25:41])
    defparam i48977_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48574_3_lut (.I0(n65635), .I1(n455[14]), .I2(n29), .I3(GND_net), 
            .O(n65636));   // verilog/motorControl.v(62[14:31])
    defparam i48574_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut (.I0(n66039), .I1(n4_adj_4966), .I2(n455[23]), .I3(n535[23]), 
            .O(n57934));
    defparam i2_4_lut.LUT_INIT = 16'hdfcd;
    SB_LUT4 i1_2_lut_4_lut (.I0(n66019), .I1(setpoint[23]), .I2(n535[23]), 
            .I3(n25015), .O(n7062));   // verilog/motorControl.v(47[25:43])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h7100;
    SB_LUT4 i46699_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n63783), 
            .O(n63761));
    defparam i46699_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48907_4_lut (.I0(n30_adj_4614), .I1(n10_adj_4613), .I2(n35), 
            .I3(n63757), .O(n65969));   // verilog/motorControl.v(62[14:31])
    defparam i48907_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_2_lut_4_lut_adj_957 (.I0(n66019), .I1(setpoint[23]), .I2(n535[23]), 
            .I3(n25015), .O(n25017));   // verilog/motorControl.v(47[25:43])
    defparam i1_2_lut_4_lut_adj_957.LUT_INIT = 16'h8e00;
    SB_LUT4 i4428_4_lut (.I0(n7062), .I1(n4744), .I2(n57934), .I3(n25017), 
            .O(n9972));
    defparam i4428_4_lut.LUT_INIT = 16'hbbab;
    SB_LUT4 i47292_3_lut (.I0(n65636), .I1(n455[15]), .I2(n31), .I3(GND_net), 
            .O(n64354));   // verilog/motorControl.v(62[14:31])
    defparam i47292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49118_4_lut (.I0(n64354), .I1(n65969), .I2(n35), .I3(n63761), 
            .O(n66180));   // verilog/motorControl.v(62[14:31])
    defparam i49118_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i49119_3_lut (.I0(n66180), .I1(n455[18]), .I2(n37), .I3(GND_net), 
            .O(n66181));   // verilog/motorControl.v(62[14:31])
    defparam i49119_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46250_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[13]), 
            .I3(GND_net), .O(n62945));
    defparam i46250_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i49083_3_lut (.I0(n66181), .I1(n455[19]), .I2(n39_adj_4708), 
            .I3(GND_net), .O(n66145));   // verilog/motorControl.v(62[14:31])
    defparam i49083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46183_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[14]), 
            .I3(GND_net), .O(n63019));
    defparam i46183_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i46675_4_lut (.I0(n43), .I1(n41_adj_4967), .I2(n39_adj_4708), 
            .I3(n66074), .O(n63737));
    defparam i46675_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46420_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[15]), 
            .I3(GND_net), .O(n63054));
    defparam i46420_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i48967_4_lut (.I0(n64352), .I1(n65476), .I2(n45_adj_4654), 
            .I3(n63724), .O(n66029));   // verilog/motorControl.v(62[14:31])
    defparam i48967_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i46506_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[23]), 
            .I3(GND_net), .O(n63132));
    defparam i46506_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i46368_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[9]), 
            .I3(GND_net), .O(n63175));
    defparam i46368_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i46367_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[10]), 
            .I3(GND_net), .O(n63176));
    defparam i46367_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i46383_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[11]), 
            .I3(GND_net), .O(n63177));
    defparam i46383_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i46366_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[12]), 
            .I3(GND_net), .O(n63178));
    defparam i46366_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i46357_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[16]), 
            .I3(GND_net), .O(n63055));
    defparam i46357_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i46133_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[17]), 
            .I3(GND_net), .O(n63111));
    defparam i46133_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i46470_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[18]), 
            .I3(GND_net), .O(n63114));
    defparam i46470_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i47106_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[6]), 
            .I3(GND_net), .O(n63172));
    defparam i47106_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i46370_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[7]), 
            .I3(GND_net), .O(n63173));
    defparam i46370_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i46906_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[4]), 
            .I3(GND_net), .O(n63167));
    defparam i46906_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i46461_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[3]), 
            .I3(GND_net), .O(n63160));
    defparam i46461_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i47003_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[2]), 
            .I3(GND_net), .O(n63142));
    defparam i47003_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i46353_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[22]), 
            .I3(GND_net), .O(n63118));
    defparam i46353_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i46222_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[1]), 
            .I3(GND_net), .O(n63140));
    defparam i46222_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i46363_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[19]), 
            .I3(GND_net), .O(n63115));
    defparam i46363_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i46354_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[20]), 
            .I3(GND_net), .O(n63116));
    defparam i46354_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i46362_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n63117));
    defparam i46362_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i46967_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[0]), 
            .I3(GND_net), .O(n63139));
    defparam i46967_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i46369_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[8]), 
            .I3(GND_net), .O(n63174));
    defparam i46369_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i1_2_lut_4_lut_adj_958 (.I0(n66037), .I1(PWMLimit[23]), .I2(n455[23]), 
            .I3(n24981), .O(n24983));   // verilog/motorControl.v(63[16:31])
    defparam i1_2_lut_4_lut_adj_958.LUT_INIT = 16'hff71;
    SB_LUT4 i46372_2_lut_3_lut (.I0(n7064), .I1(n24983), .I2(PWMLimit[5]), 
            .I3(GND_net), .O(n63168));
    defparam i46372_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 n9972_bdd_4_lut_49592 (.I0(n9972), .I1(n63054), .I2(setpoint[15]), 
            .I3(n4744), .O(n66663));
    defparam n9972_bdd_4_lut_49592.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_959 (.I0(n66037), .I1(PWMLimit[23]), .I2(n455[23]), 
            .I3(n24981), .O(n4_adj_4966));   // verilog/motorControl.v(63[16:31])
    defparam i1_2_lut_4_lut_adj_959.LUT_INIT = 16'hff8e;
    SB_LUT4 i47298_3_lut (.I0(n66145), .I1(n455[20]), .I2(n41_adj_4967), 
            .I3(GND_net), .O(n64360));   // verilog/motorControl.v(62[14:31])
    defparam i47298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n66663_bdd_4_lut (.I0(n66663), .I1(n535[15]), .I2(n455[15]), 
            .I3(n4744), .O(n66666));
    defparam n66663_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i48974_3_lut (.I0(n66035), .I1(n455[23]), .I2(n47_adj_4780), 
            .I3(GND_net), .O(n66036));   // verilog/motorControl.v(62[35:55])
    defparam i48974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48969_4_lut (.I0(n64360), .I1(n66029), .I2(n45_adj_4654), 
            .I3(n63737), .O(n66031));   // verilog/motorControl.v(62[14:31])
    defparam i48969_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 n9972_bdd_4_lut_49577 (.I0(n9972), .I1(n63019), .I2(setpoint[14]), 
            .I3(n4744), .O(n66657));
    defparam n9972_bdd_4_lut_49577.LUT_INIT = 16'he4aa;
    SB_LUT4 i46869_3_lut_4_lut (.I0(n233[3]), .I1(n285[3]), .I2(n285[2]), 
            .I3(n233[2]), .O(n63931));   // verilog/motorControl.v(58[23:46])
    defparam i46869_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 n66657_bdd_4_lut (.I0(n66657), .I1(n535[14]), .I2(n455[14]), 
            .I3(n4744), .O(n66660));
    defparam n66657_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 LessThan_19_i6_3_lut_3_lut (.I0(n233[3]), .I1(n285[3]), .I2(n285[2]), 
            .I3(GND_net), .O(n6_adj_4555));   // verilog/motorControl.v(58[23:46])
    defparam LessThan_19_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i22587_4_lut (.I0(n66031), .I1(n66036), .I2(deadband[23]), 
            .I3(n455[23]), .O(n38328));
    defparam i22587_4_lut.LUT_INIT = 16'hecfe;
    SB_LUT4 i3_4_lut_adj_960 (.I0(counter[6]), .I1(counter[4]), .I2(counter[0]), 
            .I3(counter[3]), .O(n58117));   // verilog/motorControl.v(27[8:42])
    defparam i3_4_lut_adj_960.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(n58117), .I1(counter[2]), .I2(counter[5]), .I3(counter[8]), 
            .O(n18_adj_4968));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(counter[7]), .I1(n18_adj_4968), .I2(counter[1]), 
            .I3(counter[10]), .O(n20_adj_4969));
    defparam i9_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i2_2_lut (.I0(counter[9]), .I1(counter[11]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_4970));   // verilog/motorControl.v(27[8:42])
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_961 (.I0(n7_adj_4970), .I1(counter[12]), .I2(counter[13]), 
            .I3(n20_adj_4969), .O(counter_31__N_3714));   // verilog/motorControl.v(27[8:42])
    defparam i4_4_lut_adj_961.LUT_INIT = 16'h0080;
    SB_LUT4 mult_23_i316_2_lut (.I0(\Kp[6] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_4451));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i365_2_lut (.I0(\Kp[7] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_4450));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32297_2_lut_3_lut (.I0(\Kp[0] ), .I1(n207[23]), .I2(\Kp[1] ), 
            .I3(GND_net), .O(n48010));   // verilog/motorControl.v(61[20:26])
    defparam i32297_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i32303_2_lut_3_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\Kp[2] ), 
            .I3(GND_net), .O(n49517));   // verilog/motorControl.v(61[20:26])
    defparam i32303_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 mult_23_i414_2_lut (.I0(\Kp[8] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n615));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_21_i12_3_lut (.I0(n233[11]), .I1(n285[11]), .I2(n284), 
            .I3(GND_net), .O(n310[11]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_21_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_22_i12_3_lut (.I0(n310[11]), .I1(IntegralLimit[11]), .I2(n258), 
            .I3(GND_net), .O(n335[11]));   // verilog/motorControl.v(58[20] 60[14])
    defparam mux_22_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_24_i71_2_lut (.I0(\Ki[1] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i24_2_lut (.I0(\Ki[0] ), .I1(n335[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4432));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i463_2_lut (.I0(\Kp[9] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i512_2_lut (.I0(\Kp[10] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i561_2_lut (.I0(\Kp[11] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46402_2_lut_4_lut (.I0(n455[21]), .I1(n535[21]), .I2(n455[9]), 
            .I3(n535[9]), .O(n63464));
    defparam i46402_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i120_2_lut (.I0(\Ki[2] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i610_2_lut (.I0(\Kp[12] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i659_2_lut (.I0(\Kp[13] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i69_2_lut (.I0(\Kp[1] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i22_2_lut (.I0(\Kp[0] ), .I1(n207[14]), .I2(GND_net), 
            .I3(GND_net), .O(n32));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46981_3_lut_4_lut (.I0(IntegralLimit[3]), .I1(n233[3]), .I2(n233[2]), 
            .I3(IntegralLimit[2]), .O(n64043));   // verilog/motorControl.v(56[14:36])
    defparam i46981_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_24_i169_2_lut (.I0(\Ki[3] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_17_i6_3_lut_3_lut (.I0(IntegralLimit[3]), .I1(n233[3]), 
            .I2(n233[2]), .I3(GND_net), .O(n6_adj_4498));   // verilog/motorControl.v(56[14:36])
    defparam LessThan_17_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_23_i118_2_lut (.I0(\Kp[2] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46426_2_lut_4_lut (.I0(n455[16]), .I1(n535[16]), .I2(n455[7]), 
            .I3(n535[7]), .O(n63488));
    defparam i46426_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i46656_2_lut_4_lut (.I0(deadband[21]), .I1(n455[21]), .I2(deadband[9]), 
            .I3(n455[9]), .O(n63718));
    defparam i46656_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i167_2_lut (.I0(\Kp[3] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n247));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i216_2_lut (.I0(\Kp[4] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n320));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46695_2_lut_4_lut (.I0(deadband[16]), .I1(n455[16]), .I2(deadband[7]), 
            .I3(n455[7]), .O(n63757));
    defparam i46695_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i32243_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[22]), .I2(n335[21]), 
            .I3(\Ki[1] ), .O(n20596[0]));   // verilog/motorControl.v(61[29:40])
    defparam i32243_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i32245_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[22]), .I2(n335[21]), 
            .I3(\Ki[1] ), .O(n47955));   // verilog/motorControl.v(61[29:40])
    defparam i32245_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i46984_2_lut_4_lut (.I0(setpoint[21]), .I1(n535[21]), .I2(setpoint[9]), 
            .I3(n535[9]), .O(n64046));
    defparam i46984_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i32272_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[21]), .I2(n335[20]), 
            .I3(\Ki[1] ), .O(n20575[0]));   // verilog/motorControl.v(61[29:40])
    defparam i32272_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i32274_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[21]), .I2(n335[20]), 
            .I3(\Ki[1] ), .O(n47985));   // verilog/motorControl.v(61[29:40])
    defparam i32274_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_24_i218_2_lut (.I0(\Ki[4] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_962 (.I0(\Ki[3] ), .I1(n335[19]), .I2(n4_adj_4972), 
            .I3(n20575[1]), .O(n20538[2]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_962.LUT_INIT = 16'h8778;
    SB_LUT4 mult_23_i265_2_lut (.I0(\Kp[5] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32340_3_lut_4_lut (.I0(\Ki[3] ), .I1(n335[19]), .I2(n4_adj_4972), 
            .I3(n20575[1]), .O(n6_adj_4955));   // verilog/motorControl.v(61[29:40])
    defparam i32340_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i32332_3_lut_4_lut (.I0(\Ki[2] ), .I1(n335[19]), .I2(n48038), 
            .I3(n20575[0]), .O(n4_adj_4972));   // verilog/motorControl.v(61[29:40])
    defparam i32332_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i46756_2_lut_4_lut (.I0(n233[21]), .I1(n285[21]), .I2(n233[9]), 
            .I3(n285[9]), .O(n63818));
    defparam i46756_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_3_lut_4_lut_adj_963 (.I0(\Ki[2] ), .I1(n335[19]), .I2(n48038), 
            .I3(n20575[0]), .O(n20538[1]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_963.LUT_INIT = 16'h8778;
    SB_LUT4 i32319_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[20]), .I2(n335[19]), 
            .I3(\Ki[1] ), .O(n20538[0]));   // verilog/motorControl.v(61[29:40])
    defparam i32319_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i32321_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[20]), .I2(n335[19]), 
            .I3(\Ki[1] ), .O(n48038));   // verilog/motorControl.v(61[29:40])
    defparam i32321_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i47014_2_lut_4_lut (.I0(setpoint[16]), .I1(n535[16]), .I2(setpoint[7]), 
            .I3(n535[7]), .O(n64076));
    defparam i47014_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i46810_2_lut_4_lut (.I0(n233[16]), .I1(n285[16]), .I2(n233[7]), 
            .I3(n285[7]), .O(n63872));
    defparam i46810_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_23_i314_2_lut (.I0(\Kp[6] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n466));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32415_3_lut_4_lut (.I0(\Ki[3] ), .I1(n335[18]), .I2(n4_adj_4973), 
            .I3(n20538[1]), .O(n6_adj_4949));   // verilog/motorControl.v(61[29:40])
    defparam i32415_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_23_i363_2_lut (.I0(\Kp[7] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n539));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i412_2_lut (.I0(\Kp[8] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n612));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i267_2_lut (.I0(\Ki[5] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i461_2_lut (.I0(\Kp[9] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_23_i510_2_lut (.I0(\Kp[10] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_964 (.I0(\Ki[3] ), .I1(n335[18]), .I2(n4_adj_4973), 
            .I3(n20538[1]), .O(n20481[2]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_964.LUT_INIT = 16'h8778;
    SB_LUT4 i1_3_lut_4_lut_adj_965 (.I0(\Ki[2] ), .I1(n335[18]), .I2(n48119), 
            .I3(n20538[0]), .O(n20481[1]));   // verilog/motorControl.v(61[29:40])
    defparam i1_3_lut_4_lut_adj_965.LUT_INIT = 16'h8778;
    SB_LUT4 i32407_3_lut_4_lut (.I0(\Ki[2] ), .I1(n335[18]), .I2(n48119), 
            .I3(n20538[0]), .O(n4_adj_4973));   // verilog/motorControl.v(61[29:40])
    defparam i32407_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i32394_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[19]), .I2(n335[18]), 
            .I3(\Ki[1] ), .O(n20481[0]));   // verilog/motorControl.v(61[29:40])
    defparam i32394_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i32396_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(n335[19]), .I2(n335[18]), 
            .I3(\Ki[1] ), .O(n48119));   // verilog/motorControl.v(61[29:40])
    defparam i32396_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_23_i559_2_lut (.I0(\Kp[11] ), .I1(n207[13]), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(61[20:26])
    defparam mult_23_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_24_i316_2_lut (.I0(\Ki[6] ), .I1(n335[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_4430));   // verilog/motorControl.v(61[29:40])
    defparam mult_24_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i46873_2_lut_4_lut (.I0(IntegralLimit[21]), .I1(n233[21]), .I2(IntegralLimit[9]), 
            .I3(n233[9]), .O(n63935));
    defparam i46873_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i46928_2_lut_4_lut (.I0(IntegralLimit[16]), .I1(n233[16]), .I2(IntegralLimit[7]), 
            .I3(n233[7]), .O(n63990));
    defparam i46928_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i4_4_lut_adj_966 (.I0(control_mode[7]), .I1(control_mode[0]), 
            .I2(control_mode[1]), .I3(control_mode[4]), .O(n10_adj_4974));
    defparam i4_4_lut_adj_966.LUT_INIT = 16'h0040;
    SB_LUT4 LessThan_30_i45_2_lut (.I0(PWMLimit[22]), .I1(n455[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut (.I0(control_mode[6]), .I1(n10_adj_4974), .I2(control_mode[5]), 
            .I3(GND_net), .O(n55181));
    defparam i5_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 LessThan_9_i31_2_lut (.I0(PWMLimit[15]), .I1(setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4975));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i37_2_lut (.I0(PWMLimit[18]), .I1(n455[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4487));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i29_2_lut (.I0(PWMLimit[14]), .I1(setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4976));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i27_2_lut (.I0(PWMLimit[13]), .I1(setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4977));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i19_2_lut (.I0(PWMLimit[9]), .I1(setpoint[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4978));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i23_2_lut (.I0(PWMLimit[11]), .I1(setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4979));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i39_2_lut (.I0(PWMLimit[19]), .I1(n455[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4503));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i15_2_lut (.I0(PWMLimit[7]), .I1(setpoint[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4980));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i41_2_lut (.I0(PWMLimit[20]), .I1(n455[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4507));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i17_2_lut (.I0(PWMLimit[8]), .I1(setpoint[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4981));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i7_2_lut (.I0(PWMLimit[3]), .I1(setpoint[3]), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_4982));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i9_2_lut (.I0(PWMLimit[4]), .I1(setpoint[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4983));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i11_2_lut (.I0(PWMLimit[5]), .I1(setpoint[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4984));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i13_2_lut (.I0(PWMLimit[6]), .I1(setpoint[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4985));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i43_2_lut (.I0(PWMLimit[21]), .I1(n455[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4431));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i5_2_lut (.I0(PWMLimit[2]), .I1(setpoint[2]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4986));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i46206_4_lut (.I0(n11_adj_4984), .I1(n9_adj_4983), .I2(n7_adj_4982), 
            .I3(n5_adj_4986), .O(n63268));
    defparam i46206_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i46191_4_lut (.I0(n17_adj_4981), .I1(n15_adj_4980), .I2(n13_adj_4985), 
            .I3(n63268), .O(n63253));
    defparam i46191_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48379_4_lut (.I0(n23_adj_4979), .I1(n21), .I2(n19_adj_4978), 
            .I3(n63253), .O(n65441));
    defparam i48379_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_9_i4_4_lut (.I0(PWMLimit[0]), .I1(setpoint[1]), .I2(PWMLimit[1]), 
            .I3(setpoint[0]), .O(n4_adj_4988));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i48428_3_lut (.I0(n4_adj_4988), .I1(setpoint[13]), .I2(n27_adj_4977), 
            .I3(GND_net), .O(n65490));   // verilog/motorControl.v(45[16:33])
    defparam i48428_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48429_3_lut (.I0(n65490), .I1(setpoint[14]), .I2(n29_adj_4976), 
            .I3(GND_net), .O(n65491));   // verilog/motorControl.v(45[16:33])
    defparam i48429_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47140_4_lut (.I0(n29_adj_4976), .I1(n27_adj_4977), .I2(n15_adj_4980), 
            .I3(n63259), .O(n64202));
    defparam i47140_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i48041_3_lut (.I0(n10_adj_4959), .I1(setpoint[7]), .I2(n15_adj_4980), 
            .I3(GND_net), .O(n65103));   // verilog/motorControl.v(45[16:33])
    defparam i48041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i35_2_lut (.I0(PWMLimit[17]), .I1(n455[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4486));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48402_3_lut (.I0(n65491), .I1(setpoint[15]), .I2(n31_adj_4975), 
            .I3(GND_net), .O(n65464));   // verilog/motorControl.v(45[16:33])
    defparam i48402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i29_2_lut (.I0(PWMLimit[14]), .I1(n455[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4467));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_9_i16_3_lut (.I0(n8_adj_4958), .I1(setpoint[9]), .I2(n19_adj_4978), 
            .I3(GND_net), .O(n16_adj_4989));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i49037_4_lut (.I0(n16_adj_4989), .I1(n6_adj_4957), .I2(n19_adj_4978), 
            .I3(n63239), .O(n66099));   // verilog/motorControl.v(45[16:33])
    defparam i49037_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i49038_3_lut (.I0(n66099), .I1(setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n66100));   // verilog/motorControl.v(45[16:33])
    defparam i49038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48946_3_lut (.I0(n66100), .I1(setpoint[11]), .I2(n23_adj_4979), 
            .I3(GND_net), .O(n66008));   // verilog/motorControl.v(45[16:33])
    defparam i48946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i31_2_lut (.I0(PWMLimit[15]), .I1(n455[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4473));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 n9972_bdd_4_lut_49572 (.I0(n9972), .I1(n62945), .I2(setpoint[13]), 
            .I3(n4744), .O(n66567));
    defparam n9972_bdd_4_lut_49572.LUT_INIT = 16'he4aa;
    SB_LUT4 i47142_4_lut (.I0(n29_adj_4976), .I1(n27_adj_4977), .I2(n25), 
            .I3(n65441), .O(n64204));
    defparam i47142_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i48426_4_lut (.I0(n65464), .I1(n65103), .I2(n31_adj_4975), 
            .I3(n64202), .O(n65488));   // verilog/motorControl.v(45[16:33])
    defparam i48426_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i48744_3_lut (.I0(n66008), .I1(setpoint[12]), .I2(n25), .I3(GND_net), 
            .O(n65806));   // verilog/motorControl.v(45[16:33])
    defparam i48744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i48979_4_lut (.I0(n65806), .I1(n65488), .I2(n31_adj_4975), 
            .I3(n64204), .O(n66041));   // verilog/motorControl.v(45[16:33])
    defparam i48979_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i48980_3_lut (.I0(n66041), .I1(setpoint[16]), .I2(PWMLimit[16]), 
            .I3(GND_net), .O(n66042));   // verilog/motorControl.v(45[16:33])
    defparam i48980_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_9_i36_3_lut (.I0(n66042), .I1(setpoint[17]), .I2(PWMLimit[17]), 
            .I3(GND_net), .O(n36));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i36_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_9_i40_3_lut (.I0(n33833), .I1(setpoint[19]), .I2(PWMLimit[19]), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(45[16:33])
    defparam LessThan_9_i40_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_30_i33_2_lut (.I0(PWMLimit[16]), .I1(n455[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4472));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i48424_3_lut (.I0(n33791), .I1(setpoint[21]), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n65486));   // verilog/motorControl.v(45[16:33])
    defparam i48424_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i46554_4_lut (.I0(n21_c), .I1(n19_adj_4947), .I2(n17), .I3(n9_adj_4943), 
            .O(n63616));
    defparam i46554_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i48425_3_lut (.I0(n65486), .I1(setpoint[22]), .I2(PWMLimit[22]), 
            .I3(GND_net), .O(n65487));   // verilog/motorControl.v(45[16:33])
    defparam i48425_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i48407_3_lut (.I0(n65487), .I1(PWMLimit[23]), .I2(setpoint[23]), 
            .I3(GND_net), .O(n105));   // verilog/motorControl.v(45[16:33])
    defparam i48407_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 n66567_bdd_4_lut (.I0(n66567), .I1(n535[13]), .I2(n455[13]), 
            .I3(n4744), .O(n66570));
    defparam n66567_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i46534_4_lut (.I0(n27), .I1(n15_adj_4946), .I2(n13_adj_4945), 
            .I3(n11_adj_4944), .O(n63596));
    defparam i46534_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_30_i12_3_lut (.I0(n455[7]), .I1(n455[16]), .I2(n33_adj_4472), 
            .I3(GND_net), .O(n12_adj_4991));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i10_3_lut (.I0(n455[5]), .I1(n455[6]), .I2(n13_adj_4945), 
            .I3(GND_net), .O(n10));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_30_i30_3_lut (.I0(n12_adj_4991), .I1(n455[17]), .I2(n35_adj_4486), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i47554_4_lut (.I0(n13_adj_4945), .I1(n11_adj_4944), .I2(n9_adj_4943), 
            .I3(n63644), .O(n64616));
    defparam i47554_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i47546_4_lut (.I0(n19_adj_4947), .I1(n17), .I2(n15_adj_4946), 
            .I3(n64616), .O(n64608));
    defparam i47546_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i48809_4_lut (.I0(n25_c), .I1(n23), .I2(n21_c), .I3(n64608), 
            .O(n65871));
    defparam i48809_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i48119_4_lut (.I0(n31_adj_4473), .I1(n29_adj_4467), .I2(n27), 
            .I3(n65871), .O(n65181));
    defparam i48119_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i48998_4_lut (.I0(n37_adj_4487), .I1(n35_adj_4486), .I2(n33_adj_4472), 
            .I3(n65181), .O(n66060));
    defparam i48998_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_26_i41_2_lut (.I0(deadband[20]), .I1(n455[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4967));   // verilog/motorControl.v(62[14:31])
    defparam LessThan_26_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_30_i16_3_lut (.I0(n455[9]), .I1(n455[21]), .I2(n43_adj_4431), 
            .I3(GND_net), .O(n16));   // verilog/motorControl.v(63[16:31])
    defparam LessThan_30_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i46487_2_lut_4_lut (.I0(PWMLimit[21]), .I1(n455[21]), .I2(PWMLimit[9]), 
            .I3(n455[9]), .O(n63549));
    defparam i46487_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    
endmodule
