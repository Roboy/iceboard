// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Jan 29 2020 19:19:01

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    TX,
    SDA,
    SCL,
    RX,
    NEOPXL,
    LED,
    INLC,
    INLB,
    INLA,
    INHC,
    INHB,
    INHA,
    HALL3,
    HALL2,
    HALL1,
    FAULT_N,
    ENCODER1_B,
    ENCODER1_A,
    ENCODER0_B,
    ENCODER0_A,
    DE,
    CS_MISO,
    CS_CLK,
    CS,
    CLK);

    output USBPU;
    output TX;
    inout SDA;
    inout SCL;
    input RX;
    output NEOPXL;
    output LED;
    output INLC;
    output INLB;
    output INLA;
    output INHC;
    output INHB;
    output INHA;
    input HALL3;
    input HALL2;
    input HALL1;
    input FAULT_N;
    input ENCODER1_B;
    input ENCODER1_A;
    input ENCODER0_B;
    input ENCODER0_A;
    output DE;
    input CS_MISO;
    output CS_CLK;
    output CS;
    input CLK;

    wire N__6589;
    wire N__6588;
    wire N__6587;
    wire N__6580;
    wire N__6579;
    wire N__6578;
    wire N__6571;
    wire N__6570;
    wire N__6569;
    wire N__6562;
    wire N__6561;
    wire N__6560;
    wire N__6553;
    wire N__6552;
    wire N__6551;
    wire N__6544;
    wire N__6543;
    wire N__6542;
    wire N__6535;
    wire N__6534;
    wire N__6533;
    wire N__6526;
    wire N__6525;
    wire N__6524;
    wire N__6517;
    wire N__6516;
    wire N__6515;
    wire N__6508;
    wire N__6507;
    wire N__6506;
    wire N__6499;
    wire N__6498;
    wire N__6497;
    wire N__6490;
    wire N__6489;
    wire N__6488;
    wire N__6481;
    wire N__6480;
    wire N__6479;
    wire N__6472;
    wire N__6471;
    wire N__6470;
    wire N__6463;
    wire N__6462;
    wire N__6461;
    wire N__6454;
    wire N__6453;
    wire N__6452;
    wire N__6435;
    wire N__6434;
    wire N__6433;
    wire N__6428;
    wire N__6425;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6408;
    wire N__6405;
    wire N__6402;
    wire N__6399;
    wire N__6396;
    wire N__6393;
    wire N__6390;
    wire N__6387;
    wire N__6384;
    wire N__6383;
    wire N__6382;
    wire N__6381;
    wire N__6380;
    wire N__6379;
    wire N__6374;
    wire N__6371;
    wire N__6366;
    wire N__6363;
    wire N__6354;
    wire N__6353;
    wire N__6352;
    wire N__6349;
    wire N__6348;
    wire N__6347;
    wire N__6346;
    wire N__6341;
    wire N__6338;
    wire N__6335;
    wire N__6332;
    wire N__6329;
    wire N__6318;
    wire N__6315;
    wire N__6312;
    wire N__6311;
    wire N__6310;
    wire N__6307;
    wire N__6306;
    wire N__6301;
    wire N__6296;
    wire N__6293;
    wire N__6290;
    wire N__6285;
    wire N__6282;
    wire N__6279;
    wire N__6276;
    wire N__6273;
    wire N__6270;
    wire N__6269;
    wire N__6268;
    wire N__6267;
    wire N__6266;
    wire N__6265;
    wire N__6262;
    wire N__6259;
    wire N__6258;
    wire N__6257;
    wire N__6256;
    wire N__6247;
    wire N__6246;
    wire N__6245;
    wire N__6242;
    wire N__6239;
    wire N__6232;
    wire N__6229;
    wire N__6224;
    wire N__6213;
    wire N__6210;
    wire N__6207;
    wire N__6204;
    wire N__6201;
    wire N__6198;
    wire N__6195;
    wire N__6194;
    wire N__6191;
    wire N__6188;
    wire N__6183;
    wire N__6182;
    wire N__6181;
    wire N__6180;
    wire N__6177;
    wire N__6174;
    wire N__6171;
    wire N__6170;
    wire N__6169;
    wire N__6166;
    wire N__6165;
    wire N__6162;
    wire N__6157;
    wire N__6154;
    wire N__6153;
    wire N__6150;
    wire N__6147;
    wire N__6144;
    wire N__6137;
    wire N__6134;
    wire N__6131;
    wire N__6130;
    wire N__6129;
    wire N__6126;
    wire N__6123;
    wire N__6118;
    wire N__6117;
    wire N__6114;
    wire N__6111;
    wire N__6110;
    wire N__6107;
    wire N__6106;
    wire N__6103;
    wire N__6100;
    wire N__6097;
    wire N__6094;
    wire N__6089;
    wire N__6086;
    wire N__6083;
    wire N__6080;
    wire N__6063;
    wire N__6060;
    wire N__6057;
    wire N__6054;
    wire N__6051;
    wire N__6050;
    wire N__6047;
    wire N__6044;
    wire N__6039;
    wire N__6036;
    wire N__6033;
    wire N__6032;
    wire N__6029;
    wire N__6026;
    wire N__6021;
    wire N__6018;
    wire N__6015;
    wire N__6014;
    wire N__6011;
    wire N__6008;
    wire N__6003;
    wire N__6000;
    wire N__5997;
    wire N__5994;
    wire N__5991;
    wire N__5988;
    wire N__5987;
    wire N__5986;
    wire N__5985;
    wire N__5984;
    wire N__5981;
    wire N__5980;
    wire N__5977;
    wire N__5976;
    wire N__5973;
    wire N__5958;
    wire N__5955;
    wire N__5952;
    wire N__5951;
    wire N__5948;
    wire N__5947;
    wire N__5946;
    wire N__5945;
    wire N__5944;
    wire N__5939;
    wire N__5936;
    wire N__5933;
    wire N__5930;
    wire N__5929;
    wire N__5926;
    wire N__5923;
    wire N__5920;
    wire N__5917;
    wire N__5910;
    wire N__5909;
    wire N__5908;
    wire N__5905;
    wire N__5902;
    wire N__5897;
    wire N__5894;
    wire N__5891;
    wire N__5880;
    wire N__5877;
    wire N__5876;
    wire N__5875;
    wire N__5874;
    wire N__5873;
    wire N__5872;
    wire N__5871;
    wire N__5870;
    wire N__5867;
    wire N__5862;
    wire N__5861;
    wire N__5860;
    wire N__5859;
    wire N__5858;
    wire N__5857;
    wire N__5854;
    wire N__5845;
    wire N__5844;
    wire N__5843;
    wire N__5842;
    wire N__5841;
    wire N__5840;
    wire N__5839;
    wire N__5838;
    wire N__5837;
    wire N__5834;
    wire N__5831;
    wire N__5828;
    wire N__5825;
    wire N__5818;
    wire N__5813;
    wire N__5804;
    wire N__5795;
    wire N__5778;
    wire N__5777;
    wire N__5776;
    wire N__5773;
    wire N__5772;
    wire N__5771;
    wire N__5770;
    wire N__5769;
    wire N__5768;
    wire N__5767;
    wire N__5766;
    wire N__5765;
    wire N__5762;
    wire N__5761;
    wire N__5760;
    wire N__5759;
    wire N__5758;
    wire N__5751;
    wire N__5746;
    wire N__5745;
    wire N__5744;
    wire N__5743;
    wire N__5742;
    wire N__5741;
    wire N__5738;
    wire N__5735;
    wire N__5728;
    wire N__5727;
    wire N__5726;
    wire N__5725;
    wire N__5724;
    wire N__5721;
    wire N__5718;
    wire N__5715;
    wire N__5710;
    wire N__5705;
    wire N__5694;
    wire N__5687;
    wire N__5678;
    wire N__5661;
    wire N__5660;
    wire N__5657;
    wire N__5654;
    wire N__5653;
    wire N__5652;
    wire N__5651;
    wire N__5650;
    wire N__5649;
    wire N__5648;
    wire N__5645;
    wire N__5640;
    wire N__5639;
    wire N__5638;
    wire N__5637;
    wire N__5632;
    wire N__5631;
    wire N__5630;
    wire N__5629;
    wire N__5626;
    wire N__5625;
    wire N__5624;
    wire N__5623;
    wire N__5620;
    wire N__5619;
    wire N__5618;
    wire N__5617;
    wire N__5616;
    wire N__5615;
    wire N__5612;
    wire N__5607;
    wire N__5600;
    wire N__5597;
    wire N__5588;
    wire N__5581;
    wire N__5578;
    wire N__5565;
    wire N__5550;
    wire N__5549;
    wire N__5548;
    wire N__5545;
    wire N__5540;
    wire N__5539;
    wire N__5538;
    wire N__5537;
    wire N__5536;
    wire N__5535;
    wire N__5534;
    wire N__5533;
    wire N__5532;
    wire N__5529;
    wire N__5526;
    wire N__5525;
    wire N__5524;
    wire N__5523;
    wire N__5522;
    wire N__5521;
    wire N__5518;
    wire N__5517;
    wire N__5516;
    wire N__5515;
    wire N__5510;
    wire N__5505;
    wire N__5498;
    wire N__5493;
    wire N__5490;
    wire N__5481;
    wire N__5472;
    wire N__5457;
    wire N__5456;
    wire N__5453;
    wire N__5450;
    wire N__5447;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5430;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5418;
    wire N__5415;
    wire N__5414;
    wire N__5413;
    wire N__5406;
    wire N__5403;
    wire N__5400;
    wire N__5397;
    wire N__5396;
    wire N__5393;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5373;
    wire N__5372;
    wire N__5369;
    wire N__5366;
    wire N__5363;
    wire N__5358;
    wire N__5355;
    wire N__5354;
    wire N__5351;
    wire N__5348;
    wire N__5343;
    wire N__5342;
    wire N__5337;
    wire N__5336;
    wire N__5335;
    wire N__5334;
    wire N__5331;
    wire N__5328;
    wire N__5325;
    wire N__5322;
    wire N__5313;
    wire N__5310;
    wire N__5307;
    wire N__5304;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5292;
    wire N__5289;
    wire N__5288;
    wire N__5285;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5271;
    wire N__5268;
    wire N__5265;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5253;
    wire N__5250;
    wire N__5247;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5199;
    wire N__5196;
    wire N__5195;
    wire N__5192;
    wire N__5189;
    wire N__5184;
    wire N__5181;
    wire N__5180;
    wire N__5177;
    wire N__5174;
    wire N__5169;
    wire N__5166;
    wire N__5165;
    wire N__5162;
    wire N__5159;
    wire N__5154;
    wire N__5151;
    wire N__5148;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5136;
    wire N__5135;
    wire N__5134;
    wire N__5133;
    wire N__5132;
    wire N__5131;
    wire N__5130;
    wire N__5129;
    wire N__5128;
    wire N__5127;
    wire N__5126;
    wire N__5125;
    wire N__5124;
    wire N__5123;
    wire N__5122;
    wire N__5121;
    wire N__5120;
    wire N__5119;
    wire N__5118;
    wire N__5117;
    wire N__5076;
    wire N__5073;
    wire N__5070;
    wire N__5067;
    wire N__5066;
    wire N__5065;
    wire N__5062;
    wire N__5059;
    wire N__5056;
    wire N__5049;
    wire N__5046;
    wire N__5043;
    wire N__5040;
    wire N__5039;
    wire N__5038;
    wire N__5035;
    wire N__5030;
    wire N__5025;
    wire N__5022;
    wire N__5021;
    wire N__5018;
    wire N__5015;
    wire N__5010;
    wire N__5007;
    wire N__5004;
    wire N__5001;
    wire N__4998;
    wire N__4995;
    wire N__4992;
    wire N__4989;
    wire N__4986;
    wire N__4985;
    wire N__4982;
    wire N__4979;
    wire N__4976;
    wire N__4971;
    wire N__4968;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4958;
    wire N__4957;
    wire N__4954;
    wire N__4951;
    wire N__4948;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4928;
    wire N__4925;
    wire N__4924;
    wire N__4923;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4899;
    wire N__4896;
    wire N__4893;
    wire N__4890;
    wire N__4887;
    wire N__4884;
    wire N__4883;
    wire N__4880;
    wire N__4877;
    wire N__4872;
    wire N__4869;
    wire N__4866;
    wire N__4863;
    wire N__4860;
    wire N__4857;
    wire N__4856;
    wire N__4853;
    wire N__4850;
    wire N__4849;
    wire N__4846;
    wire N__4843;
    wire N__4840;
    wire N__4837;
    wire N__4834;
    wire N__4831;
    wire N__4824;
    wire N__4821;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4809;
    wire N__4806;
    wire N__4803;
    wire N__4800;
    wire N__4799;
    wire N__4798;
    wire N__4795;
    wire N__4792;
    wire N__4789;
    wire N__4782;
    wire N__4779;
    wire N__4776;
    wire N__4773;
    wire N__4770;
    wire N__4767;
    wire N__4764;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4752;
    wire N__4749;
    wire N__4746;
    wire N__4743;
    wire N__4740;
    wire N__4737;
    wire N__4734;
    wire N__4731;
    wire N__4730;
    wire N__4725;
    wire N__4722;
    wire N__4719;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4707;
    wire N__4704;
    wire N__4701;
    wire N__4700;
    wire N__4699;
    wire N__4696;
    wire N__4693;
    wire N__4690;
    wire N__4687;
    wire N__4680;
    wire N__4677;
    wire N__4674;
    wire N__4671;
    wire N__4668;
    wire N__4665;
    wire N__4664;
    wire N__4663;
    wire N__4660;
    wire N__4655;
    wire N__4650;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4642;
    wire N__4639;
    wire N__4636;
    wire N__4633;
    wire N__4626;
    wire N__4623;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4610;
    wire N__4609;
    wire N__4604;
    wire N__4601;
    wire N__4596;
    wire N__4593;
    wire N__4590;
    wire N__4587;
    wire N__4584;
    wire N__4583;
    wire N__4582;
    wire N__4579;
    wire N__4574;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4562;
    wire N__4561;
    wire N__4558;
    wire N__4553;
    wire N__4548;
    wire N__4547;
    wire N__4546;
    wire N__4545;
    wire N__4544;
    wire N__4543;
    wire N__4542;
    wire N__4541;
    wire N__4540;
    wire N__4539;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4531;
    wire N__4530;
    wire N__4529;
    wire N__4528;
    wire N__4525;
    wire N__4522;
    wire N__4519;
    wire N__4518;
    wire N__4517;
    wire N__4516;
    wire N__4507;
    wire N__4504;
    wire N__4501;
    wire N__4496;
    wire N__4491;
    wire N__4486;
    wire N__4475;
    wire N__4474;
    wire N__4473;
    wire N__4472;
    wire N__4471;
    wire N__4470;
    wire N__4469;
    wire N__4468;
    wire N__4467;
    wire N__4464;
    wire N__4461;
    wire N__4458;
    wire N__4451;
    wire N__4446;
    wire N__4439;
    wire N__4428;
    wire N__4413;
    wire N__4412;
    wire N__4411;
    wire N__4410;
    wire N__4409;
    wire N__4408;
    wire N__4405;
    wire N__4404;
    wire N__4401;
    wire N__4398;
    wire N__4395;
    wire N__4392;
    wire N__4387;
    wire N__4384;
    wire N__4377;
    wire N__4374;
    wire N__4373;
    wire N__4372;
    wire N__4371;
    wire N__4370;
    wire N__4367;
    wire N__4362;
    wire N__4359;
    wire N__4358;
    wire N__4357;
    wire N__4356;
    wire N__4353;
    wire N__4350;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4342;
    wire N__4339;
    wire N__4336;
    wire N__4333;
    wire N__4322;
    wire N__4319;
    wire N__4312;
    wire N__4299;
    wire N__4296;
    wire N__4293;
    wire N__4292;
    wire N__4289;
    wire N__4288;
    wire N__4285;
    wire N__4282;
    wire N__4279;
    wire N__4272;
    wire N__4271;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4257;
    wire N__4254;
    wire N__4251;
    wire N__4248;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4238;
    wire N__4233;
    wire N__4230;
    wire N__4227;
    wire N__4224;
    wire N__4221;
    wire N__4220;
    wire N__4219;
    wire N__4218;
    wire N__4215;
    wire N__4210;
    wire N__4207;
    wire N__4204;
    wire N__4201;
    wire N__4198;
    wire N__4193;
    wire N__4188;
    wire N__4187;
    wire N__4184;
    wire N__4181;
    wire N__4176;
    wire N__4175;
    wire N__4172;
    wire N__4169;
    wire N__4164;
    wire N__4163;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4149;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4137;
    wire N__4136;
    wire N__4135;
    wire N__4130;
    wire N__4127;
    wire N__4124;
    wire N__4119;
    wire N__4116;
    wire N__4113;
    wire N__4112;
    wire N__4111;
    wire N__4108;
    wire N__4105;
    wire N__4102;
    wire N__4101;
    wire N__4096;
    wire N__4093;
    wire N__4090;
    wire N__4087;
    wire N__4084;
    wire N__4081;
    wire N__4074;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4062;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4050;
    wire N__4049;
    wire N__4044;
    wire N__4041;
    wire N__4038;
    wire N__4037;
    wire N__4034;
    wire N__4031;
    wire N__4026;
    wire N__4025;
    wire N__4022;
    wire N__4019;
    wire N__4014;
    wire N__4013;
    wire N__4010;
    wire N__4007;
    wire N__4004;
    wire N__3999;
    wire N__3998;
    wire N__3995;
    wire N__3992;
    wire N__3987;
    wire N__3984;
    wire N__3983;
    wire N__3980;
    wire N__3977;
    wire N__3974;
    wire N__3971;
    wire N__3966;
    wire N__3963;
    wire N__3960;
    wire N__3957;
    wire N__3954;
    wire N__3953;
    wire N__3952;
    wire N__3951;
    wire N__3950;
    wire N__3949;
    wire N__3948;
    wire N__3947;
    wire N__3944;
    wire N__3941;
    wire N__3936;
    wire N__3927;
    wire N__3918;
    wire N__3915;
    wire N__3912;
    wire N__3909;
    wire N__3908;
    wire N__3905;
    wire N__3902;
    wire N__3897;
    wire N__3896;
    wire N__3893;
    wire N__3890;
    wire N__3885;
    wire N__3884;
    wire N__3881;
    wire N__3878;
    wire N__3875;
    wire N__3870;
    wire N__3869;
    wire N__3866;
    wire N__3863;
    wire N__3858;
    wire N__3857;
    wire N__3854;
    wire N__3851;
    wire N__3846;
    wire N__3845;
    wire N__3842;
    wire N__3839;
    wire N__3834;
    wire N__3833;
    wire N__3830;
    wire N__3827;
    wire N__3824;
    wire N__3819;
    wire N__3818;
    wire N__3815;
    wire N__3812;
    wire N__3807;
    wire N__3804;
    wire N__3803;
    wire N__3800;
    wire N__3797;
    wire N__3792;
    wire N__3791;
    wire N__3788;
    wire N__3785;
    wire N__3780;
    wire N__3777;
    wire N__3776;
    wire N__3773;
    wire N__3770;
    wire N__3765;
    wire N__3764;
    wire N__3761;
    wire N__3758;
    wire N__3753;
    wire N__3752;
    wire N__3749;
    wire N__3746;
    wire N__3741;
    wire N__3740;
    wire N__3737;
    wire N__3734;
    wire N__3731;
    wire N__3726;
    wire N__3725;
    wire N__3722;
    wire N__3719;
    wire N__3714;
    wire N__3713;
    wire N__3710;
    wire N__3707;
    wire N__3702;
    wire N__3701;
    wire N__3698;
    wire N__3695;
    wire N__3690;
    wire N__3689;
    wire N__3686;
    wire N__3683;
    wire N__3678;
    wire N__3675;
    wire N__3672;
    wire N__3671;
    wire N__3668;
    wire N__3665;
    wire N__3660;
    wire N__3659;
    wire N__3656;
    wire N__3653;
    wire N__3648;
    wire N__3645;
    wire N__3642;
    wire N__3639;
    wire N__3636;
    wire N__3633;
    wire N__3630;
    wire N__3627;
    wire N__3626;
    wire N__3625;
    wire N__3622;
    wire N__3617;
    wire N__3612;
    wire N__3609;
    wire N__3606;
    wire N__3605;
    wire N__3604;
    wire N__3603;
    wire N__3600;
    wire N__3597;
    wire N__3592;
    wire N__3585;
    wire N__3582;
    wire N__3579;
    wire N__3576;
    wire N__3573;
    wire N__3570;
    wire N__3567;
    wire N__3564;
    wire N__3561;
    wire N__3558;
    wire N__3555;
    wire N__3554;
    wire N__3553;
    wire N__3552;
    wire N__3551;
    wire N__3550;
    wire N__3549;
    wire N__3548;
    wire N__3547;
    wire N__3544;
    wire N__3543;
    wire N__3540;
    wire N__3539;
    wire N__3536;
    wire N__3535;
    wire N__3532;
    wire N__3529;
    wire N__3528;
    wire N__3525;
    wire N__3524;
    wire N__3521;
    wire N__3520;
    wire N__3517;
    wire N__3516;
    wire N__3499;
    wire N__3482;
    wire N__3477;
    wire N__3474;
    wire N__3471;
    wire N__3468;
    wire N__3465;
    wire N__3462;
    wire N__3459;
    wire N__3456;
    wire N__3453;
    wire N__3450;
    wire N__3449;
    wire N__3448;
    wire N__3445;
    wire N__3440;
    wire N__3435;
    wire N__3432;
    wire N__3429;
    wire N__3426;
    wire N__3423;
    wire N__3420;
    wire N__3419;
    wire N__3418;
    wire N__3415;
    wire N__3410;
    wire N__3405;
    wire N__3402;
    wire N__3399;
    wire N__3396;
    wire N__3393;
    wire N__3392;
    wire N__3391;
    wire N__3388;
    wire N__3383;
    wire N__3378;
    wire N__3375;
    wire N__3372;
    wire N__3371;
    wire N__3370;
    wire N__3367;
    wire N__3364;
    wire N__3359;
    wire N__3354;
    wire N__3351;
    wire N__3348;
    wire N__3347;
    wire N__3344;
    wire N__3343;
    wire N__3340;
    wire N__3337;
    wire N__3332;
    wire N__3327;
    wire N__3324;
    wire N__3321;
    wire N__3318;
    wire N__3315;
    wire N__3312;
    wire N__3311;
    wire N__3310;
    wire N__3307;
    wire N__3302;
    wire N__3297;
    wire N__3294;
    wire N__3291;
    wire N__3288;
    wire N__3285;
    wire N__3282;
    wire N__3279;
    wire N__3278;
    wire N__3277;
    wire N__3274;
    wire N__3269;
    wire N__3264;
    wire N__3261;
    wire N__3258;
    wire N__3255;
    wire N__3252;
    wire N__3249;
    wire N__3246;
    wire N__3243;
    wire N__3240;
    wire N__3237;
    wire N__3234;
    wire N__3231;
    wire N__3228;
    wire N__3227;
    wire N__3226;
    wire N__3223;
    wire N__3218;
    wire N__3213;
    wire N__3210;
    wire N__3207;
    wire N__3204;
    wire N__3201;
    wire N__3198;
    wire N__3195;
    wire N__3192;
    wire N__3189;
    wire N__3186;
    wire N__3183;
    wire N__3180;
    wire N__3177;
    wire N__3174;
    wire N__3171;
    wire N__3168;
    wire N__3165;
    wire N__3162;
    wire N__3159;
    wire N__3156;
    wire N__3153;
    wire N__3150;
    wire N__3147;
    wire N__3144;
    wire N__3141;
    wire N__3138;
    wire N__3135;
    wire N__3132;
    wire N__3129;
    wire N__3126;
    wire N__3123;
    wire N__3120;
    wire N__3117;
    wire N__3114;
    wire N__3111;
    wire N__3108;
    wire N__3105;
    wire N__3102;
    wire N__3099;
    wire N__3096;
    wire N__3093;
    wire N__3090;
    wire N__3087;
    wire N__3086;
    wire N__3085;
    wire N__3080;
    wire N__3077;
    wire N__3072;
    wire N__3069;
    wire N__3068;
    wire N__3067;
    wire N__3062;
    wire N__3059;
    wire N__3054;
    wire N__3051;
    wire N__3050;
    wire N__3047;
    wire N__3044;
    wire N__3043;
    wire N__3038;
    wire N__3035;
    wire N__3030;
    wire N__3027;
    wire N__3026;
    wire N__3025;
    wire N__3020;
    wire N__3017;
    wire N__3012;
    wire N__3009;
    wire N__3006;
    wire N__3005;
    wire N__3002;
    wire N__2999;
    wire N__2994;
    wire N__2991;
    wire N__2988;
    wire N__2985;
    wire N__2982;
    wire N__2979;
    wire N__2976;
    wire N__2973;
    wire N__2970;
    wire N__2967;
    wire N__2964;
    wire N__2961;
    wire N__2958;
    wire N__2955;
    wire N__2952;
    wire N__2949;
    wire N__2946;
    wire N__2943;
    wire N__2940;
    wire N__2937;
    wire N__2934;
    wire N__2931;
    wire N__2928;
    wire N__2925;
    wire N__2922;
    wire N__2919;
    wire N__2916;
    wire N__2913;
    wire N__2910;
    wire N__2907;
    wire N__2904;
    wire N__2901;
    wire N__2898;
    wire N__2895;
    wire N__2892;
    wire N__2889;
    wire N__2886;
    wire N__2883;
    wire N__2880;
    wire N__2877;
    wire N__2874;
    wire N__2871;
    wire N__2868;
    wire N__2865;
    wire N__2862;
    wire N__2859;
    wire N__2856;
    wire N__2853;
    wire N__2850;
    wire N__2847;
    wire N__2844;
    wire N__2841;
    wire N__2838;
    wire N__2835;
    wire N__2832;
    wire N__2829;
    wire N__2826;
    wire N__2823;
    wire N__2820;
    wire N__2817;
    wire N__2814;
    wire N__2811;
    wire N__2808;
    wire N__2805;
    wire N__2802;
    wire N__2799;
    wire N__2796;
    wire N__2793;
    wire N__2790;
    wire N__2787;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire GNDG0;
    wire n2553_cascade_;
    wire LED_c;
    wire n2554;
    wire n26;
    wire bfn_14_21_0_;
    wire n25;
    wire n2294;
    wire n24;
    wire n2295;
    wire n23;
    wire n2296;
    wire n22;
    wire n2297;
    wire n21;
    wire n2298;
    wire n20;
    wire n2299;
    wire n19;
    wire n2300;
    wire n2301;
    wire n18;
    wire bfn_14_22_0_;
    wire n17;
    wire n2302;
    wire n16;
    wire n2303;
    wire n15;
    wire n2304;
    wire n14;
    wire n2305;
    wire n13;
    wire n2306;
    wire n12;
    wire n2307;
    wire n11;
    wire n2308;
    wire n2309;
    wire n10;
    wire bfn_14_23_0_;
    wire n9;
    wire n2310;
    wire n8_adj_409;
    wire n2311;
    wire n7;
    wire n2312;
    wire n6_adj_410;
    wire n2313;
    wire blink_counter_21;
    wire n2314;
    wire blink_counter_22;
    wire n2315;
    wire blink_counter_23;
    wire n2316;
    wire n2317;
    wire blink_counter_24;
    wire bfn_14_24_0_;
    wire n2318;
    wire blink_counter_25;
    wire n693_cascade_;
    wire bfn_17_21_0_;
    wire n2263;
    wire n2264;
    wire n2265;
    wire n2266;
    wire n2267;
    wire n2268;
    wire n2269;
    wire n2270;
    wire bfn_17_22_0_;
    wire n2271;
    wire n2272;
    wire n2273;
    wire n2274;
    wire n2275;
    wire n2276;
    wire n2277;
    wire n2278;
    wire bfn_17_23_0_;
    wire n2279;
    wire n2280;
    wire n2281;
    wire n2282;
    wire n2283;
    wire n2284;
    wire n2285;
    wire n2286;
    wire bfn_17_24_0_;
    wire n2287;
    wire n2288;
    wire n2289;
    wire n2290;
    wire n2291;
    wire n2292;
    wire n2293;
    wire bfn_18_17_0_;
    wire \eeprom.n2241 ;
    wire \eeprom.delay_counter_2 ;
    wire \eeprom.delay_counter_15_N_171_2 ;
    wire \eeprom.n2242 ;
    wire \eeprom.n2243 ;
    wire \eeprom.n2244 ;
    wire \eeprom.n2245 ;
    wire \eeprom.delay_counter_6 ;
    wire \eeprom.delay_counter_15_N_171_6 ;
    wire \eeprom.n2246 ;
    wire \eeprom.n2247 ;
    wire \eeprom.n2248 ;
    wire \eeprom.delay_counter_8 ;
    wire \eeprom.delay_counter_15_N_171_8 ;
    wire bfn_18_18_0_;
    wire \eeprom.n2249 ;
    wire \eeprom.n2250 ;
    wire \eeprom.n2251 ;
    wire \eeprom.delay_counter_12 ;
    wire \eeprom.delay_counter_15_N_171_12 ;
    wire \eeprom.n2252 ;
    wire \eeprom.n2253 ;
    wire \eeprom.n2254 ;
    wire \eeprom.n642 ;
    wire \eeprom.n2255 ;
    wire \eeprom.n14 ;
    wire \eeprom.n13_cascade_ ;
    wire \eeprom.n7_cascade_ ;
    wire \eeprom.delay_counter_15_N_171_1 ;
    wire \eeprom.delay_counter_1 ;
    wire \eeprom.delay_counter_15_N_171_0 ;
    wire \eeprom.delay_counter_0 ;
    wire \eeprom.delay_counter_15_N_171_5 ;
    wire \eeprom.delay_counter_5 ;
    wire \eeprom.delay_counter_15_N_171_10 ;
    wire \eeprom.delay_counter_10 ;
    wire \eeprom.delay_counter_15_N_171_4 ;
    wire \eeprom.delay_counter_4 ;
    wire n324;
    wire \eeprom.n1500 ;
    wire n6_adj_405_cascade_;
    wire n41;
    wire \eeprom.n1018 ;
    wire n2483_cascade_;
    wire \eeprom.n2453 ;
    wire n1568_cascade_;
    wire state_1;
    wire n1568;
    wire delay_counter_7;
    wire delay_counter_8;
    wire delay_counter_1;
    wire delay_counter_4;
    wire delay_counter_10;
    wire delay_counter_12;
    wire delay_counter_11;
    wire delay_counter_13;
    wire n2512_cascade_;
    wire delay_counter_16;
    wire delay_counter_18;
    wire n2495_cascade_;
    wire delay_counter_19;
    wire delay_counter_9;
    wire delay_counter_6;
    wire delay_counter_3;
    wire delay_counter_0;
    wire delay_counter_17;
    wire delay_counter_15;
    wire delay_counter_14;
    wire n8;
    wire delay_counter_21;
    wire delay_counter_23;
    wire n6_adj_413;
    wire delay_counter_5;
    wire n16_adj_407;
    wire delay_counter_2;
    wire n17_adj_406;
    wire n2536;
    wire read_N;
    wire delay_counter_22;
    wire delay_counter_25;
    wire delay_counter_20;
    wire n8_adj_412;
    wire n9_adj_404;
    wire delay_counter_31;
    wire n9_adj_404_cascade_;
    wire addr_10__N_70;
    wire delay_counter_29;
    wire delay_counter_28;
    wire n10_adj_403;
    wire delay_counter_26;
    wire delay_counter_30;
    wire delay_counter_27;
    wire delay_counter_24;
    wire n14_adj_401;
    wire \eeprom.delay_counter_15_N_171_7 ;
    wire \eeprom.delay_counter_15_N_171_3 ;
    wire \eeprom.delay_counter_3 ;
    wire \eeprom.delay_counter_15_N_171_11 ;
    wire \eeprom.delay_counter_15_N_171_9 ;
    wire \eeprom.delay_counter_11 ;
    wire \eeprom.delay_counter_7 ;
    wire \eeprom.n6_cascade_ ;
    wire \eeprom.delay_counter_9 ;
    wire \eeprom.n8 ;
    wire \eeprom.delay_counter_15_N_171_15 ;
    wire \eeprom.delay_counter_15 ;
    wire \eeprom.delay_counter_15_N_171_14 ;
    wire \eeprom.delay_counter_14 ;
    wire state_0;
    wire \eeprom.n1601 ;
    wire \eeprom.delay_counter_15_N_171_13 ;
    wire \eeprom.delay_counter_13 ;
    wire \INVeeprom.i2c.write_enable_132C_net ;
    wire n11_adj_399_cascade_;
    wire \eeprom.i2c.n1669 ;
    wire \eeprom.i2c.n37_cascade_ ;
    wire \eeprom.i2c.n33 ;
    wire \eeprom.i2c.n39_cascade_ ;
    wire \eeprom.i2c.n1027 ;
    wire \eeprom.i2c.n11_adj_379 ;
    wire \INVeeprom.i2c.sda_out_133C_net ;
    wire \eeprom.i2c.n6_cascade_ ;
    wire \eeprom.i2c.counter2_7__N_256_cascade_ ;
    wire \eeprom.i2c.n1580 ;
    wire rw;
    wire n1835_cascade_;
    wire n2569;
    wire n949_cascade_;
    wire n949;
    wire n2547_cascade_;
    wire \eeprom.i2c.n2574_cascade_ ;
    wire \eeprom.i2c.n2557 ;
    wire \eeprom.enable ;
    wire n2538_cascade_;
    wire n4_adj_411_cascade_;
    wire n1835;
    wire n2507_cascade_;
    wire n10_adj_394;
    wire saved_addr_0;
    wire n11_adj_399;
    wire n2566;
    wire \eeprom.i2c.n39 ;
    wire \eeprom.i2c.n2406 ;
    wire \eeprom.i2c.n37 ;
    wire \eeprom.i2c.n1051_cascade_ ;
    wire \eeprom.i2c.n13 ;
    wire sda_out;
    wire sda_enable;
    wire state_7_N_285_3_cascade_;
    wire \eeprom.i2c.n2475 ;
    wire \eeprom.i2c.n2475_cascade_ ;
    wire \eeprom.i2c.n9 ;
    wire \eeprom.i2c.counter2_0 ;
    wire bfn_21_18_0_;
    wire \eeprom.i2c.counter2_1 ;
    wire \eeprom.i2c.n2319 ;
    wire \eeprom.i2c.counter2_2 ;
    wire \eeprom.i2c.n2320 ;
    wire \eeprom.i2c.counter2_3 ;
    wire \eeprom.i2c.n2321 ;
    wire \eeprom.i2c.n2322 ;
    wire \eeprom.i2c.counter2_4 ;
    wire CLK_N;
    wire \eeprom.i2c.counter2_7__N_256 ;
    wire n306;
    wire n10_adj_398_cascade_;
    wire state_7_N_269_0;
    wire n2460_cascade_;
    wire n2560;
    wire n308;
    wire n320;
    wire n318;
    wire n1817;
    wire \eeprom.i2c.n12_cascade_ ;
    wire n4_adj_408;
    wire \eeprom.i2c.n942 ;
    wire n10_adj_398;
    wire n11_adj_400;
    wire \eeprom.i2c.n942_cascade_ ;
    wire n1532;
    wire \eeprom.i2c.counter_0 ;
    wire bfn_21_22_0_;
    wire \eeprom.i2c.n2256 ;
    wire \eeprom.i2c.n2257 ;
    wire \eeprom.i2c.counter_3 ;
    wire \eeprom.i2c.n2258 ;
    wire \eeprom.i2c.counter_4 ;
    wire \eeprom.i2c.n2259 ;
    wire \eeprom.i2c.counter_5 ;
    wire \eeprom.i2c.n2260 ;
    wire \eeprom.i2c.counter_6 ;
    wire \eeprom.i2c.n2261 ;
    wire \eeprom.i2c.n2262 ;
    wire \eeprom.i2c.counter_7 ;
    wire \eeprom.i2c.n1548 ;
    wire \eeprom.i2c.n1655 ;
    wire CONSTANT_ONE_NET;
    wire n15_adj_393;
    wire \eeprom.i2c.n10_cascade_ ;
    wire \INVeeprom.i2c.i2c_scl_enable_124C_net ;
    wire state_2;
    wire state_0_adj_397;
    wire state_1_adj_396;
    wire state_3;
    wire n1826;
    wire n314;
    wire n1518;
    wire n4_adj_395_cascade_;
    wire n310;
    wire n4_adj_395;
    wire n312;
    wire \eeprom.i2c.counter_1 ;
    wire \eeprom.i2c.counter_2 ;
    wire n4;
    wire n1523;
    wire n4_cascade_;
    wire state_7_N_285_3;
    wire n316;
    wire scl_enable;
    wire \eeprom.i2c.i2c_clk ;
    wire scl_c;
    wire _gnd_net_;

    defparam CS_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CS_CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CS_CLK_pad_iopad (
            .OE(N__6589),
            .DIN(N__6588),
            .DOUT(N__6587),
            .PACKAGEPIN(CS_CLK));
    defparam CS_CLK_pad_preio.PIN_TYPE=6'b011001;
    defparam CS_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CS_CLK_pad_preio (
            .PADOEN(N__6589),
            .PADOUT(N__6588),
            .PADIN(N__6587),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam CS_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CS_pad_iopad.PULLUP=1'b0;
    IO_PAD CS_pad_iopad (
            .OE(N__6580),
            .DIN(N__6579),
            .DOUT(N__6578),
            .PACKAGEPIN(CS));
    defparam CS_pad_preio.PIN_TYPE=6'b011001;
    defparam CS_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CS_pad_preio (
            .PADOEN(N__6580),
            .PADOUT(N__6579),
            .PADIN(N__6578),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam DE_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DE_pad_iopad.PULLUP=1'b0;
    IO_PAD DE_pad_iopad (
            .OE(N__6571),
            .DIN(N__6570),
            .DOUT(N__6569),
            .PACKAGEPIN(DE));
    defparam DE_pad_preio.PIN_TYPE=6'b011001;
    defparam DE_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DE_pad_preio (
            .PADOEN(N__6571),
            .PADOUT(N__6570),
            .PADIN(N__6569),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHA_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHA_pad_iopad.PULLUP=1'b0;
    IO_PAD INHA_pad_iopad (
            .OE(N__6562),
            .DIN(N__6561),
            .DOUT(N__6560),
            .PACKAGEPIN(INHA));
    defparam INHA_pad_preio.PIN_TYPE=6'b011001;
    defparam INHA_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHA_pad_preio (
            .PADOEN(N__6562),
            .PADOUT(N__6561),
            .PADIN(N__6560),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHB_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHB_pad_iopad.PULLUP=1'b0;
    IO_PAD INHB_pad_iopad (
            .OE(N__6553),
            .DIN(N__6552),
            .DOUT(N__6551),
            .PACKAGEPIN(INHB));
    defparam INHB_pad_preio.PIN_TYPE=6'b011001;
    defparam INHB_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHB_pad_preio (
            .PADOEN(N__6553),
            .PADOUT(N__6552),
            .PADIN(N__6551),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHC_pad_iopad.PULLUP=1'b0;
    IO_PAD INHC_pad_iopad (
            .OE(N__6544),
            .DIN(N__6543),
            .DOUT(N__6542),
            .PACKAGEPIN(INHC));
    defparam INHC_pad_preio.PIN_TYPE=6'b011001;
    defparam INHC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHC_pad_preio (
            .PADOEN(N__6544),
            .PADOUT(N__6543),
            .PADIN(N__6542),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLA_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLA_pad_iopad.PULLUP=1'b0;
    IO_PAD INLA_pad_iopad (
            .OE(N__6535),
            .DIN(N__6534),
            .DOUT(N__6533),
            .PACKAGEPIN(INLA));
    defparam INLA_pad_preio.PIN_TYPE=6'b011001;
    defparam INLA_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLA_pad_preio (
            .PADOEN(N__6535),
            .PADOUT(N__6534),
            .PADIN(N__6533),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLB_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLB_pad_iopad.PULLUP=1'b0;
    IO_PAD INLB_pad_iopad (
            .OE(N__6526),
            .DIN(N__6525),
            .DOUT(N__6524),
            .PACKAGEPIN(INLB));
    defparam INLB_pad_preio.PIN_TYPE=6'b011001;
    defparam INLB_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLB_pad_preio (
            .PADOEN(N__6526),
            .PADOUT(N__6525),
            .PADIN(N__6524),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLC_pad_iopad.PULLUP=1'b0;
    IO_PAD INLC_pad_iopad (
            .OE(N__6517),
            .DIN(N__6516),
            .DOUT(N__6515),
            .PACKAGEPIN(INLC));
    defparam INLC_pad_preio.PIN_TYPE=6'b011001;
    defparam INLC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLC_pad_preio (
            .PADOEN(N__6517),
            .PADOUT(N__6516),
            .PADIN(N__6515),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__6508),
            .DIN(N__6507),
            .DOUT(N__6506),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__6508),
            .PADOUT(N__6507),
            .PADIN(N__6506),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__2838),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam NEOPXL_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam NEOPXL_pad_iopad.PULLUP=1'b0;
    IO_PAD NEOPXL_pad_iopad (
            .OE(N__6499),
            .DIN(N__6498),
            .DOUT(N__6497),
            .PACKAGEPIN(NEOPXL));
    defparam NEOPXL_pad_preio.PIN_TYPE=6'b011001;
    defparam NEOPXL_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO NEOPXL_pad_preio (
            .PADOEN(N__6499),
            .PADOUT(N__6498),
            .PADIN(N__6497),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam TX_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TX_pad_iopad.PULLUP=1'b0;
    IO_PAD TX_pad_iopad (
            .OE(N__6490),
            .DIN(N__6489),
            .DOUT(N__6488),
            .PACKAGEPIN(TX));
    defparam TX_pad_preio.PIN_TYPE=6'b011001;
    defparam TX_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO TX_pad_preio (
            .PADOEN(N__6490),
            .PADOUT(N__6489),
            .PADIN(N__6488),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__6481),
            .DIN(N__6480),
            .DOUT(N__6479),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__6481),
            .PADOUT(N__6480),
            .PADIN(N__6479),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam scl_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam scl_output_iopad.PULLUP=1'b1;
    IO_PAD scl_output_iopad (
            .OE(N__6472),
            .DIN(N__6471),
            .DOUT(N__6470),
            .PACKAGEPIN(SCL));
    defparam scl_output_preio.PIN_TYPE=6'b101001;
    defparam scl_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO scl_output_preio (
            .PADOEN(N__6472),
            .PADOUT(N__6471),
            .PADIN(N__6470),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__6063),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__6207));
    defparam sda_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam sda_output_iopad.PULLUP=1'b1;
    IO_PAD sda_output_iopad (
            .OE(N__6463),
            .DIN(N__6462),
            .DOUT(N__6461),
            .PACKAGEPIN(SDA));
    defparam sda_output_preio.PIN_TYPE=6'b101001;
    defparam sda_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO sda_output_preio (
            .PADOEN(N__6463),
            .PADOUT(N__6462),
            .PADIN(N__6461),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__6282),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__4941));
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__6454),
            .DIN(N__6453),
            .DOUT(N__6452),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__6454),
            .PADOUT(N__6453),
            .PADIN(N__6452),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__1455 (
            .O(N__6435),
            .I(N__6428));
    InMux I__1454 (
            .O(N__6434),
            .I(N__6428));
    InMux I__1453 (
            .O(N__6433),
            .I(N__6425));
    LocalMux I__1452 (
            .O(N__6428),
            .I(N__6421));
    LocalMux I__1451 (
            .O(N__6425),
            .I(N__6418));
    InMux I__1450 (
            .O(N__6424),
            .I(N__6415));
    Odrv4 I__1449 (
            .O(N__6421),
            .I(n1518));
    Odrv4 I__1448 (
            .O(N__6418),
            .I(n1518));
    LocalMux I__1447 (
            .O(N__6415),
            .I(n1518));
    CascadeMux I__1446 (
            .O(N__6408),
            .I(n4_adj_395_cascade_));
    InMux I__1445 (
            .O(N__6405),
            .I(N__6402));
    LocalMux I__1444 (
            .O(N__6402),
            .I(n310));
    InMux I__1443 (
            .O(N__6399),
            .I(N__6396));
    LocalMux I__1442 (
            .O(N__6396),
            .I(n4_adj_395));
    CascadeMux I__1441 (
            .O(N__6393),
            .I(N__6390));
    InMux I__1440 (
            .O(N__6390),
            .I(N__6387));
    LocalMux I__1439 (
            .O(N__6387),
            .I(n312));
    InMux I__1438 (
            .O(N__6384),
            .I(N__6374));
    InMux I__1437 (
            .O(N__6383),
            .I(N__6374));
    InMux I__1436 (
            .O(N__6382),
            .I(N__6371));
    InMux I__1435 (
            .O(N__6381),
            .I(N__6366));
    InMux I__1434 (
            .O(N__6380),
            .I(N__6366));
    InMux I__1433 (
            .O(N__6379),
            .I(N__6363));
    LocalMux I__1432 (
            .O(N__6374),
            .I(\eeprom.i2c.counter_1 ));
    LocalMux I__1431 (
            .O(N__6371),
            .I(\eeprom.i2c.counter_1 ));
    LocalMux I__1430 (
            .O(N__6366),
            .I(\eeprom.i2c.counter_1 ));
    LocalMux I__1429 (
            .O(N__6363),
            .I(\eeprom.i2c.counter_1 ));
    CascadeMux I__1428 (
            .O(N__6354),
            .I(N__6349));
    InMux I__1427 (
            .O(N__6353),
            .I(N__6341));
    InMux I__1426 (
            .O(N__6352),
            .I(N__6341));
    InMux I__1425 (
            .O(N__6349),
            .I(N__6338));
    InMux I__1424 (
            .O(N__6348),
            .I(N__6335));
    InMux I__1423 (
            .O(N__6347),
            .I(N__6332));
    InMux I__1422 (
            .O(N__6346),
            .I(N__6329));
    LocalMux I__1421 (
            .O(N__6341),
            .I(\eeprom.i2c.counter_2 ));
    LocalMux I__1420 (
            .O(N__6338),
            .I(\eeprom.i2c.counter_2 ));
    LocalMux I__1419 (
            .O(N__6335),
            .I(\eeprom.i2c.counter_2 ));
    LocalMux I__1418 (
            .O(N__6332),
            .I(\eeprom.i2c.counter_2 ));
    LocalMux I__1417 (
            .O(N__6329),
            .I(\eeprom.i2c.counter_2 ));
    InMux I__1416 (
            .O(N__6318),
            .I(N__6315));
    LocalMux I__1415 (
            .O(N__6315),
            .I(n4));
    CascadeMux I__1414 (
            .O(N__6312),
            .I(N__6307));
    InMux I__1413 (
            .O(N__6311),
            .I(N__6301));
    InMux I__1412 (
            .O(N__6310),
            .I(N__6301));
    InMux I__1411 (
            .O(N__6307),
            .I(N__6296));
    InMux I__1410 (
            .O(N__6306),
            .I(N__6296));
    LocalMux I__1409 (
            .O(N__6301),
            .I(N__6293));
    LocalMux I__1408 (
            .O(N__6296),
            .I(N__6290));
    Odrv4 I__1407 (
            .O(N__6293),
            .I(n1523));
    Odrv4 I__1406 (
            .O(N__6290),
            .I(n1523));
    CascadeMux I__1405 (
            .O(N__6285),
            .I(n4_cascade_));
    IoInMux I__1404 (
            .O(N__6282),
            .I(N__6279));
    LocalMux I__1403 (
            .O(N__6279),
            .I(N__6276));
    Span4Mux_s0_h I__1402 (
            .O(N__6276),
            .I(N__6273));
    Sp12to4 I__1401 (
            .O(N__6273),
            .I(N__6270));
    Span12Mux_v I__1400 (
            .O(N__6270),
            .I(N__6262));
    InMux I__1399 (
            .O(N__6269),
            .I(N__6259));
    InMux I__1398 (
            .O(N__6268),
            .I(N__6247));
    InMux I__1397 (
            .O(N__6267),
            .I(N__6247));
    InMux I__1396 (
            .O(N__6266),
            .I(N__6247));
    InMux I__1395 (
            .O(N__6265),
            .I(N__6247));
    Span12Mux_h I__1394 (
            .O(N__6262),
            .I(N__6242));
    LocalMux I__1393 (
            .O(N__6259),
            .I(N__6239));
    InMux I__1392 (
            .O(N__6258),
            .I(N__6232));
    InMux I__1391 (
            .O(N__6257),
            .I(N__6232));
    InMux I__1390 (
            .O(N__6256),
            .I(N__6232));
    LocalMux I__1389 (
            .O(N__6247),
            .I(N__6229));
    InMux I__1388 (
            .O(N__6246),
            .I(N__6224));
    InMux I__1387 (
            .O(N__6245),
            .I(N__6224));
    Odrv12 I__1386 (
            .O(N__6242),
            .I(state_7_N_285_3));
    Odrv4 I__1385 (
            .O(N__6239),
            .I(state_7_N_285_3));
    LocalMux I__1384 (
            .O(N__6232),
            .I(state_7_N_285_3));
    Odrv4 I__1383 (
            .O(N__6229),
            .I(state_7_N_285_3));
    LocalMux I__1382 (
            .O(N__6224),
            .I(state_7_N_285_3));
    InMux I__1381 (
            .O(N__6213),
            .I(N__6210));
    LocalMux I__1380 (
            .O(N__6210),
            .I(n316));
    IoInMux I__1379 (
            .O(N__6207),
            .I(N__6204));
    LocalMux I__1378 (
            .O(N__6204),
            .I(N__6201));
    IoSpan4Mux I__1377 (
            .O(N__6201),
            .I(N__6198));
    Span4Mux_s2_h I__1376 (
            .O(N__6198),
            .I(N__6195));
    Span4Mux_h I__1375 (
            .O(N__6195),
            .I(N__6191));
    InMux I__1374 (
            .O(N__6194),
            .I(N__6188));
    Odrv4 I__1373 (
            .O(N__6191),
            .I(scl_enable));
    LocalMux I__1372 (
            .O(N__6188),
            .I(scl_enable));
    ClkMux I__1371 (
            .O(N__6183),
            .I(N__6177));
    InMux I__1370 (
            .O(N__6182),
            .I(N__6174));
    ClkMux I__1369 (
            .O(N__6181),
            .I(N__6171));
    ClkMux I__1368 (
            .O(N__6180),
            .I(N__6166));
    LocalMux I__1367 (
            .O(N__6177),
            .I(N__6162));
    LocalMux I__1366 (
            .O(N__6174),
            .I(N__6157));
    LocalMux I__1365 (
            .O(N__6171),
            .I(N__6157));
    ClkMux I__1364 (
            .O(N__6170),
            .I(N__6154));
    ClkMux I__1363 (
            .O(N__6169),
            .I(N__6150));
    LocalMux I__1362 (
            .O(N__6166),
            .I(N__6147));
    ClkMux I__1361 (
            .O(N__6165),
            .I(N__6144));
    Span4Mux_v I__1360 (
            .O(N__6162),
            .I(N__6137));
    Span4Mux_v I__1359 (
            .O(N__6157),
            .I(N__6137));
    LocalMux I__1358 (
            .O(N__6154),
            .I(N__6137));
    ClkMux I__1357 (
            .O(N__6153),
            .I(N__6134));
    LocalMux I__1356 (
            .O(N__6150),
            .I(N__6131));
    Span4Mux_v I__1355 (
            .O(N__6147),
            .I(N__6126));
    LocalMux I__1354 (
            .O(N__6144),
            .I(N__6123));
    Span4Mux_h I__1353 (
            .O(N__6137),
            .I(N__6118));
    LocalMux I__1352 (
            .O(N__6134),
            .I(N__6118));
    Span4Mux_h I__1351 (
            .O(N__6131),
            .I(N__6114));
    ClkMux I__1350 (
            .O(N__6130),
            .I(N__6111));
    ClkMux I__1349 (
            .O(N__6129),
            .I(N__6107));
    Span4Mux_h I__1348 (
            .O(N__6126),
            .I(N__6103));
    Span4Mux_h I__1347 (
            .O(N__6123),
            .I(N__6100));
    Sp12to4 I__1346 (
            .O(N__6118),
            .I(N__6097));
    InMux I__1345 (
            .O(N__6117),
            .I(N__6094));
    Span4Mux_v I__1344 (
            .O(N__6114),
            .I(N__6089));
    LocalMux I__1343 (
            .O(N__6111),
            .I(N__6089));
    InMux I__1342 (
            .O(N__6110),
            .I(N__6086));
    LocalMux I__1341 (
            .O(N__6107),
            .I(N__6083));
    InMux I__1340 (
            .O(N__6106),
            .I(N__6080));
    Odrv4 I__1339 (
            .O(N__6103),
            .I(\eeprom.i2c.i2c_clk ));
    Odrv4 I__1338 (
            .O(N__6100),
            .I(\eeprom.i2c.i2c_clk ));
    Odrv12 I__1337 (
            .O(N__6097),
            .I(\eeprom.i2c.i2c_clk ));
    LocalMux I__1336 (
            .O(N__6094),
            .I(\eeprom.i2c.i2c_clk ));
    Odrv4 I__1335 (
            .O(N__6089),
            .I(\eeprom.i2c.i2c_clk ));
    LocalMux I__1334 (
            .O(N__6086),
            .I(\eeprom.i2c.i2c_clk ));
    Odrv4 I__1333 (
            .O(N__6083),
            .I(\eeprom.i2c.i2c_clk ));
    LocalMux I__1332 (
            .O(N__6080),
            .I(\eeprom.i2c.i2c_clk ));
    IoInMux I__1331 (
            .O(N__6063),
            .I(N__6060));
    LocalMux I__1330 (
            .O(N__6060),
            .I(N__6057));
    Sp12to4 I__1329 (
            .O(N__6057),
            .I(N__6054));
    Odrv12 I__1328 (
            .O(N__6054),
            .I(scl_c));
    InMux I__1327 (
            .O(N__6051),
            .I(N__6047));
    InMux I__1326 (
            .O(N__6050),
            .I(N__6044));
    LocalMux I__1325 (
            .O(N__6047),
            .I(\eeprom.i2c.counter_5 ));
    LocalMux I__1324 (
            .O(N__6044),
            .I(\eeprom.i2c.counter_5 ));
    InMux I__1323 (
            .O(N__6039),
            .I(\eeprom.i2c.n2260 ));
    CascadeMux I__1322 (
            .O(N__6036),
            .I(N__6033));
    InMux I__1321 (
            .O(N__6033),
            .I(N__6029));
    InMux I__1320 (
            .O(N__6032),
            .I(N__6026));
    LocalMux I__1319 (
            .O(N__6029),
            .I(\eeprom.i2c.counter_6 ));
    LocalMux I__1318 (
            .O(N__6026),
            .I(\eeprom.i2c.counter_6 ));
    InMux I__1317 (
            .O(N__6021),
            .I(\eeprom.i2c.n2261 ));
    InMux I__1316 (
            .O(N__6018),
            .I(\eeprom.i2c.n2262 ));
    InMux I__1315 (
            .O(N__6015),
            .I(N__6011));
    InMux I__1314 (
            .O(N__6014),
            .I(N__6008));
    LocalMux I__1313 (
            .O(N__6011),
            .I(\eeprom.i2c.counter_7 ));
    LocalMux I__1312 (
            .O(N__6008),
            .I(\eeprom.i2c.counter_7 ));
    CEMux I__1311 (
            .O(N__6003),
            .I(N__6000));
    LocalMux I__1310 (
            .O(N__6000),
            .I(\eeprom.i2c.n1548 ));
    SRMux I__1309 (
            .O(N__5997),
            .I(N__5994));
    LocalMux I__1308 (
            .O(N__5994),
            .I(N__5991));
    Odrv4 I__1307 (
            .O(N__5991),
            .I(\eeprom.i2c.n1655 ));
    CascadeMux I__1306 (
            .O(N__5988),
            .I(N__5981));
    CascadeMux I__1305 (
            .O(N__5987),
            .I(N__5977));
    CascadeMux I__1304 (
            .O(N__5986),
            .I(N__5973));
    InMux I__1303 (
            .O(N__5985),
            .I(N__5958));
    InMux I__1302 (
            .O(N__5984),
            .I(N__5958));
    InMux I__1301 (
            .O(N__5981),
            .I(N__5958));
    InMux I__1300 (
            .O(N__5980),
            .I(N__5958));
    InMux I__1299 (
            .O(N__5977),
            .I(N__5958));
    InMux I__1298 (
            .O(N__5976),
            .I(N__5958));
    InMux I__1297 (
            .O(N__5973),
            .I(N__5958));
    LocalMux I__1296 (
            .O(N__5958),
            .I(N__5955));
    Odrv4 I__1295 (
            .O(N__5955),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__1294 (
            .O(N__5952),
            .I(N__5948));
    InMux I__1293 (
            .O(N__5951),
            .I(N__5939));
    InMux I__1292 (
            .O(N__5948),
            .I(N__5939));
    InMux I__1291 (
            .O(N__5947),
            .I(N__5936));
    CascadeMux I__1290 (
            .O(N__5946),
            .I(N__5933));
    CascadeMux I__1289 (
            .O(N__5945),
            .I(N__5930));
    CascadeMux I__1288 (
            .O(N__5944),
            .I(N__5926));
    LocalMux I__1287 (
            .O(N__5939),
            .I(N__5923));
    LocalMux I__1286 (
            .O(N__5936),
            .I(N__5920));
    InMux I__1285 (
            .O(N__5933),
            .I(N__5917));
    InMux I__1284 (
            .O(N__5930),
            .I(N__5910));
    InMux I__1283 (
            .O(N__5929),
            .I(N__5910));
    InMux I__1282 (
            .O(N__5926),
            .I(N__5910));
    Span4Mux_h I__1281 (
            .O(N__5923),
            .I(N__5905));
    Span4Mux_v I__1280 (
            .O(N__5920),
            .I(N__5902));
    LocalMux I__1279 (
            .O(N__5917),
            .I(N__5897));
    LocalMux I__1278 (
            .O(N__5910),
            .I(N__5897));
    InMux I__1277 (
            .O(N__5909),
            .I(N__5894));
    InMux I__1276 (
            .O(N__5908),
            .I(N__5891));
    Odrv4 I__1275 (
            .O(N__5905),
            .I(n15_adj_393));
    Odrv4 I__1274 (
            .O(N__5902),
            .I(n15_adj_393));
    Odrv12 I__1273 (
            .O(N__5897),
            .I(n15_adj_393));
    LocalMux I__1272 (
            .O(N__5894),
            .I(n15_adj_393));
    LocalMux I__1271 (
            .O(N__5891),
            .I(n15_adj_393));
    CascadeMux I__1270 (
            .O(N__5880),
            .I(\eeprom.i2c.n10_cascade_ ));
    InMux I__1269 (
            .O(N__5877),
            .I(N__5867));
    InMux I__1268 (
            .O(N__5876),
            .I(N__5862));
    InMux I__1267 (
            .O(N__5875),
            .I(N__5862));
    InMux I__1266 (
            .O(N__5874),
            .I(N__5854));
    InMux I__1265 (
            .O(N__5873),
            .I(N__5845));
    InMux I__1264 (
            .O(N__5872),
            .I(N__5845));
    InMux I__1263 (
            .O(N__5871),
            .I(N__5845));
    InMux I__1262 (
            .O(N__5870),
            .I(N__5845));
    LocalMux I__1261 (
            .O(N__5867),
            .I(N__5834));
    LocalMux I__1260 (
            .O(N__5862),
            .I(N__5831));
    InMux I__1259 (
            .O(N__5861),
            .I(N__5828));
    InMux I__1258 (
            .O(N__5860),
            .I(N__5825));
    InMux I__1257 (
            .O(N__5859),
            .I(N__5818));
    InMux I__1256 (
            .O(N__5858),
            .I(N__5818));
    InMux I__1255 (
            .O(N__5857),
            .I(N__5818));
    LocalMux I__1254 (
            .O(N__5854),
            .I(N__5813));
    LocalMux I__1253 (
            .O(N__5845),
            .I(N__5813));
    InMux I__1252 (
            .O(N__5844),
            .I(N__5804));
    InMux I__1251 (
            .O(N__5843),
            .I(N__5804));
    InMux I__1250 (
            .O(N__5842),
            .I(N__5804));
    InMux I__1249 (
            .O(N__5841),
            .I(N__5804));
    InMux I__1248 (
            .O(N__5840),
            .I(N__5795));
    InMux I__1247 (
            .O(N__5839),
            .I(N__5795));
    InMux I__1246 (
            .O(N__5838),
            .I(N__5795));
    InMux I__1245 (
            .O(N__5837),
            .I(N__5795));
    Odrv4 I__1244 (
            .O(N__5834),
            .I(state_2));
    Odrv4 I__1243 (
            .O(N__5831),
            .I(state_2));
    LocalMux I__1242 (
            .O(N__5828),
            .I(state_2));
    LocalMux I__1241 (
            .O(N__5825),
            .I(state_2));
    LocalMux I__1240 (
            .O(N__5818),
            .I(state_2));
    Odrv4 I__1239 (
            .O(N__5813),
            .I(state_2));
    LocalMux I__1238 (
            .O(N__5804),
            .I(state_2));
    LocalMux I__1237 (
            .O(N__5795),
            .I(state_2));
    CascadeMux I__1236 (
            .O(N__5778),
            .I(N__5773));
    InMux I__1235 (
            .O(N__5777),
            .I(N__5762));
    InMux I__1234 (
            .O(N__5776),
            .I(N__5751));
    InMux I__1233 (
            .O(N__5773),
            .I(N__5751));
    InMux I__1232 (
            .O(N__5772),
            .I(N__5751));
    InMux I__1231 (
            .O(N__5771),
            .I(N__5746));
    InMux I__1230 (
            .O(N__5770),
            .I(N__5746));
    InMux I__1229 (
            .O(N__5769),
            .I(N__5738));
    InMux I__1228 (
            .O(N__5768),
            .I(N__5735));
    InMux I__1227 (
            .O(N__5767),
            .I(N__5728));
    InMux I__1226 (
            .O(N__5766),
            .I(N__5728));
    InMux I__1225 (
            .O(N__5765),
            .I(N__5728));
    LocalMux I__1224 (
            .O(N__5762),
            .I(N__5721));
    InMux I__1223 (
            .O(N__5761),
            .I(N__5718));
    InMux I__1222 (
            .O(N__5760),
            .I(N__5715));
    InMux I__1221 (
            .O(N__5759),
            .I(N__5710));
    InMux I__1220 (
            .O(N__5758),
            .I(N__5710));
    LocalMux I__1219 (
            .O(N__5751),
            .I(N__5705));
    LocalMux I__1218 (
            .O(N__5746),
            .I(N__5705));
    InMux I__1217 (
            .O(N__5745),
            .I(N__5694));
    InMux I__1216 (
            .O(N__5744),
            .I(N__5694));
    InMux I__1215 (
            .O(N__5743),
            .I(N__5694));
    InMux I__1214 (
            .O(N__5742),
            .I(N__5694));
    InMux I__1213 (
            .O(N__5741),
            .I(N__5694));
    LocalMux I__1212 (
            .O(N__5738),
            .I(N__5687));
    LocalMux I__1211 (
            .O(N__5735),
            .I(N__5687));
    LocalMux I__1210 (
            .O(N__5728),
            .I(N__5687));
    InMux I__1209 (
            .O(N__5727),
            .I(N__5678));
    InMux I__1208 (
            .O(N__5726),
            .I(N__5678));
    InMux I__1207 (
            .O(N__5725),
            .I(N__5678));
    InMux I__1206 (
            .O(N__5724),
            .I(N__5678));
    Odrv4 I__1205 (
            .O(N__5721),
            .I(state_0_adj_397));
    LocalMux I__1204 (
            .O(N__5718),
            .I(state_0_adj_397));
    LocalMux I__1203 (
            .O(N__5715),
            .I(state_0_adj_397));
    LocalMux I__1202 (
            .O(N__5710),
            .I(state_0_adj_397));
    Odrv4 I__1201 (
            .O(N__5705),
            .I(state_0_adj_397));
    LocalMux I__1200 (
            .O(N__5694),
            .I(state_0_adj_397));
    Odrv4 I__1199 (
            .O(N__5687),
            .I(state_0_adj_397));
    LocalMux I__1198 (
            .O(N__5678),
            .I(state_0_adj_397));
    InMux I__1197 (
            .O(N__5661),
            .I(N__5657));
    CascadeMux I__1196 (
            .O(N__5660),
            .I(N__5654));
    LocalMux I__1195 (
            .O(N__5657),
            .I(N__5645));
    InMux I__1194 (
            .O(N__5654),
            .I(N__5640));
    InMux I__1193 (
            .O(N__5653),
            .I(N__5640));
    InMux I__1192 (
            .O(N__5652),
            .I(N__5632));
    InMux I__1191 (
            .O(N__5651),
            .I(N__5632));
    CascadeMux I__1190 (
            .O(N__5650),
            .I(N__5626));
    CascadeMux I__1189 (
            .O(N__5649),
            .I(N__5620));
    CascadeMux I__1188 (
            .O(N__5648),
            .I(N__5612));
    Span4Mux_h I__1187 (
            .O(N__5645),
            .I(N__5607));
    LocalMux I__1186 (
            .O(N__5640),
            .I(N__5607));
    InMux I__1185 (
            .O(N__5639),
            .I(N__5600));
    InMux I__1184 (
            .O(N__5638),
            .I(N__5600));
    InMux I__1183 (
            .O(N__5637),
            .I(N__5600));
    LocalMux I__1182 (
            .O(N__5632),
            .I(N__5597));
    InMux I__1181 (
            .O(N__5631),
            .I(N__5588));
    InMux I__1180 (
            .O(N__5630),
            .I(N__5588));
    InMux I__1179 (
            .O(N__5629),
            .I(N__5588));
    InMux I__1178 (
            .O(N__5626),
            .I(N__5588));
    InMux I__1177 (
            .O(N__5625),
            .I(N__5581));
    InMux I__1176 (
            .O(N__5624),
            .I(N__5581));
    InMux I__1175 (
            .O(N__5623),
            .I(N__5581));
    InMux I__1174 (
            .O(N__5620),
            .I(N__5578));
    InMux I__1173 (
            .O(N__5619),
            .I(N__5565));
    InMux I__1172 (
            .O(N__5618),
            .I(N__5565));
    InMux I__1171 (
            .O(N__5617),
            .I(N__5565));
    InMux I__1170 (
            .O(N__5616),
            .I(N__5565));
    InMux I__1169 (
            .O(N__5615),
            .I(N__5565));
    InMux I__1168 (
            .O(N__5612),
            .I(N__5565));
    Odrv4 I__1167 (
            .O(N__5607),
            .I(state_1_adj_396));
    LocalMux I__1166 (
            .O(N__5600),
            .I(state_1_adj_396));
    Odrv4 I__1165 (
            .O(N__5597),
            .I(state_1_adj_396));
    LocalMux I__1164 (
            .O(N__5588),
            .I(state_1_adj_396));
    LocalMux I__1163 (
            .O(N__5581),
            .I(state_1_adj_396));
    LocalMux I__1162 (
            .O(N__5578),
            .I(state_1_adj_396));
    LocalMux I__1161 (
            .O(N__5565),
            .I(state_1_adj_396));
    InMux I__1160 (
            .O(N__5550),
            .I(N__5545));
    InMux I__1159 (
            .O(N__5549),
            .I(N__5540));
    InMux I__1158 (
            .O(N__5548),
            .I(N__5540));
    LocalMux I__1157 (
            .O(N__5545),
            .I(N__5529));
    LocalMux I__1156 (
            .O(N__5540),
            .I(N__5526));
    CascadeMux I__1155 (
            .O(N__5539),
            .I(N__5518));
    InMux I__1154 (
            .O(N__5538),
            .I(N__5510));
    InMux I__1153 (
            .O(N__5537),
            .I(N__5510));
    InMux I__1152 (
            .O(N__5536),
            .I(N__5505));
    InMux I__1151 (
            .O(N__5535),
            .I(N__5505));
    InMux I__1150 (
            .O(N__5534),
            .I(N__5498));
    InMux I__1149 (
            .O(N__5533),
            .I(N__5498));
    InMux I__1148 (
            .O(N__5532),
            .I(N__5498));
    Span4Mux_h I__1147 (
            .O(N__5529),
            .I(N__5493));
    Span4Mux_h I__1146 (
            .O(N__5526),
            .I(N__5493));
    InMux I__1145 (
            .O(N__5525),
            .I(N__5490));
    InMux I__1144 (
            .O(N__5524),
            .I(N__5481));
    InMux I__1143 (
            .O(N__5523),
            .I(N__5481));
    InMux I__1142 (
            .O(N__5522),
            .I(N__5481));
    InMux I__1141 (
            .O(N__5521),
            .I(N__5481));
    InMux I__1140 (
            .O(N__5518),
            .I(N__5472));
    InMux I__1139 (
            .O(N__5517),
            .I(N__5472));
    InMux I__1138 (
            .O(N__5516),
            .I(N__5472));
    InMux I__1137 (
            .O(N__5515),
            .I(N__5472));
    LocalMux I__1136 (
            .O(N__5510),
            .I(state_3));
    LocalMux I__1135 (
            .O(N__5505),
            .I(state_3));
    LocalMux I__1134 (
            .O(N__5498),
            .I(state_3));
    Odrv4 I__1133 (
            .O(N__5493),
            .I(state_3));
    LocalMux I__1132 (
            .O(N__5490),
            .I(state_3));
    LocalMux I__1131 (
            .O(N__5481),
            .I(state_3));
    LocalMux I__1130 (
            .O(N__5472),
            .I(state_3));
    CascadeMux I__1129 (
            .O(N__5457),
            .I(N__5453));
    InMux I__1128 (
            .O(N__5456),
            .I(N__5450));
    InMux I__1127 (
            .O(N__5453),
            .I(N__5447));
    LocalMux I__1126 (
            .O(N__5450),
            .I(N__5442));
    LocalMux I__1125 (
            .O(N__5447),
            .I(N__5442));
    Odrv4 I__1124 (
            .O(N__5442),
            .I(n1826));
    CascadeMux I__1123 (
            .O(N__5439),
            .I(N__5436));
    InMux I__1122 (
            .O(N__5436),
            .I(N__5433));
    LocalMux I__1121 (
            .O(N__5433),
            .I(n314));
    InMux I__1120 (
            .O(N__5430),
            .I(N__5426));
    InMux I__1119 (
            .O(N__5429),
            .I(N__5423));
    LocalMux I__1118 (
            .O(N__5426),
            .I(n1817));
    LocalMux I__1117 (
            .O(N__5423),
            .I(n1817));
    CascadeMux I__1116 (
            .O(N__5418),
            .I(\eeprom.i2c.n12_cascade_ ));
    InMux I__1115 (
            .O(N__5415),
            .I(N__5406));
    InMux I__1114 (
            .O(N__5414),
            .I(N__5406));
    InMux I__1113 (
            .O(N__5413),
            .I(N__5406));
    LocalMux I__1112 (
            .O(N__5406),
            .I(n4_adj_408));
    InMux I__1111 (
            .O(N__5403),
            .I(N__5400));
    LocalMux I__1110 (
            .O(N__5400),
            .I(\eeprom.i2c.n942 ));
    CascadeMux I__1109 (
            .O(N__5397),
            .I(N__5393));
    InMux I__1108 (
            .O(N__5396),
            .I(N__5389));
    InMux I__1107 (
            .O(N__5393),
            .I(N__5386));
    InMux I__1106 (
            .O(N__5392),
            .I(N__5383));
    LocalMux I__1105 (
            .O(N__5389),
            .I(N__5380));
    LocalMux I__1104 (
            .O(N__5386),
            .I(n10_adj_398));
    LocalMux I__1103 (
            .O(N__5383),
            .I(n10_adj_398));
    Odrv4 I__1102 (
            .O(N__5380),
            .I(n10_adj_398));
    InMux I__1101 (
            .O(N__5373),
            .I(N__5369));
    InMux I__1100 (
            .O(N__5372),
            .I(N__5366));
    LocalMux I__1099 (
            .O(N__5369),
            .I(N__5363));
    LocalMux I__1098 (
            .O(N__5366),
            .I(n11_adj_400));
    Odrv4 I__1097 (
            .O(N__5363),
            .I(n11_adj_400));
    CascadeMux I__1096 (
            .O(N__5358),
            .I(\eeprom.i2c.n942_cascade_ ));
    InMux I__1095 (
            .O(N__5355),
            .I(N__5351));
    InMux I__1094 (
            .O(N__5354),
            .I(N__5348));
    LocalMux I__1093 (
            .O(N__5351),
            .I(n1532));
    LocalMux I__1092 (
            .O(N__5348),
            .I(n1532));
    InMux I__1091 (
            .O(N__5343),
            .I(N__5337));
    InMux I__1090 (
            .O(N__5342),
            .I(N__5337));
    LocalMux I__1089 (
            .O(N__5337),
            .I(N__5331));
    InMux I__1088 (
            .O(N__5336),
            .I(N__5328));
    InMux I__1087 (
            .O(N__5335),
            .I(N__5325));
    InMux I__1086 (
            .O(N__5334),
            .I(N__5322));
    Odrv4 I__1085 (
            .O(N__5331),
            .I(\eeprom.i2c.counter_0 ));
    LocalMux I__1084 (
            .O(N__5328),
            .I(\eeprom.i2c.counter_0 ));
    LocalMux I__1083 (
            .O(N__5325),
            .I(\eeprom.i2c.counter_0 ));
    LocalMux I__1082 (
            .O(N__5322),
            .I(\eeprom.i2c.counter_0 ));
    InMux I__1081 (
            .O(N__5313),
            .I(bfn_21_22_0_));
    InMux I__1080 (
            .O(N__5310),
            .I(\eeprom.i2c.n2256 ));
    InMux I__1079 (
            .O(N__5307),
            .I(\eeprom.i2c.n2257 ));
    InMux I__1078 (
            .O(N__5304),
            .I(N__5300));
    InMux I__1077 (
            .O(N__5303),
            .I(N__5297));
    LocalMux I__1076 (
            .O(N__5300),
            .I(\eeprom.i2c.counter_3 ));
    LocalMux I__1075 (
            .O(N__5297),
            .I(\eeprom.i2c.counter_3 ));
    InMux I__1074 (
            .O(N__5292),
            .I(\eeprom.i2c.n2258 ));
    CascadeMux I__1073 (
            .O(N__5289),
            .I(N__5285));
    CascadeMux I__1072 (
            .O(N__5288),
            .I(N__5282));
    InMux I__1071 (
            .O(N__5285),
            .I(N__5279));
    InMux I__1070 (
            .O(N__5282),
            .I(N__5276));
    LocalMux I__1069 (
            .O(N__5279),
            .I(\eeprom.i2c.counter_4 ));
    LocalMux I__1068 (
            .O(N__5276),
            .I(\eeprom.i2c.counter_4 ));
    InMux I__1067 (
            .O(N__5271),
            .I(\eeprom.i2c.n2259 ));
    CascadeMux I__1066 (
            .O(N__5268),
            .I(n10_adj_398_cascade_));
    InMux I__1065 (
            .O(N__5265),
            .I(N__5261));
    InMux I__1064 (
            .O(N__5264),
            .I(N__5258));
    LocalMux I__1063 (
            .O(N__5261),
            .I(state_7_N_269_0));
    LocalMux I__1062 (
            .O(N__5258),
            .I(state_7_N_269_0));
    CascadeMux I__1061 (
            .O(N__5253),
            .I(n2460_cascade_));
    InMux I__1060 (
            .O(N__5250),
            .I(N__5247));
    LocalMux I__1059 (
            .O(N__5247),
            .I(N__5244));
    Odrv4 I__1058 (
            .O(N__5244),
            .I(n2560));
    InMux I__1057 (
            .O(N__5241),
            .I(N__5238));
    LocalMux I__1056 (
            .O(N__5238),
            .I(n308));
    CascadeMux I__1055 (
            .O(N__5235),
            .I(N__5232));
    InMux I__1054 (
            .O(N__5232),
            .I(N__5229));
    LocalMux I__1053 (
            .O(N__5229),
            .I(n320));
    CascadeMux I__1052 (
            .O(N__5226),
            .I(N__5223));
    InMux I__1051 (
            .O(N__5223),
            .I(N__5220));
    LocalMux I__1050 (
            .O(N__5220),
            .I(n318));
    InMux I__1049 (
            .O(N__5217),
            .I(N__5214));
    LocalMux I__1048 (
            .O(N__5214),
            .I(\eeprom.i2c.n9 ));
    InMux I__1047 (
            .O(N__5211),
            .I(N__5207));
    InMux I__1046 (
            .O(N__5210),
            .I(N__5204));
    LocalMux I__1045 (
            .O(N__5207),
            .I(\eeprom.i2c.counter2_0 ));
    LocalMux I__1044 (
            .O(N__5204),
            .I(\eeprom.i2c.counter2_0 ));
    InMux I__1043 (
            .O(N__5199),
            .I(bfn_21_18_0_));
    InMux I__1042 (
            .O(N__5196),
            .I(N__5192));
    InMux I__1041 (
            .O(N__5195),
            .I(N__5189));
    LocalMux I__1040 (
            .O(N__5192),
            .I(\eeprom.i2c.counter2_1 ));
    LocalMux I__1039 (
            .O(N__5189),
            .I(\eeprom.i2c.counter2_1 ));
    InMux I__1038 (
            .O(N__5184),
            .I(\eeprom.i2c.n2319 ));
    InMux I__1037 (
            .O(N__5181),
            .I(N__5177));
    InMux I__1036 (
            .O(N__5180),
            .I(N__5174));
    LocalMux I__1035 (
            .O(N__5177),
            .I(\eeprom.i2c.counter2_2 ));
    LocalMux I__1034 (
            .O(N__5174),
            .I(\eeprom.i2c.counter2_2 ));
    InMux I__1033 (
            .O(N__5169),
            .I(\eeprom.i2c.n2320 ));
    InMux I__1032 (
            .O(N__5166),
            .I(N__5162));
    InMux I__1031 (
            .O(N__5165),
            .I(N__5159));
    LocalMux I__1030 (
            .O(N__5162),
            .I(\eeprom.i2c.counter2_3 ));
    LocalMux I__1029 (
            .O(N__5159),
            .I(\eeprom.i2c.counter2_3 ));
    InMux I__1028 (
            .O(N__5154),
            .I(\eeprom.i2c.n2321 ));
    InMux I__1027 (
            .O(N__5151),
            .I(\eeprom.i2c.n2322 ));
    InMux I__1026 (
            .O(N__5148),
            .I(N__5144));
    InMux I__1025 (
            .O(N__5147),
            .I(N__5141));
    LocalMux I__1024 (
            .O(N__5144),
            .I(\eeprom.i2c.counter2_4 ));
    LocalMux I__1023 (
            .O(N__5141),
            .I(\eeprom.i2c.counter2_4 ));
    ClkMux I__1022 (
            .O(N__5136),
            .I(N__5076));
    ClkMux I__1021 (
            .O(N__5135),
            .I(N__5076));
    ClkMux I__1020 (
            .O(N__5134),
            .I(N__5076));
    ClkMux I__1019 (
            .O(N__5133),
            .I(N__5076));
    ClkMux I__1018 (
            .O(N__5132),
            .I(N__5076));
    ClkMux I__1017 (
            .O(N__5131),
            .I(N__5076));
    ClkMux I__1016 (
            .O(N__5130),
            .I(N__5076));
    ClkMux I__1015 (
            .O(N__5129),
            .I(N__5076));
    ClkMux I__1014 (
            .O(N__5128),
            .I(N__5076));
    ClkMux I__1013 (
            .O(N__5127),
            .I(N__5076));
    ClkMux I__1012 (
            .O(N__5126),
            .I(N__5076));
    ClkMux I__1011 (
            .O(N__5125),
            .I(N__5076));
    ClkMux I__1010 (
            .O(N__5124),
            .I(N__5076));
    ClkMux I__1009 (
            .O(N__5123),
            .I(N__5076));
    ClkMux I__1008 (
            .O(N__5122),
            .I(N__5076));
    ClkMux I__1007 (
            .O(N__5121),
            .I(N__5076));
    ClkMux I__1006 (
            .O(N__5120),
            .I(N__5076));
    ClkMux I__1005 (
            .O(N__5119),
            .I(N__5076));
    ClkMux I__1004 (
            .O(N__5118),
            .I(N__5076));
    ClkMux I__1003 (
            .O(N__5117),
            .I(N__5076));
    GlobalMux I__1002 (
            .O(N__5076),
            .I(N__5073));
    gio2CtrlBuf I__1001 (
            .O(N__5073),
            .I(CLK_N));
    SRMux I__1000 (
            .O(N__5070),
            .I(N__5067));
    LocalMux I__999 (
            .O(N__5067),
            .I(N__5062));
    InMux I__998 (
            .O(N__5066),
            .I(N__5059));
    InMux I__997 (
            .O(N__5065),
            .I(N__5056));
    Odrv4 I__996 (
            .O(N__5062),
            .I(\eeprom.i2c.counter2_7__N_256 ));
    LocalMux I__995 (
            .O(N__5059),
            .I(\eeprom.i2c.counter2_7__N_256 ));
    LocalMux I__994 (
            .O(N__5056),
            .I(\eeprom.i2c.counter2_7__N_256 ));
    CascadeMux I__993 (
            .O(N__5049),
            .I(N__5046));
    InMux I__992 (
            .O(N__5046),
            .I(N__5043));
    LocalMux I__991 (
            .O(N__5043),
            .I(n306));
    InMux I__990 (
            .O(N__5040),
            .I(N__5035));
    InMux I__989 (
            .O(N__5039),
            .I(N__5030));
    InMux I__988 (
            .O(N__5038),
            .I(N__5030));
    LocalMux I__987 (
            .O(N__5035),
            .I(saved_addr_0));
    LocalMux I__986 (
            .O(N__5030),
            .I(saved_addr_0));
    CascadeMux I__985 (
            .O(N__5025),
            .I(N__5022));
    InMux I__984 (
            .O(N__5022),
            .I(N__5018));
    InMux I__983 (
            .O(N__5021),
            .I(N__5015));
    LocalMux I__982 (
            .O(N__5018),
            .I(n11_adj_399));
    LocalMux I__981 (
            .O(N__5015),
            .I(n11_adj_399));
    InMux I__980 (
            .O(N__5010),
            .I(N__5007));
    LocalMux I__979 (
            .O(N__5007),
            .I(n2566));
    InMux I__978 (
            .O(N__5004),
            .I(N__5001));
    LocalMux I__977 (
            .O(N__5001),
            .I(\eeprom.i2c.n39 ));
    CEMux I__976 (
            .O(N__4998),
            .I(N__4995));
    LocalMux I__975 (
            .O(N__4995),
            .I(N__4992));
    Span4Mux_v I__974 (
            .O(N__4992),
            .I(N__4989));
    Odrv4 I__973 (
            .O(N__4989),
            .I(\eeprom.i2c.n2406 ));
    InMux I__972 (
            .O(N__4986),
            .I(N__4982));
    InMux I__971 (
            .O(N__4985),
            .I(N__4979));
    LocalMux I__970 (
            .O(N__4982),
            .I(N__4976));
    LocalMux I__969 (
            .O(N__4979),
            .I(\eeprom.i2c.n37 ));
    Odrv4 I__968 (
            .O(N__4976),
            .I(\eeprom.i2c.n37 ));
    CascadeMux I__967 (
            .O(N__4971),
            .I(\eeprom.i2c.n1051_cascade_ ));
    CascadeMux I__966 (
            .O(N__4968),
            .I(N__4965));
    InMux I__965 (
            .O(N__4965),
            .I(N__4962));
    LocalMux I__964 (
            .O(N__4962),
            .I(\eeprom.i2c.n13 ));
    InMux I__963 (
            .O(N__4959),
            .I(N__4954));
    InMux I__962 (
            .O(N__4958),
            .I(N__4951));
    InMux I__961 (
            .O(N__4957),
            .I(N__4948));
    LocalMux I__960 (
            .O(N__4954),
            .I(sda_out));
    LocalMux I__959 (
            .O(N__4951),
            .I(sda_out));
    LocalMux I__958 (
            .O(N__4948),
            .I(sda_out));
    IoInMux I__957 (
            .O(N__4941),
            .I(N__4938));
    LocalMux I__956 (
            .O(N__4938),
            .I(N__4935));
    Span4Mux_s1_h I__955 (
            .O(N__4935),
            .I(N__4932));
    Sp12to4 I__954 (
            .O(N__4932),
            .I(N__4929));
    Span12Mux_v I__953 (
            .O(N__4929),
            .I(N__4925));
    InMux I__952 (
            .O(N__4928),
            .I(N__4920));
    Span12Mux_h I__951 (
            .O(N__4925),
            .I(N__4917));
    InMux I__950 (
            .O(N__4924),
            .I(N__4914));
    InMux I__949 (
            .O(N__4923),
            .I(N__4911));
    LocalMux I__948 (
            .O(N__4920),
            .I(N__4908));
    Odrv12 I__947 (
            .O(N__4917),
            .I(sda_enable));
    LocalMux I__946 (
            .O(N__4914),
            .I(sda_enable));
    LocalMux I__945 (
            .O(N__4911),
            .I(sda_enable));
    Odrv4 I__944 (
            .O(N__4908),
            .I(sda_enable));
    CascadeMux I__943 (
            .O(N__4899),
            .I(state_7_N_285_3_cascade_));
    InMux I__942 (
            .O(N__4896),
            .I(N__4893));
    LocalMux I__941 (
            .O(N__4893),
            .I(\eeprom.i2c.n2475 ));
    CascadeMux I__940 (
            .O(N__4890),
            .I(\eeprom.i2c.n2475_cascade_ ));
    CascadeMux I__939 (
            .O(N__4887),
            .I(n949_cascade_));
    InMux I__938 (
            .O(N__4884),
            .I(N__4880));
    InMux I__937 (
            .O(N__4883),
            .I(N__4877));
    LocalMux I__936 (
            .O(N__4880),
            .I(n949));
    LocalMux I__935 (
            .O(N__4877),
            .I(n949));
    CascadeMux I__934 (
            .O(N__4872),
            .I(n2547_cascade_));
    CascadeMux I__933 (
            .O(N__4869),
            .I(\eeprom.i2c.n2574_cascade_ ));
    InMux I__932 (
            .O(N__4866),
            .I(N__4863));
    LocalMux I__931 (
            .O(N__4863),
            .I(\eeprom.i2c.n2557 ));
    CascadeMux I__930 (
            .O(N__4860),
            .I(N__4857));
    InMux I__929 (
            .O(N__4857),
            .I(N__4853));
    SRMux I__928 (
            .O(N__4856),
            .I(N__4850));
    LocalMux I__927 (
            .O(N__4853),
            .I(N__4846));
    LocalMux I__926 (
            .O(N__4850),
            .I(N__4843));
    InMux I__925 (
            .O(N__4849),
            .I(N__4840));
    Span4Mux_v I__924 (
            .O(N__4846),
            .I(N__4837));
    Span4Mux_h I__923 (
            .O(N__4843),
            .I(N__4834));
    LocalMux I__922 (
            .O(N__4840),
            .I(N__4831));
    Odrv4 I__921 (
            .O(N__4837),
            .I(\eeprom.enable ));
    Odrv4 I__920 (
            .O(N__4834),
            .I(\eeprom.enable ));
    Odrv4 I__919 (
            .O(N__4831),
            .I(\eeprom.enable ));
    CascadeMux I__918 (
            .O(N__4824),
            .I(n2538_cascade_));
    CascadeMux I__917 (
            .O(N__4821),
            .I(n4_adj_411_cascade_));
    InMux I__916 (
            .O(N__4818),
            .I(N__4815));
    LocalMux I__915 (
            .O(N__4815),
            .I(n1835));
    CascadeMux I__914 (
            .O(N__4812),
            .I(n2507_cascade_));
    InMux I__913 (
            .O(N__4809),
            .I(N__4806));
    LocalMux I__912 (
            .O(N__4806),
            .I(n10_adj_394));
    CascadeMux I__911 (
            .O(N__4803),
            .I(N__4800));
    InMux I__910 (
            .O(N__4800),
            .I(N__4795));
    InMux I__909 (
            .O(N__4799),
            .I(N__4792));
    InMux I__908 (
            .O(N__4798),
            .I(N__4789));
    LocalMux I__907 (
            .O(N__4795),
            .I(\eeprom.i2c.n11_adj_379 ));
    LocalMux I__906 (
            .O(N__4792),
            .I(\eeprom.i2c.n11_adj_379 ));
    LocalMux I__905 (
            .O(N__4789),
            .I(\eeprom.i2c.n11_adj_379 ));
    CascadeMux I__904 (
            .O(N__4782),
            .I(\eeprom.i2c.n6_cascade_ ));
    CascadeMux I__903 (
            .O(N__4779),
            .I(\eeprom.i2c.counter2_7__N_256_cascade_ ));
    CEMux I__902 (
            .O(N__4776),
            .I(N__4773));
    LocalMux I__901 (
            .O(N__4773),
            .I(\eeprom.i2c.n1580 ));
    CascadeMux I__900 (
            .O(N__4770),
            .I(N__4767));
    InMux I__899 (
            .O(N__4767),
            .I(N__4764));
    LocalMux I__898 (
            .O(N__4764),
            .I(N__4760));
    InMux I__897 (
            .O(N__4763),
            .I(N__4757));
    Odrv4 I__896 (
            .O(N__4760),
            .I(rw));
    LocalMux I__895 (
            .O(N__4757),
            .I(rw));
    CascadeMux I__894 (
            .O(N__4752),
            .I(n1835_cascade_));
    InMux I__893 (
            .O(N__4749),
            .I(N__4746));
    LocalMux I__892 (
            .O(N__4746),
            .I(n2569));
    CascadeMux I__891 (
            .O(N__4743),
            .I(n11_adj_399_cascade_));
    SRMux I__890 (
            .O(N__4740),
            .I(N__4737));
    LocalMux I__889 (
            .O(N__4737),
            .I(\eeprom.i2c.n1669 ));
    CascadeMux I__888 (
            .O(N__4734),
            .I(\eeprom.i2c.n37_cascade_ ));
    InMux I__887 (
            .O(N__4731),
            .I(N__4725));
    InMux I__886 (
            .O(N__4730),
            .I(N__4725));
    LocalMux I__885 (
            .O(N__4725),
            .I(\eeprom.i2c.n33 ));
    CascadeMux I__884 (
            .O(N__4722),
            .I(\eeprom.i2c.n39_cascade_ ));
    CEMux I__883 (
            .O(N__4719),
            .I(N__4716));
    LocalMux I__882 (
            .O(N__4716),
            .I(N__4713));
    Odrv4 I__881 (
            .O(N__4713),
            .I(\eeprom.i2c.n1027 ));
    InMux I__880 (
            .O(N__4710),
            .I(N__4707));
    LocalMux I__879 (
            .O(N__4707),
            .I(\eeprom.delay_counter_15_N_171_3 ));
    InMux I__878 (
            .O(N__4704),
            .I(N__4701));
    LocalMux I__877 (
            .O(N__4701),
            .I(N__4696));
    InMux I__876 (
            .O(N__4700),
            .I(N__4693));
    InMux I__875 (
            .O(N__4699),
            .I(N__4690));
    Span4Mux_v I__874 (
            .O(N__4696),
            .I(N__4687));
    LocalMux I__873 (
            .O(N__4693),
            .I(\eeprom.delay_counter_3 ));
    LocalMux I__872 (
            .O(N__4690),
            .I(\eeprom.delay_counter_3 ));
    Odrv4 I__871 (
            .O(N__4687),
            .I(\eeprom.delay_counter_3 ));
    InMux I__870 (
            .O(N__4680),
            .I(N__4677));
    LocalMux I__869 (
            .O(N__4677),
            .I(\eeprom.delay_counter_15_N_171_11 ));
    InMux I__868 (
            .O(N__4674),
            .I(N__4671));
    LocalMux I__867 (
            .O(N__4671),
            .I(\eeprom.delay_counter_15_N_171_9 ));
    CascadeMux I__866 (
            .O(N__4668),
            .I(N__4665));
    InMux I__865 (
            .O(N__4665),
            .I(N__4660));
    InMux I__864 (
            .O(N__4664),
            .I(N__4655));
    InMux I__863 (
            .O(N__4663),
            .I(N__4655));
    LocalMux I__862 (
            .O(N__4660),
            .I(\eeprom.delay_counter_11 ));
    LocalMux I__861 (
            .O(N__4655),
            .I(\eeprom.delay_counter_11 ));
    CascadeMux I__860 (
            .O(N__4650),
            .I(N__4646));
    InMux I__859 (
            .O(N__4649),
            .I(N__4643));
    InMux I__858 (
            .O(N__4646),
            .I(N__4639));
    LocalMux I__857 (
            .O(N__4643),
            .I(N__4636));
    InMux I__856 (
            .O(N__4642),
            .I(N__4633));
    LocalMux I__855 (
            .O(N__4639),
            .I(\eeprom.delay_counter_7 ));
    Odrv4 I__854 (
            .O(N__4636),
            .I(\eeprom.delay_counter_7 ));
    LocalMux I__853 (
            .O(N__4633),
            .I(\eeprom.delay_counter_7 ));
    CascadeMux I__852 (
            .O(N__4626),
            .I(\eeprom.n6_cascade_ ));
    CascadeMux I__851 (
            .O(N__4623),
            .I(N__4619));
    CascadeMux I__850 (
            .O(N__4622),
            .I(N__4616));
    InMux I__849 (
            .O(N__4619),
            .I(N__4613));
    InMux I__848 (
            .O(N__4616),
            .I(N__4610));
    LocalMux I__847 (
            .O(N__4613),
            .I(N__4604));
    LocalMux I__846 (
            .O(N__4610),
            .I(N__4604));
    InMux I__845 (
            .O(N__4609),
            .I(N__4601));
    Odrv4 I__844 (
            .O(N__4604),
            .I(\eeprom.delay_counter_9 ));
    LocalMux I__843 (
            .O(N__4601),
            .I(\eeprom.delay_counter_9 ));
    InMux I__842 (
            .O(N__4596),
            .I(N__4593));
    LocalMux I__841 (
            .O(N__4593),
            .I(\eeprom.n8 ));
    InMux I__840 (
            .O(N__4590),
            .I(N__4587));
    LocalMux I__839 (
            .O(N__4587),
            .I(\eeprom.delay_counter_15_N_171_15 ));
    InMux I__838 (
            .O(N__4584),
            .I(N__4579));
    InMux I__837 (
            .O(N__4583),
            .I(N__4574));
    InMux I__836 (
            .O(N__4582),
            .I(N__4574));
    LocalMux I__835 (
            .O(N__4579),
            .I(\eeprom.delay_counter_15 ));
    LocalMux I__834 (
            .O(N__4574),
            .I(\eeprom.delay_counter_15 ));
    InMux I__833 (
            .O(N__4569),
            .I(N__4566));
    LocalMux I__832 (
            .O(N__4566),
            .I(\eeprom.delay_counter_15_N_171_14 ));
    InMux I__831 (
            .O(N__4563),
            .I(N__4558));
    InMux I__830 (
            .O(N__4562),
            .I(N__4553));
    InMux I__829 (
            .O(N__4561),
            .I(N__4553));
    LocalMux I__828 (
            .O(N__4558),
            .I(\eeprom.delay_counter_14 ));
    LocalMux I__827 (
            .O(N__4553),
            .I(\eeprom.delay_counter_14 ));
    InMux I__826 (
            .O(N__4548),
            .I(N__4535));
    InMux I__825 (
            .O(N__4547),
            .I(N__4532));
    CascadeMux I__824 (
            .O(N__4546),
            .I(N__4525));
    CascadeMux I__823 (
            .O(N__4545),
            .I(N__4522));
    CascadeMux I__822 (
            .O(N__4544),
            .I(N__4519));
    InMux I__821 (
            .O(N__4543),
            .I(N__4507));
    InMux I__820 (
            .O(N__4542),
            .I(N__4507));
    InMux I__819 (
            .O(N__4541),
            .I(N__4507));
    InMux I__818 (
            .O(N__4540),
            .I(N__4507));
    InMux I__817 (
            .O(N__4539),
            .I(N__4504));
    InMux I__816 (
            .O(N__4538),
            .I(N__4501));
    LocalMux I__815 (
            .O(N__4535),
            .I(N__4496));
    LocalMux I__814 (
            .O(N__4532),
            .I(N__4496));
    InMux I__813 (
            .O(N__4531),
            .I(N__4491));
    InMux I__812 (
            .O(N__4530),
            .I(N__4491));
    InMux I__811 (
            .O(N__4529),
            .I(N__4486));
    InMux I__810 (
            .O(N__4528),
            .I(N__4486));
    InMux I__809 (
            .O(N__4525),
            .I(N__4475));
    InMux I__808 (
            .O(N__4522),
            .I(N__4475));
    InMux I__807 (
            .O(N__4519),
            .I(N__4475));
    InMux I__806 (
            .O(N__4518),
            .I(N__4475));
    InMux I__805 (
            .O(N__4517),
            .I(N__4475));
    InMux I__804 (
            .O(N__4516),
            .I(N__4464));
    LocalMux I__803 (
            .O(N__4507),
            .I(N__4461));
    LocalMux I__802 (
            .O(N__4504),
            .I(N__4458));
    LocalMux I__801 (
            .O(N__4501),
            .I(N__4451));
    Span4Mux_h I__800 (
            .O(N__4496),
            .I(N__4451));
    LocalMux I__799 (
            .O(N__4491),
            .I(N__4451));
    LocalMux I__798 (
            .O(N__4486),
            .I(N__4446));
    LocalMux I__797 (
            .O(N__4475),
            .I(N__4446));
    InMux I__796 (
            .O(N__4474),
            .I(N__4439));
    InMux I__795 (
            .O(N__4473),
            .I(N__4439));
    InMux I__794 (
            .O(N__4472),
            .I(N__4439));
    InMux I__793 (
            .O(N__4471),
            .I(N__4428));
    InMux I__792 (
            .O(N__4470),
            .I(N__4428));
    InMux I__791 (
            .O(N__4469),
            .I(N__4428));
    InMux I__790 (
            .O(N__4468),
            .I(N__4428));
    InMux I__789 (
            .O(N__4467),
            .I(N__4428));
    LocalMux I__788 (
            .O(N__4464),
            .I(state_0));
    Odrv4 I__787 (
            .O(N__4461),
            .I(state_0));
    Odrv4 I__786 (
            .O(N__4458),
            .I(state_0));
    Odrv4 I__785 (
            .O(N__4451),
            .I(state_0));
    Odrv4 I__784 (
            .O(N__4446),
            .I(state_0));
    LocalMux I__783 (
            .O(N__4439),
            .I(state_0));
    LocalMux I__782 (
            .O(N__4428),
            .I(state_0));
    CascadeMux I__781 (
            .O(N__4413),
            .I(N__4405));
    CascadeMux I__780 (
            .O(N__4412),
            .I(N__4401));
    CascadeMux I__779 (
            .O(N__4411),
            .I(N__4398));
    CascadeMux I__778 (
            .O(N__4410),
            .I(N__4395));
    CascadeMux I__777 (
            .O(N__4409),
            .I(N__4392));
    InMux I__776 (
            .O(N__4408),
            .I(N__4387));
    InMux I__775 (
            .O(N__4405),
            .I(N__4387));
    InMux I__774 (
            .O(N__4404),
            .I(N__4384));
    InMux I__773 (
            .O(N__4401),
            .I(N__4377));
    InMux I__772 (
            .O(N__4398),
            .I(N__4377));
    InMux I__771 (
            .O(N__4395),
            .I(N__4377));
    InMux I__770 (
            .O(N__4392),
            .I(N__4374));
    LocalMux I__769 (
            .O(N__4387),
            .I(N__4367));
    LocalMux I__768 (
            .O(N__4384),
            .I(N__4362));
    LocalMux I__767 (
            .O(N__4377),
            .I(N__4362));
    LocalMux I__766 (
            .O(N__4374),
            .I(N__4359));
    CascadeMux I__765 (
            .O(N__4373),
            .I(N__4353));
    CascadeMux I__764 (
            .O(N__4372),
            .I(N__4350));
    CascadeMux I__763 (
            .O(N__4371),
            .I(N__4346));
    CascadeMux I__762 (
            .O(N__4370),
            .I(N__4343));
    Span4Mux_v I__761 (
            .O(N__4367),
            .I(N__4339));
    Span4Mux_h I__760 (
            .O(N__4362),
            .I(N__4336));
    Span4Mux_h I__759 (
            .O(N__4359),
            .I(N__4333));
    InMux I__758 (
            .O(N__4358),
            .I(N__4322));
    InMux I__757 (
            .O(N__4357),
            .I(N__4322));
    InMux I__756 (
            .O(N__4356),
            .I(N__4322));
    InMux I__755 (
            .O(N__4353),
            .I(N__4322));
    InMux I__754 (
            .O(N__4350),
            .I(N__4322));
    InMux I__753 (
            .O(N__4349),
            .I(N__4319));
    InMux I__752 (
            .O(N__4346),
            .I(N__4312));
    InMux I__751 (
            .O(N__4343),
            .I(N__4312));
    InMux I__750 (
            .O(N__4342),
            .I(N__4312));
    Odrv4 I__749 (
            .O(N__4339),
            .I(\eeprom.n1601 ));
    Odrv4 I__748 (
            .O(N__4336),
            .I(\eeprom.n1601 ));
    Odrv4 I__747 (
            .O(N__4333),
            .I(\eeprom.n1601 ));
    LocalMux I__746 (
            .O(N__4322),
            .I(\eeprom.n1601 ));
    LocalMux I__745 (
            .O(N__4319),
            .I(\eeprom.n1601 ));
    LocalMux I__744 (
            .O(N__4312),
            .I(\eeprom.n1601 ));
    InMux I__743 (
            .O(N__4299),
            .I(N__4296));
    LocalMux I__742 (
            .O(N__4296),
            .I(\eeprom.delay_counter_15_N_171_13 ));
    CascadeMux I__741 (
            .O(N__4293),
            .I(N__4289));
    InMux I__740 (
            .O(N__4292),
            .I(N__4285));
    InMux I__739 (
            .O(N__4289),
            .I(N__4282));
    InMux I__738 (
            .O(N__4288),
            .I(N__4279));
    LocalMux I__737 (
            .O(N__4285),
            .I(\eeprom.delay_counter_13 ));
    LocalMux I__736 (
            .O(N__4282),
            .I(\eeprom.delay_counter_13 ));
    LocalMux I__735 (
            .O(N__4279),
            .I(\eeprom.delay_counter_13 ));
    InMux I__734 (
            .O(N__4272),
            .I(N__4268));
    InMux I__733 (
            .O(N__4271),
            .I(N__4265));
    LocalMux I__732 (
            .O(N__4268),
            .I(N__4262));
    LocalMux I__731 (
            .O(N__4265),
            .I(delay_counter_5));
    Odrv4 I__730 (
            .O(N__4262),
            .I(delay_counter_5));
    InMux I__729 (
            .O(N__4257),
            .I(N__4254));
    LocalMux I__728 (
            .O(N__4254),
            .I(n16_adj_407));
    CascadeMux I__727 (
            .O(N__4251),
            .I(N__4248));
    InMux I__726 (
            .O(N__4248),
            .I(N__4244));
    InMux I__725 (
            .O(N__4247),
            .I(N__4241));
    LocalMux I__724 (
            .O(N__4244),
            .I(N__4238));
    LocalMux I__723 (
            .O(N__4241),
            .I(delay_counter_2));
    Odrv4 I__722 (
            .O(N__4238),
            .I(delay_counter_2));
    InMux I__721 (
            .O(N__4233),
            .I(N__4230));
    LocalMux I__720 (
            .O(N__4230),
            .I(n17_adj_406));
    InMux I__719 (
            .O(N__4227),
            .I(N__4224));
    LocalMux I__718 (
            .O(N__4224),
            .I(n2536));
    InMux I__717 (
            .O(N__4221),
            .I(N__4215));
    InMux I__716 (
            .O(N__4220),
            .I(N__4210));
    InMux I__715 (
            .O(N__4219),
            .I(N__4210));
    InMux I__714 (
            .O(N__4218),
            .I(N__4207));
    LocalMux I__713 (
            .O(N__4215),
            .I(N__4204));
    LocalMux I__712 (
            .O(N__4210),
            .I(N__4201));
    LocalMux I__711 (
            .O(N__4207),
            .I(N__4198));
    Span4Mux_v I__710 (
            .O(N__4204),
            .I(N__4193));
    Span4Mux_h I__709 (
            .O(N__4201),
            .I(N__4193));
    Odrv4 I__708 (
            .O(N__4198),
            .I(read_N));
    Odrv4 I__707 (
            .O(N__4193),
            .I(read_N));
    InMux I__706 (
            .O(N__4188),
            .I(N__4184));
    InMux I__705 (
            .O(N__4187),
            .I(N__4181));
    LocalMux I__704 (
            .O(N__4184),
            .I(delay_counter_22));
    LocalMux I__703 (
            .O(N__4181),
            .I(delay_counter_22));
    InMux I__702 (
            .O(N__4176),
            .I(N__4172));
    InMux I__701 (
            .O(N__4175),
            .I(N__4169));
    LocalMux I__700 (
            .O(N__4172),
            .I(delay_counter_25));
    LocalMux I__699 (
            .O(N__4169),
            .I(delay_counter_25));
    CascadeMux I__698 (
            .O(N__4164),
            .I(N__4160));
    InMux I__697 (
            .O(N__4163),
            .I(N__4157));
    InMux I__696 (
            .O(N__4160),
            .I(N__4154));
    LocalMux I__695 (
            .O(N__4157),
            .I(delay_counter_20));
    LocalMux I__694 (
            .O(N__4154),
            .I(delay_counter_20));
    InMux I__693 (
            .O(N__4149),
            .I(N__4146));
    LocalMux I__692 (
            .O(N__4146),
            .I(n8_adj_412));
    InMux I__691 (
            .O(N__4143),
            .I(N__4140));
    LocalMux I__690 (
            .O(N__4140),
            .I(n9_adj_404));
    InMux I__689 (
            .O(N__4137),
            .I(N__4130));
    InMux I__688 (
            .O(N__4136),
            .I(N__4130));
    InMux I__687 (
            .O(N__4135),
            .I(N__4127));
    LocalMux I__686 (
            .O(N__4130),
            .I(N__4124));
    LocalMux I__685 (
            .O(N__4127),
            .I(delay_counter_31));
    Odrv4 I__684 (
            .O(N__4124),
            .I(delay_counter_31));
    CascadeMux I__683 (
            .O(N__4119),
            .I(n9_adj_404_cascade_));
    SRMux I__682 (
            .O(N__4116),
            .I(N__4113));
    LocalMux I__681 (
            .O(N__4113),
            .I(N__4108));
    SRMux I__680 (
            .O(N__4112),
            .I(N__4105));
    SRMux I__679 (
            .O(N__4111),
            .I(N__4102));
    Span4Mux_v I__678 (
            .O(N__4108),
            .I(N__4096));
    LocalMux I__677 (
            .O(N__4105),
            .I(N__4096));
    LocalMux I__676 (
            .O(N__4102),
            .I(N__4093));
    SRMux I__675 (
            .O(N__4101),
            .I(N__4090));
    Span4Mux_h I__674 (
            .O(N__4096),
            .I(N__4087));
    Span4Mux_h I__673 (
            .O(N__4093),
            .I(N__4084));
    LocalMux I__672 (
            .O(N__4090),
            .I(N__4081));
    Odrv4 I__671 (
            .O(N__4087),
            .I(addr_10__N_70));
    Odrv4 I__670 (
            .O(N__4084),
            .I(addr_10__N_70));
    Odrv12 I__669 (
            .O(N__4081),
            .I(addr_10__N_70));
    InMux I__668 (
            .O(N__4074),
            .I(N__4070));
    InMux I__667 (
            .O(N__4073),
            .I(N__4067));
    LocalMux I__666 (
            .O(N__4070),
            .I(delay_counter_29));
    LocalMux I__665 (
            .O(N__4067),
            .I(delay_counter_29));
    InMux I__664 (
            .O(N__4062),
            .I(N__4058));
    InMux I__663 (
            .O(N__4061),
            .I(N__4055));
    LocalMux I__662 (
            .O(N__4058),
            .I(delay_counter_28));
    LocalMux I__661 (
            .O(N__4055),
            .I(delay_counter_28));
    InMux I__660 (
            .O(N__4050),
            .I(N__4044));
    InMux I__659 (
            .O(N__4049),
            .I(N__4044));
    LocalMux I__658 (
            .O(N__4044),
            .I(N__4041));
    Odrv4 I__657 (
            .O(N__4041),
            .I(n10_adj_403));
    InMux I__656 (
            .O(N__4038),
            .I(N__4034));
    InMux I__655 (
            .O(N__4037),
            .I(N__4031));
    LocalMux I__654 (
            .O(N__4034),
            .I(delay_counter_26));
    LocalMux I__653 (
            .O(N__4031),
            .I(delay_counter_26));
    InMux I__652 (
            .O(N__4026),
            .I(N__4022));
    InMux I__651 (
            .O(N__4025),
            .I(N__4019));
    LocalMux I__650 (
            .O(N__4022),
            .I(delay_counter_30));
    LocalMux I__649 (
            .O(N__4019),
            .I(delay_counter_30));
    CascadeMux I__648 (
            .O(N__4014),
            .I(N__4010));
    InMux I__647 (
            .O(N__4013),
            .I(N__4007));
    InMux I__646 (
            .O(N__4010),
            .I(N__4004));
    LocalMux I__645 (
            .O(N__4007),
            .I(delay_counter_27));
    LocalMux I__644 (
            .O(N__4004),
            .I(delay_counter_27));
    InMux I__643 (
            .O(N__3999),
            .I(N__3995));
    InMux I__642 (
            .O(N__3998),
            .I(N__3992));
    LocalMux I__641 (
            .O(N__3995),
            .I(delay_counter_24));
    LocalMux I__640 (
            .O(N__3992),
            .I(delay_counter_24));
    CascadeMux I__639 (
            .O(N__3987),
            .I(N__3984));
    InMux I__638 (
            .O(N__3984),
            .I(N__3980));
    InMux I__637 (
            .O(N__3983),
            .I(N__3977));
    LocalMux I__636 (
            .O(N__3980),
            .I(N__3974));
    LocalMux I__635 (
            .O(N__3977),
            .I(N__3971));
    Odrv4 I__634 (
            .O(N__3974),
            .I(n14_adj_401));
    Odrv4 I__633 (
            .O(N__3971),
            .I(n14_adj_401));
    InMux I__632 (
            .O(N__3966),
            .I(N__3963));
    LocalMux I__631 (
            .O(N__3963),
            .I(\eeprom.delay_counter_15_N_171_7 ));
    SRMux I__630 (
            .O(N__3960),
            .I(N__3957));
    LocalMux I__629 (
            .O(N__3957),
            .I(N__3954));
    Span4Mux_h I__628 (
            .O(N__3954),
            .I(N__3944));
    InMux I__627 (
            .O(N__3953),
            .I(N__3941));
    InMux I__626 (
            .O(N__3952),
            .I(N__3936));
    InMux I__625 (
            .O(N__3951),
            .I(N__3936));
    InMux I__624 (
            .O(N__3950),
            .I(N__3927));
    InMux I__623 (
            .O(N__3949),
            .I(N__3927));
    InMux I__622 (
            .O(N__3948),
            .I(N__3927));
    InMux I__621 (
            .O(N__3947),
            .I(N__3927));
    Odrv4 I__620 (
            .O(N__3944),
            .I(state_1));
    LocalMux I__619 (
            .O(N__3941),
            .I(state_1));
    LocalMux I__618 (
            .O(N__3936),
            .I(state_1));
    LocalMux I__617 (
            .O(N__3927),
            .I(state_1));
    CEMux I__616 (
            .O(N__3918),
            .I(N__3915));
    LocalMux I__615 (
            .O(N__3915),
            .I(N__3912));
    Odrv12 I__614 (
            .O(N__3912),
            .I(n1568));
    InMux I__613 (
            .O(N__3909),
            .I(N__3905));
    InMux I__612 (
            .O(N__3908),
            .I(N__3902));
    LocalMux I__611 (
            .O(N__3905),
            .I(delay_counter_7));
    LocalMux I__610 (
            .O(N__3902),
            .I(delay_counter_7));
    InMux I__609 (
            .O(N__3897),
            .I(N__3893));
    InMux I__608 (
            .O(N__3896),
            .I(N__3890));
    LocalMux I__607 (
            .O(N__3893),
            .I(delay_counter_8));
    LocalMux I__606 (
            .O(N__3890),
            .I(delay_counter_8));
    CascadeMux I__605 (
            .O(N__3885),
            .I(N__3881));
    InMux I__604 (
            .O(N__3884),
            .I(N__3878));
    InMux I__603 (
            .O(N__3881),
            .I(N__3875));
    LocalMux I__602 (
            .O(N__3878),
            .I(delay_counter_1));
    LocalMux I__601 (
            .O(N__3875),
            .I(delay_counter_1));
    InMux I__600 (
            .O(N__3870),
            .I(N__3866));
    InMux I__599 (
            .O(N__3869),
            .I(N__3863));
    LocalMux I__598 (
            .O(N__3866),
            .I(delay_counter_4));
    LocalMux I__597 (
            .O(N__3863),
            .I(delay_counter_4));
    InMux I__596 (
            .O(N__3858),
            .I(N__3854));
    InMux I__595 (
            .O(N__3857),
            .I(N__3851));
    LocalMux I__594 (
            .O(N__3854),
            .I(delay_counter_10));
    LocalMux I__593 (
            .O(N__3851),
            .I(delay_counter_10));
    InMux I__592 (
            .O(N__3846),
            .I(N__3842));
    InMux I__591 (
            .O(N__3845),
            .I(N__3839));
    LocalMux I__590 (
            .O(N__3842),
            .I(delay_counter_12));
    LocalMux I__589 (
            .O(N__3839),
            .I(delay_counter_12));
    CascadeMux I__588 (
            .O(N__3834),
            .I(N__3830));
    InMux I__587 (
            .O(N__3833),
            .I(N__3827));
    InMux I__586 (
            .O(N__3830),
            .I(N__3824));
    LocalMux I__585 (
            .O(N__3827),
            .I(delay_counter_11));
    LocalMux I__584 (
            .O(N__3824),
            .I(delay_counter_11));
    InMux I__583 (
            .O(N__3819),
            .I(N__3815));
    InMux I__582 (
            .O(N__3818),
            .I(N__3812));
    LocalMux I__581 (
            .O(N__3815),
            .I(delay_counter_13));
    LocalMux I__580 (
            .O(N__3812),
            .I(delay_counter_13));
    CascadeMux I__579 (
            .O(N__3807),
            .I(n2512_cascade_));
    InMux I__578 (
            .O(N__3804),
            .I(N__3800));
    InMux I__577 (
            .O(N__3803),
            .I(N__3797));
    LocalMux I__576 (
            .O(N__3800),
            .I(delay_counter_16));
    LocalMux I__575 (
            .O(N__3797),
            .I(delay_counter_16));
    InMux I__574 (
            .O(N__3792),
            .I(N__3788));
    InMux I__573 (
            .O(N__3791),
            .I(N__3785));
    LocalMux I__572 (
            .O(N__3788),
            .I(delay_counter_18));
    LocalMux I__571 (
            .O(N__3785),
            .I(delay_counter_18));
    CascadeMux I__570 (
            .O(N__3780),
            .I(n2495_cascade_));
    InMux I__569 (
            .O(N__3777),
            .I(N__3773));
    InMux I__568 (
            .O(N__3776),
            .I(N__3770));
    LocalMux I__567 (
            .O(N__3773),
            .I(delay_counter_19));
    LocalMux I__566 (
            .O(N__3770),
            .I(delay_counter_19));
    InMux I__565 (
            .O(N__3765),
            .I(N__3761));
    InMux I__564 (
            .O(N__3764),
            .I(N__3758));
    LocalMux I__563 (
            .O(N__3761),
            .I(delay_counter_9));
    LocalMux I__562 (
            .O(N__3758),
            .I(delay_counter_9));
    InMux I__561 (
            .O(N__3753),
            .I(N__3749));
    InMux I__560 (
            .O(N__3752),
            .I(N__3746));
    LocalMux I__559 (
            .O(N__3749),
            .I(delay_counter_6));
    LocalMux I__558 (
            .O(N__3746),
            .I(delay_counter_6));
    CascadeMux I__557 (
            .O(N__3741),
            .I(N__3737));
    InMux I__556 (
            .O(N__3740),
            .I(N__3734));
    InMux I__555 (
            .O(N__3737),
            .I(N__3731));
    LocalMux I__554 (
            .O(N__3734),
            .I(delay_counter_3));
    LocalMux I__553 (
            .O(N__3731),
            .I(delay_counter_3));
    InMux I__552 (
            .O(N__3726),
            .I(N__3722));
    InMux I__551 (
            .O(N__3725),
            .I(N__3719));
    LocalMux I__550 (
            .O(N__3722),
            .I(delay_counter_0));
    LocalMux I__549 (
            .O(N__3719),
            .I(delay_counter_0));
    InMux I__548 (
            .O(N__3714),
            .I(N__3710));
    InMux I__547 (
            .O(N__3713),
            .I(N__3707));
    LocalMux I__546 (
            .O(N__3710),
            .I(delay_counter_17));
    LocalMux I__545 (
            .O(N__3707),
            .I(delay_counter_17));
    InMux I__544 (
            .O(N__3702),
            .I(N__3698));
    InMux I__543 (
            .O(N__3701),
            .I(N__3695));
    LocalMux I__542 (
            .O(N__3698),
            .I(delay_counter_15));
    LocalMux I__541 (
            .O(N__3695),
            .I(delay_counter_15));
    InMux I__540 (
            .O(N__3690),
            .I(N__3686));
    InMux I__539 (
            .O(N__3689),
            .I(N__3683));
    LocalMux I__538 (
            .O(N__3686),
            .I(delay_counter_14));
    LocalMux I__537 (
            .O(N__3683),
            .I(delay_counter_14));
    InMux I__536 (
            .O(N__3678),
            .I(N__3675));
    LocalMux I__535 (
            .O(N__3675),
            .I(n8));
    InMux I__534 (
            .O(N__3672),
            .I(N__3668));
    InMux I__533 (
            .O(N__3671),
            .I(N__3665));
    LocalMux I__532 (
            .O(N__3668),
            .I(delay_counter_21));
    LocalMux I__531 (
            .O(N__3665),
            .I(delay_counter_21));
    InMux I__530 (
            .O(N__3660),
            .I(N__3656));
    InMux I__529 (
            .O(N__3659),
            .I(N__3653));
    LocalMux I__528 (
            .O(N__3656),
            .I(delay_counter_23));
    LocalMux I__527 (
            .O(N__3653),
            .I(delay_counter_23));
    InMux I__526 (
            .O(N__3648),
            .I(N__3645));
    LocalMux I__525 (
            .O(N__3645),
            .I(n6_adj_413));
    InMux I__524 (
            .O(N__3642),
            .I(N__3639));
    LocalMux I__523 (
            .O(N__3639),
            .I(N__3636));
    Odrv4 I__522 (
            .O(N__3636),
            .I(\eeprom.delay_counter_15_N_171_4 ));
    CascadeMux I__521 (
            .O(N__3633),
            .I(N__3630));
    InMux I__520 (
            .O(N__3630),
            .I(N__3627));
    LocalMux I__519 (
            .O(N__3627),
            .I(N__3622));
    InMux I__518 (
            .O(N__3626),
            .I(N__3617));
    InMux I__517 (
            .O(N__3625),
            .I(N__3617));
    Odrv4 I__516 (
            .O(N__3622),
            .I(\eeprom.delay_counter_4 ));
    LocalMux I__515 (
            .O(N__3617),
            .I(\eeprom.delay_counter_4 ));
    InMux I__514 (
            .O(N__3612),
            .I(N__3609));
    LocalMux I__513 (
            .O(N__3609),
            .I(n324));
    InMux I__512 (
            .O(N__3606),
            .I(N__3600));
    InMux I__511 (
            .O(N__3605),
            .I(N__3597));
    InMux I__510 (
            .O(N__3604),
            .I(N__3592));
    InMux I__509 (
            .O(N__3603),
            .I(N__3592));
    LocalMux I__508 (
            .O(N__3600),
            .I(\eeprom.n1500 ));
    LocalMux I__507 (
            .O(N__3597),
            .I(\eeprom.n1500 ));
    LocalMux I__506 (
            .O(N__3592),
            .I(\eeprom.n1500 ));
    CascadeMux I__505 (
            .O(N__3585),
            .I(n6_adj_405_cascade_));
    InMux I__504 (
            .O(N__3582),
            .I(N__3579));
    LocalMux I__503 (
            .O(N__3579),
            .I(n41));
    InMux I__502 (
            .O(N__3576),
            .I(N__3573));
    LocalMux I__501 (
            .O(N__3573),
            .I(\eeprom.n1018 ));
    CascadeMux I__500 (
            .O(N__3570),
            .I(n2483_cascade_));
    InMux I__499 (
            .O(N__3567),
            .I(N__3564));
    LocalMux I__498 (
            .O(N__3564),
            .I(\eeprom.n2453 ));
    CascadeMux I__497 (
            .O(N__3561),
            .I(n1568_cascade_));
    InMux I__496 (
            .O(N__3558),
            .I(\eeprom.n2254 ));
    CascadeMux I__495 (
            .O(N__3555),
            .I(N__3544));
    CascadeMux I__494 (
            .O(N__3554),
            .I(N__3540));
    CascadeMux I__493 (
            .O(N__3553),
            .I(N__3536));
    CascadeMux I__492 (
            .O(N__3552),
            .I(N__3532));
    CascadeMux I__491 (
            .O(N__3551),
            .I(N__3529));
    CascadeMux I__490 (
            .O(N__3550),
            .I(N__3525));
    CascadeMux I__489 (
            .O(N__3549),
            .I(N__3521));
    CascadeMux I__488 (
            .O(N__3548),
            .I(N__3517));
    InMux I__487 (
            .O(N__3547),
            .I(N__3499));
    InMux I__486 (
            .O(N__3544),
            .I(N__3499));
    InMux I__485 (
            .O(N__3543),
            .I(N__3499));
    InMux I__484 (
            .O(N__3540),
            .I(N__3499));
    InMux I__483 (
            .O(N__3539),
            .I(N__3499));
    InMux I__482 (
            .O(N__3536),
            .I(N__3499));
    InMux I__481 (
            .O(N__3535),
            .I(N__3499));
    InMux I__480 (
            .O(N__3532),
            .I(N__3499));
    InMux I__479 (
            .O(N__3529),
            .I(N__3482));
    InMux I__478 (
            .O(N__3528),
            .I(N__3482));
    InMux I__477 (
            .O(N__3525),
            .I(N__3482));
    InMux I__476 (
            .O(N__3524),
            .I(N__3482));
    InMux I__475 (
            .O(N__3521),
            .I(N__3482));
    InMux I__474 (
            .O(N__3520),
            .I(N__3482));
    InMux I__473 (
            .O(N__3517),
            .I(N__3482));
    InMux I__472 (
            .O(N__3516),
            .I(N__3482));
    LocalMux I__471 (
            .O(N__3499),
            .I(\eeprom.n642 ));
    LocalMux I__470 (
            .O(N__3482),
            .I(\eeprom.n642 ));
    InMux I__469 (
            .O(N__3477),
            .I(\eeprom.n2255 ));
    InMux I__468 (
            .O(N__3474),
            .I(N__3471));
    LocalMux I__467 (
            .O(N__3471),
            .I(\eeprom.n14 ));
    CascadeMux I__466 (
            .O(N__3468),
            .I(\eeprom.n13_cascade_ ));
    CascadeMux I__465 (
            .O(N__3465),
            .I(\eeprom.n7_cascade_ ));
    InMux I__464 (
            .O(N__3462),
            .I(N__3459));
    LocalMux I__463 (
            .O(N__3459),
            .I(N__3456));
    Odrv4 I__462 (
            .O(N__3456),
            .I(\eeprom.delay_counter_15_N_171_1 ));
    InMux I__461 (
            .O(N__3453),
            .I(N__3450));
    LocalMux I__460 (
            .O(N__3450),
            .I(N__3445));
    InMux I__459 (
            .O(N__3449),
            .I(N__3440));
    InMux I__458 (
            .O(N__3448),
            .I(N__3440));
    Odrv4 I__457 (
            .O(N__3445),
            .I(\eeprom.delay_counter_1 ));
    LocalMux I__456 (
            .O(N__3440),
            .I(\eeprom.delay_counter_1 ));
    InMux I__455 (
            .O(N__3435),
            .I(N__3432));
    LocalMux I__454 (
            .O(N__3432),
            .I(N__3429));
    Odrv4 I__453 (
            .O(N__3429),
            .I(\eeprom.delay_counter_15_N_171_0 ));
    CascadeMux I__452 (
            .O(N__3426),
            .I(N__3423));
    InMux I__451 (
            .O(N__3423),
            .I(N__3420));
    LocalMux I__450 (
            .O(N__3420),
            .I(N__3415));
    InMux I__449 (
            .O(N__3419),
            .I(N__3410));
    InMux I__448 (
            .O(N__3418),
            .I(N__3410));
    Odrv4 I__447 (
            .O(N__3415),
            .I(\eeprom.delay_counter_0 ));
    LocalMux I__446 (
            .O(N__3410),
            .I(\eeprom.delay_counter_0 ));
    InMux I__445 (
            .O(N__3405),
            .I(N__3402));
    LocalMux I__444 (
            .O(N__3402),
            .I(N__3399));
    Odrv4 I__443 (
            .O(N__3399),
            .I(\eeprom.delay_counter_15_N_171_5 ));
    InMux I__442 (
            .O(N__3396),
            .I(N__3393));
    LocalMux I__441 (
            .O(N__3393),
            .I(N__3388));
    InMux I__440 (
            .O(N__3392),
            .I(N__3383));
    InMux I__439 (
            .O(N__3391),
            .I(N__3383));
    Odrv4 I__438 (
            .O(N__3388),
            .I(\eeprom.delay_counter_5 ));
    LocalMux I__437 (
            .O(N__3383),
            .I(\eeprom.delay_counter_5 ));
    InMux I__436 (
            .O(N__3378),
            .I(N__3375));
    LocalMux I__435 (
            .O(N__3375),
            .I(\eeprom.delay_counter_15_N_171_10 ));
    CascadeMux I__434 (
            .O(N__3372),
            .I(N__3367));
    InMux I__433 (
            .O(N__3371),
            .I(N__3364));
    InMux I__432 (
            .O(N__3370),
            .I(N__3359));
    InMux I__431 (
            .O(N__3367),
            .I(N__3359));
    LocalMux I__430 (
            .O(N__3364),
            .I(\eeprom.delay_counter_10 ));
    LocalMux I__429 (
            .O(N__3359),
            .I(\eeprom.delay_counter_10 ));
    InMux I__428 (
            .O(N__3354),
            .I(\eeprom.n2245 ));
    CascadeMux I__427 (
            .O(N__3351),
            .I(N__3348));
    InMux I__426 (
            .O(N__3348),
            .I(N__3344));
    CascadeMux I__425 (
            .O(N__3347),
            .I(N__3340));
    LocalMux I__424 (
            .O(N__3344),
            .I(N__3337));
    InMux I__423 (
            .O(N__3343),
            .I(N__3332));
    InMux I__422 (
            .O(N__3340),
            .I(N__3332));
    Odrv4 I__421 (
            .O(N__3337),
            .I(\eeprom.delay_counter_6 ));
    LocalMux I__420 (
            .O(N__3332),
            .I(\eeprom.delay_counter_6 ));
    InMux I__419 (
            .O(N__3327),
            .I(N__3324));
    LocalMux I__418 (
            .O(N__3324),
            .I(N__3321));
    Odrv4 I__417 (
            .O(N__3321),
            .I(\eeprom.delay_counter_15_N_171_6 ));
    InMux I__416 (
            .O(N__3318),
            .I(\eeprom.n2246 ));
    InMux I__415 (
            .O(N__3315),
            .I(\eeprom.n2247 ));
    InMux I__414 (
            .O(N__3312),
            .I(N__3307));
    InMux I__413 (
            .O(N__3311),
            .I(N__3302));
    InMux I__412 (
            .O(N__3310),
            .I(N__3302));
    LocalMux I__411 (
            .O(N__3307),
            .I(\eeprom.delay_counter_8 ));
    LocalMux I__410 (
            .O(N__3302),
            .I(\eeprom.delay_counter_8 ));
    InMux I__409 (
            .O(N__3297),
            .I(N__3294));
    LocalMux I__408 (
            .O(N__3294),
            .I(\eeprom.delay_counter_15_N_171_8 ));
    InMux I__407 (
            .O(N__3291),
            .I(bfn_18_18_0_));
    InMux I__406 (
            .O(N__3288),
            .I(\eeprom.n2249 ));
    InMux I__405 (
            .O(N__3285),
            .I(\eeprom.n2250 ));
    InMux I__404 (
            .O(N__3282),
            .I(\eeprom.n2251 ));
    InMux I__403 (
            .O(N__3279),
            .I(N__3274));
    InMux I__402 (
            .O(N__3278),
            .I(N__3269));
    InMux I__401 (
            .O(N__3277),
            .I(N__3269));
    LocalMux I__400 (
            .O(N__3274),
            .I(\eeprom.delay_counter_12 ));
    LocalMux I__399 (
            .O(N__3269),
            .I(\eeprom.delay_counter_12 ));
    CascadeMux I__398 (
            .O(N__3264),
            .I(N__3261));
    InMux I__397 (
            .O(N__3261),
            .I(N__3258));
    LocalMux I__396 (
            .O(N__3258),
            .I(\eeprom.delay_counter_15_N_171_12 ));
    InMux I__395 (
            .O(N__3255),
            .I(\eeprom.n2252 ));
    InMux I__394 (
            .O(N__3252),
            .I(\eeprom.n2253 ));
    InMux I__393 (
            .O(N__3249),
            .I(n2290));
    InMux I__392 (
            .O(N__3246),
            .I(n2291));
    InMux I__391 (
            .O(N__3243),
            .I(n2292));
    InMux I__390 (
            .O(N__3240),
            .I(n2293));
    InMux I__389 (
            .O(N__3237),
            .I(\eeprom.n2241 ));
    CascadeMux I__388 (
            .O(N__3234),
            .I(N__3231));
    InMux I__387 (
            .O(N__3231),
            .I(N__3228));
    LocalMux I__386 (
            .O(N__3228),
            .I(N__3223));
    InMux I__385 (
            .O(N__3227),
            .I(N__3218));
    InMux I__384 (
            .O(N__3226),
            .I(N__3218));
    Odrv4 I__383 (
            .O(N__3223),
            .I(\eeprom.delay_counter_2 ));
    LocalMux I__382 (
            .O(N__3218),
            .I(\eeprom.delay_counter_2 ));
    CascadeMux I__381 (
            .O(N__3213),
            .I(N__3210));
    InMux I__380 (
            .O(N__3210),
            .I(N__3207));
    LocalMux I__379 (
            .O(N__3207),
            .I(N__3204));
    Odrv4 I__378 (
            .O(N__3204),
            .I(\eeprom.delay_counter_15_N_171_2 ));
    InMux I__377 (
            .O(N__3201),
            .I(\eeprom.n2242 ));
    InMux I__376 (
            .O(N__3198),
            .I(\eeprom.n2243 ));
    InMux I__375 (
            .O(N__3195),
            .I(\eeprom.n2244 ));
    InMux I__374 (
            .O(N__3192),
            .I(n2281));
    InMux I__373 (
            .O(N__3189),
            .I(n2282));
    InMux I__372 (
            .O(N__3186),
            .I(n2283));
    InMux I__371 (
            .O(N__3183),
            .I(n2284));
    InMux I__370 (
            .O(N__3180),
            .I(n2285));
    InMux I__369 (
            .O(N__3177),
            .I(bfn_17_24_0_));
    InMux I__368 (
            .O(N__3174),
            .I(n2287));
    InMux I__367 (
            .O(N__3171),
            .I(n2288));
    InMux I__366 (
            .O(N__3168),
            .I(n2289));
    InMux I__365 (
            .O(N__3165),
            .I(n2272));
    InMux I__364 (
            .O(N__3162),
            .I(n2273));
    InMux I__363 (
            .O(N__3159),
            .I(n2274));
    InMux I__362 (
            .O(N__3156),
            .I(n2275));
    InMux I__361 (
            .O(N__3153),
            .I(n2276));
    InMux I__360 (
            .O(N__3150),
            .I(n2277));
    InMux I__359 (
            .O(N__3147),
            .I(bfn_17_23_0_));
    InMux I__358 (
            .O(N__3144),
            .I(n2279));
    InMux I__357 (
            .O(N__3141),
            .I(n2280));
    InMux I__356 (
            .O(N__3138),
            .I(n2263));
    InMux I__355 (
            .O(N__3135),
            .I(n2264));
    InMux I__354 (
            .O(N__3132),
            .I(n2265));
    InMux I__353 (
            .O(N__3129),
            .I(n2266));
    InMux I__352 (
            .O(N__3126),
            .I(n2267));
    InMux I__351 (
            .O(N__3123),
            .I(n2268));
    InMux I__350 (
            .O(N__3120),
            .I(n2269));
    InMux I__349 (
            .O(N__3117),
            .I(bfn_17_22_0_));
    InMux I__348 (
            .O(N__3114),
            .I(n2271));
    CascadeMux I__347 (
            .O(N__3111),
            .I(n693_cascade_));
    InMux I__346 (
            .O(N__3108),
            .I(bfn_17_21_0_));
    InMux I__345 (
            .O(N__3105),
            .I(N__3102));
    LocalMux I__344 (
            .O(N__3102),
            .I(n7));
    InMux I__343 (
            .O(N__3099),
            .I(n2312));
    InMux I__342 (
            .O(N__3096),
            .I(N__3093));
    LocalMux I__341 (
            .O(N__3093),
            .I(n6_adj_410));
    InMux I__340 (
            .O(N__3090),
            .I(n2313));
    InMux I__339 (
            .O(N__3087),
            .I(N__3080));
    InMux I__338 (
            .O(N__3086),
            .I(N__3080));
    InMux I__337 (
            .O(N__3085),
            .I(N__3077));
    LocalMux I__336 (
            .O(N__3080),
            .I(blink_counter_21));
    LocalMux I__335 (
            .O(N__3077),
            .I(blink_counter_21));
    InMux I__334 (
            .O(N__3072),
            .I(n2314));
    InMux I__333 (
            .O(N__3069),
            .I(N__3062));
    InMux I__332 (
            .O(N__3068),
            .I(N__3062));
    InMux I__331 (
            .O(N__3067),
            .I(N__3059));
    LocalMux I__330 (
            .O(N__3062),
            .I(blink_counter_22));
    LocalMux I__329 (
            .O(N__3059),
            .I(blink_counter_22));
    InMux I__328 (
            .O(N__3054),
            .I(n2315));
    CascadeMux I__327 (
            .O(N__3051),
            .I(N__3047));
    CascadeMux I__326 (
            .O(N__3050),
            .I(N__3044));
    InMux I__325 (
            .O(N__3047),
            .I(N__3038));
    InMux I__324 (
            .O(N__3044),
            .I(N__3038));
    InMux I__323 (
            .O(N__3043),
            .I(N__3035));
    LocalMux I__322 (
            .O(N__3038),
            .I(blink_counter_23));
    LocalMux I__321 (
            .O(N__3035),
            .I(blink_counter_23));
    InMux I__320 (
            .O(N__3030),
            .I(n2316));
    InMux I__319 (
            .O(N__3027),
            .I(N__3020));
    InMux I__318 (
            .O(N__3026),
            .I(N__3020));
    InMux I__317 (
            .O(N__3025),
            .I(N__3017));
    LocalMux I__316 (
            .O(N__3020),
            .I(blink_counter_24));
    LocalMux I__315 (
            .O(N__3017),
            .I(blink_counter_24));
    InMux I__314 (
            .O(N__3012),
            .I(bfn_14_24_0_));
    InMux I__313 (
            .O(N__3009),
            .I(n2318));
    InMux I__312 (
            .O(N__3006),
            .I(N__3002));
    InMux I__311 (
            .O(N__3005),
            .I(N__2999));
    LocalMux I__310 (
            .O(N__3002),
            .I(blink_counter_25));
    LocalMux I__309 (
            .O(N__2999),
            .I(blink_counter_25));
    InMux I__308 (
            .O(N__2994),
            .I(N__2991));
    LocalMux I__307 (
            .O(N__2991),
            .I(n16));
    InMux I__306 (
            .O(N__2988),
            .I(n2303));
    InMux I__305 (
            .O(N__2985),
            .I(N__2982));
    LocalMux I__304 (
            .O(N__2982),
            .I(n15));
    InMux I__303 (
            .O(N__2979),
            .I(n2304));
    InMux I__302 (
            .O(N__2976),
            .I(N__2973));
    LocalMux I__301 (
            .O(N__2973),
            .I(n14));
    InMux I__300 (
            .O(N__2970),
            .I(n2305));
    InMux I__299 (
            .O(N__2967),
            .I(N__2964));
    LocalMux I__298 (
            .O(N__2964),
            .I(n13));
    InMux I__297 (
            .O(N__2961),
            .I(n2306));
    InMux I__296 (
            .O(N__2958),
            .I(N__2955));
    LocalMux I__295 (
            .O(N__2955),
            .I(n12));
    InMux I__294 (
            .O(N__2952),
            .I(n2307));
    InMux I__293 (
            .O(N__2949),
            .I(N__2946));
    LocalMux I__292 (
            .O(N__2946),
            .I(n11));
    InMux I__291 (
            .O(N__2943),
            .I(n2308));
    InMux I__290 (
            .O(N__2940),
            .I(N__2937));
    LocalMux I__289 (
            .O(N__2937),
            .I(n10));
    InMux I__288 (
            .O(N__2934),
            .I(bfn_14_23_0_));
    InMux I__287 (
            .O(N__2931),
            .I(N__2928));
    LocalMux I__286 (
            .O(N__2928),
            .I(n9));
    InMux I__285 (
            .O(N__2925),
            .I(n2310));
    InMux I__284 (
            .O(N__2922),
            .I(N__2919));
    LocalMux I__283 (
            .O(N__2919),
            .I(n8_adj_409));
    InMux I__282 (
            .O(N__2916),
            .I(n2311));
    InMux I__281 (
            .O(N__2913),
            .I(N__2910));
    LocalMux I__280 (
            .O(N__2910),
            .I(n24));
    InMux I__279 (
            .O(N__2907),
            .I(n2295));
    InMux I__278 (
            .O(N__2904),
            .I(N__2901));
    LocalMux I__277 (
            .O(N__2901),
            .I(n23));
    InMux I__276 (
            .O(N__2898),
            .I(n2296));
    InMux I__275 (
            .O(N__2895),
            .I(N__2892));
    LocalMux I__274 (
            .O(N__2892),
            .I(n22));
    InMux I__273 (
            .O(N__2889),
            .I(n2297));
    InMux I__272 (
            .O(N__2886),
            .I(N__2883));
    LocalMux I__271 (
            .O(N__2883),
            .I(n21));
    InMux I__270 (
            .O(N__2880),
            .I(n2298));
    InMux I__269 (
            .O(N__2877),
            .I(N__2874));
    LocalMux I__268 (
            .O(N__2874),
            .I(n20));
    InMux I__267 (
            .O(N__2871),
            .I(n2299));
    InMux I__266 (
            .O(N__2868),
            .I(N__2865));
    LocalMux I__265 (
            .O(N__2865),
            .I(n19));
    InMux I__264 (
            .O(N__2862),
            .I(n2300));
    InMux I__263 (
            .O(N__2859),
            .I(N__2856));
    LocalMux I__262 (
            .O(N__2856),
            .I(n18));
    InMux I__261 (
            .O(N__2853),
            .I(bfn_14_22_0_));
    InMux I__260 (
            .O(N__2850),
            .I(N__2847));
    LocalMux I__259 (
            .O(N__2847),
            .I(n17));
    InMux I__258 (
            .O(N__2844),
            .I(n2302));
    CascadeMux I__257 (
            .O(N__2841),
            .I(n2553_cascade_));
    IoInMux I__256 (
            .O(N__2838),
            .I(N__2835));
    LocalMux I__255 (
            .O(N__2835),
            .I(N__2832));
    Span12Mux_s9_v I__254 (
            .O(N__2832),
            .I(N__2829));
    Odrv12 I__253 (
            .O(N__2829),
            .I(LED_c));
    InMux I__252 (
            .O(N__2826),
            .I(N__2823));
    LocalMux I__251 (
            .O(N__2823),
            .I(n2554));
    InMux I__250 (
            .O(N__2820),
            .I(N__2817));
    LocalMux I__249 (
            .O(N__2817),
            .I(n26));
    InMux I__248 (
            .O(N__2814),
            .I(bfn_14_21_0_));
    InMux I__247 (
            .O(N__2811),
            .I(N__2808));
    LocalMux I__246 (
            .O(N__2808),
            .I(n25));
    InMux I__245 (
            .O(N__2805),
            .I(n2294));
    IoInMux I__244 (
            .O(N__2802),
            .I(N__2799));
    LocalMux I__243 (
            .O(N__2799),
            .I(N__2796));
    IoSpan4Mux I__242 (
            .O(N__2796),
            .I(N__2793));
    IoSpan4Mux I__241 (
            .O(N__2793),
            .I(N__2790));
    IoSpan4Mux I__240 (
            .O(N__2790),
            .I(N__2787));
    Odrv4 I__239 (
            .O(N__2787),
            .I(CLK_pad_gb_input));
    INV \INVeeprom.i2c.i2c_scl_enable_124C  (
            .O(\INVeeprom.i2c.i2c_scl_enable_124C_net ),
            .I(N__6181));
    INV \INVeeprom.i2c.sda_out_133C  (
            .O(\INVeeprom.i2c.sda_out_133C_net ),
            .I(N__6153));
    INV \INVeeprom.i2c.write_enable_132C  (
            .O(\INVeeprom.i2c.write_enable_132C_net ),
            .I(N__6129));
    defparam IN_MUX_bfv_21_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_22_0_));
    defparam IN_MUX_bfv_21_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_18_0_));
    defparam IN_MUX_bfv_18_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_17_0_));
    defparam IN_MUX_bfv_18_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_18_0_ (
            .carryinitin(\eeprom.n2248 ),
            .carryinitout(bfn_18_18_0_));
    defparam IN_MUX_bfv_17_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_21_0_));
    defparam IN_MUX_bfv_17_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_22_0_ (
            .carryinitin(n2270),
            .carryinitout(bfn_17_22_0_));
    defparam IN_MUX_bfv_17_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_23_0_ (
            .carryinitin(n2278),
            .carryinitout(bfn_17_23_0_));
    defparam IN_MUX_bfv_17_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_24_0_ (
            .carryinitin(n2286),
            .carryinitout(bfn_17_24_0_));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_21_0_));
    defparam IN_MUX_bfv_14_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_22_0_ (
            .carryinitin(n2301),
            .carryinitout(bfn_14_22_0_));
    defparam IN_MUX_bfv_14_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_23_0_ (
            .carryinitin(n2309),
            .carryinitout(bfn_14_23_0_));
    defparam IN_MUX_bfv_14_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_24_0_ (
            .carryinitin(n2317),
            .carryinitout(bfn_14_24_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__2802),
            .GLOBALBUFFEROUTPUT(CLK_N));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam i1635_4_lut_LC_13_23_3.C_ON=1'b0;
    defparam i1635_4_lut_LC_13_23_3.SEQ_MODE=4'b0000;
    defparam i1635_4_lut_LC_13_23_3.LUT_INIT=16'b1101110101000000;
    LogicCell40 i1635_4_lut_LC_13_23_3 (
            .in0(N__3026),
            .in1(N__3068),
            .in2(N__3050),
            .in3(N__3086),
            .lcout(),
            .ltout(n2553_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1637_3_lut_LC_13_23_4.C_ON=1'b0;
    defparam i1637_3_lut_LC_13_23_4.SEQ_MODE=4'b0000;
    defparam i1637_3_lut_LC_13_23_4.LUT_INIT=16'b0101010100001111;
    LogicCell40 i1637_3_lut_LC_13_23_4 (
            .in0(N__2826),
            .in1(_gnd_net_),
            .in2(N__2841),
            .in3(N__3006),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1636_4_lut_LC_13_23_5.C_ON=1'b0;
    defparam i1636_4_lut_LC_13_23_5.SEQ_MODE=4'b0000;
    defparam i1636_4_lut_LC_13_23_5.LUT_INIT=16'b1111111010110000;
    LogicCell40 i1636_4_lut_LC_13_23_5 (
            .in0(N__3027),
            .in1(N__3069),
            .in2(N__3051),
            .in3(N__3087),
            .lcout(n2554),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i0_LC_14_21_0.C_ON=1'b1;
    defparam blink_counter_363__i0_LC_14_21_0.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i0_LC_14_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i0_LC_14_21_0 (
            .in0(_gnd_net_),
            .in1(N__2820),
            .in2(_gnd_net_),
            .in3(N__2814),
            .lcout(n26),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(n2294),
            .clk(N__5117),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i1_LC_14_21_1.C_ON=1'b1;
    defparam blink_counter_363__i1_LC_14_21_1.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i1_LC_14_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i1_LC_14_21_1 (
            .in0(_gnd_net_),
            .in1(N__2811),
            .in2(_gnd_net_),
            .in3(N__2805),
            .lcout(n25),
            .ltout(),
            .carryin(n2294),
            .carryout(n2295),
            .clk(N__5117),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i2_LC_14_21_2.C_ON=1'b1;
    defparam blink_counter_363__i2_LC_14_21_2.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i2_LC_14_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i2_LC_14_21_2 (
            .in0(_gnd_net_),
            .in1(N__2913),
            .in2(_gnd_net_),
            .in3(N__2907),
            .lcout(n24),
            .ltout(),
            .carryin(n2295),
            .carryout(n2296),
            .clk(N__5117),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i3_LC_14_21_3.C_ON=1'b1;
    defparam blink_counter_363__i3_LC_14_21_3.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i3_LC_14_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i3_LC_14_21_3 (
            .in0(_gnd_net_),
            .in1(N__2904),
            .in2(_gnd_net_),
            .in3(N__2898),
            .lcout(n23),
            .ltout(),
            .carryin(n2296),
            .carryout(n2297),
            .clk(N__5117),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i4_LC_14_21_4.C_ON=1'b1;
    defparam blink_counter_363__i4_LC_14_21_4.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i4_LC_14_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i4_LC_14_21_4 (
            .in0(_gnd_net_),
            .in1(N__2895),
            .in2(_gnd_net_),
            .in3(N__2889),
            .lcout(n22),
            .ltout(),
            .carryin(n2297),
            .carryout(n2298),
            .clk(N__5117),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i5_LC_14_21_5.C_ON=1'b1;
    defparam blink_counter_363__i5_LC_14_21_5.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i5_LC_14_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i5_LC_14_21_5 (
            .in0(_gnd_net_),
            .in1(N__2886),
            .in2(_gnd_net_),
            .in3(N__2880),
            .lcout(n21),
            .ltout(),
            .carryin(n2298),
            .carryout(n2299),
            .clk(N__5117),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i6_LC_14_21_6.C_ON=1'b1;
    defparam blink_counter_363__i6_LC_14_21_6.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i6_LC_14_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i6_LC_14_21_6 (
            .in0(_gnd_net_),
            .in1(N__2877),
            .in2(_gnd_net_),
            .in3(N__2871),
            .lcout(n20),
            .ltout(),
            .carryin(n2299),
            .carryout(n2300),
            .clk(N__5117),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i7_LC_14_21_7.C_ON=1'b1;
    defparam blink_counter_363__i7_LC_14_21_7.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i7_LC_14_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i7_LC_14_21_7 (
            .in0(_gnd_net_),
            .in1(N__2868),
            .in2(_gnd_net_),
            .in3(N__2862),
            .lcout(n19),
            .ltout(),
            .carryin(n2300),
            .carryout(n2301),
            .clk(N__5117),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i8_LC_14_22_0.C_ON=1'b1;
    defparam blink_counter_363__i8_LC_14_22_0.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i8_LC_14_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i8_LC_14_22_0 (
            .in0(_gnd_net_),
            .in1(N__2859),
            .in2(_gnd_net_),
            .in3(N__2853),
            .lcout(n18),
            .ltout(),
            .carryin(bfn_14_22_0_),
            .carryout(n2302),
            .clk(N__5120),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i9_LC_14_22_1.C_ON=1'b1;
    defparam blink_counter_363__i9_LC_14_22_1.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i9_LC_14_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i9_LC_14_22_1 (
            .in0(_gnd_net_),
            .in1(N__2850),
            .in2(_gnd_net_),
            .in3(N__2844),
            .lcout(n17),
            .ltout(),
            .carryin(n2302),
            .carryout(n2303),
            .clk(N__5120),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i10_LC_14_22_2.C_ON=1'b1;
    defparam blink_counter_363__i10_LC_14_22_2.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i10_LC_14_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i10_LC_14_22_2 (
            .in0(_gnd_net_),
            .in1(N__2994),
            .in2(_gnd_net_),
            .in3(N__2988),
            .lcout(n16),
            .ltout(),
            .carryin(n2303),
            .carryout(n2304),
            .clk(N__5120),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i11_LC_14_22_3.C_ON=1'b1;
    defparam blink_counter_363__i11_LC_14_22_3.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i11_LC_14_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i11_LC_14_22_3 (
            .in0(_gnd_net_),
            .in1(N__2985),
            .in2(_gnd_net_),
            .in3(N__2979),
            .lcout(n15),
            .ltout(),
            .carryin(n2304),
            .carryout(n2305),
            .clk(N__5120),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i12_LC_14_22_4.C_ON=1'b1;
    defparam blink_counter_363__i12_LC_14_22_4.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i12_LC_14_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i12_LC_14_22_4 (
            .in0(_gnd_net_),
            .in1(N__2976),
            .in2(_gnd_net_),
            .in3(N__2970),
            .lcout(n14),
            .ltout(),
            .carryin(n2305),
            .carryout(n2306),
            .clk(N__5120),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i13_LC_14_22_5.C_ON=1'b1;
    defparam blink_counter_363__i13_LC_14_22_5.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i13_LC_14_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i13_LC_14_22_5 (
            .in0(_gnd_net_),
            .in1(N__2967),
            .in2(_gnd_net_),
            .in3(N__2961),
            .lcout(n13),
            .ltout(),
            .carryin(n2306),
            .carryout(n2307),
            .clk(N__5120),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i14_LC_14_22_6.C_ON=1'b1;
    defparam blink_counter_363__i14_LC_14_22_6.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i14_LC_14_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i14_LC_14_22_6 (
            .in0(_gnd_net_),
            .in1(N__2958),
            .in2(_gnd_net_),
            .in3(N__2952),
            .lcout(n12),
            .ltout(),
            .carryin(n2307),
            .carryout(n2308),
            .clk(N__5120),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i15_LC_14_22_7.C_ON=1'b1;
    defparam blink_counter_363__i15_LC_14_22_7.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i15_LC_14_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i15_LC_14_22_7 (
            .in0(_gnd_net_),
            .in1(N__2949),
            .in2(_gnd_net_),
            .in3(N__2943),
            .lcout(n11),
            .ltout(),
            .carryin(n2308),
            .carryout(n2309),
            .clk(N__5120),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i16_LC_14_23_0.C_ON=1'b1;
    defparam blink_counter_363__i16_LC_14_23_0.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i16_LC_14_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i16_LC_14_23_0 (
            .in0(_gnd_net_),
            .in1(N__2940),
            .in2(_gnd_net_),
            .in3(N__2934),
            .lcout(n10),
            .ltout(),
            .carryin(bfn_14_23_0_),
            .carryout(n2310),
            .clk(N__5122),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i17_LC_14_23_1.C_ON=1'b1;
    defparam blink_counter_363__i17_LC_14_23_1.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i17_LC_14_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i17_LC_14_23_1 (
            .in0(_gnd_net_),
            .in1(N__2931),
            .in2(_gnd_net_),
            .in3(N__2925),
            .lcout(n9),
            .ltout(),
            .carryin(n2310),
            .carryout(n2311),
            .clk(N__5122),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i18_LC_14_23_2.C_ON=1'b1;
    defparam blink_counter_363__i18_LC_14_23_2.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i18_LC_14_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i18_LC_14_23_2 (
            .in0(_gnd_net_),
            .in1(N__2922),
            .in2(_gnd_net_),
            .in3(N__2916),
            .lcout(n8_adj_409),
            .ltout(),
            .carryin(n2311),
            .carryout(n2312),
            .clk(N__5122),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i19_LC_14_23_3.C_ON=1'b1;
    defparam blink_counter_363__i19_LC_14_23_3.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i19_LC_14_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i19_LC_14_23_3 (
            .in0(_gnd_net_),
            .in1(N__3105),
            .in2(_gnd_net_),
            .in3(N__3099),
            .lcout(n7),
            .ltout(),
            .carryin(n2312),
            .carryout(n2313),
            .clk(N__5122),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i20_LC_14_23_4.C_ON=1'b1;
    defparam blink_counter_363__i20_LC_14_23_4.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i20_LC_14_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i20_LC_14_23_4 (
            .in0(_gnd_net_),
            .in1(N__3096),
            .in2(_gnd_net_),
            .in3(N__3090),
            .lcout(n6_adj_410),
            .ltout(),
            .carryin(n2313),
            .carryout(n2314),
            .clk(N__5122),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i21_LC_14_23_5.C_ON=1'b1;
    defparam blink_counter_363__i21_LC_14_23_5.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i21_LC_14_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i21_LC_14_23_5 (
            .in0(_gnd_net_),
            .in1(N__3085),
            .in2(_gnd_net_),
            .in3(N__3072),
            .lcout(blink_counter_21),
            .ltout(),
            .carryin(n2314),
            .carryout(n2315),
            .clk(N__5122),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i22_LC_14_23_6.C_ON=1'b1;
    defparam blink_counter_363__i22_LC_14_23_6.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i22_LC_14_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i22_LC_14_23_6 (
            .in0(_gnd_net_),
            .in1(N__3067),
            .in2(_gnd_net_),
            .in3(N__3054),
            .lcout(blink_counter_22),
            .ltout(),
            .carryin(n2315),
            .carryout(n2316),
            .clk(N__5122),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i23_LC_14_23_7.C_ON=1'b1;
    defparam blink_counter_363__i23_LC_14_23_7.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i23_LC_14_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i23_LC_14_23_7 (
            .in0(_gnd_net_),
            .in1(N__3043),
            .in2(_gnd_net_),
            .in3(N__3030),
            .lcout(blink_counter_23),
            .ltout(),
            .carryin(n2316),
            .carryout(n2317),
            .clk(N__5122),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i24_LC_14_24_0.C_ON=1'b1;
    defparam blink_counter_363__i24_LC_14_24_0.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i24_LC_14_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i24_LC_14_24_0 (
            .in0(_gnd_net_),
            .in1(N__3025),
            .in2(_gnd_net_),
            .in3(N__3012),
            .lcout(blink_counter_24),
            .ltout(),
            .carryin(bfn_14_24_0_),
            .carryout(n2318),
            .clk(N__5126),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_363__i25_LC_14_24_1.C_ON=1'b0;
    defparam blink_counter_363__i25_LC_14_24_1.SEQ_MODE=4'b1000;
    defparam blink_counter_363__i25_LC_14_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_363__i25_LC_14_24_1 (
            .in0(_gnd_net_),
            .in1(N__3005),
            .in2(_gnd_net_),
            .in3(N__3009),
            .lcout(blink_counter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5126),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.enable_39_LC_17_18_0 .C_ON=1'b0;
    defparam \eeprom.enable_39_LC_17_18_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.enable_39_LC_17_18_0 .LUT_INIT=16'b0011011100000100;
    LogicCell40 \eeprom.enable_39_LC_17_18_0  (
            .in0(N__3604),
            .in1(N__4538),
            .in2(N__5952),
            .in3(N__4221),
            .lcout(\eeprom.enable ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5118),
            .ce(),
            .sr(N__3960));
    defparam \eeprom.i1696_2_lut_LC_17_18_1 .C_ON=1'b0;
    defparam \eeprom.i1696_2_lut_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1696_2_lut_LC_17_18_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \eeprom.i1696_2_lut_LC_17_18_1  (
            .in0(_gnd_net_),
            .in1(N__5951),
            .in2(_gnd_net_),
            .in3(N__3603),
            .lcout(\eeprom.n642 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i6_4_lut_LC_17_19_0 .C_ON=1'b0;
    defparam \eeprom.i6_4_lut_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i6_4_lut_LC_17_19_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i6_4_lut_LC_17_19_0  (
            .in0(N__3226),
            .in1(N__3277),
            .in2(N__3347),
            .in3(N__3310),
            .lcout(\eeprom.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_i0_i12_LC_17_19_1 .C_ON=1'b0;
    defparam \eeprom.delay_counter_i0_i12_LC_17_19_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i12_LC_17_19_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \eeprom.delay_counter_i0_i12_LC_17_19_1  (
            .in0(N__3278),
            .in1(N__4530),
            .in2(N__3264),
            .in3(N__4342),
            .lcout(\eeprom.delay_counter_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5121),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_i0_i8_LC_17_19_2 .C_ON=1'b0;
    defparam \eeprom.delay_counter_i0_i8_LC_17_19_2 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i8_LC_17_19_2 .LUT_INIT=16'b1101111111010000;
    LogicCell40 \eeprom.delay_counter_i0_i8_LC_17_19_2  (
            .in0(N__4531),
            .in1(N__3297),
            .in2(N__4371),
            .in3(N__3311),
            .lcout(\eeprom.delay_counter_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5121),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_i0_i6_LC_17_19_4 .C_ON=1'b0;
    defparam \eeprom.delay_counter_i0_i6_LC_17_19_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i6_LC_17_19_4 .LUT_INIT=16'b1111101000111010;
    LogicCell40 \eeprom.delay_counter_i0_i6_LC_17_19_4  (
            .in0(N__3343),
            .in1(N__4529),
            .in2(N__4370),
            .in3(N__3327),
            .lcout(\eeprom.delay_counter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5121),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_i0_i2_LC_17_19_6 .C_ON=1'b0;
    defparam \eeprom.delay_counter_i0_i2_LC_17_19_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i2_LC_17_19_6 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \eeprom.delay_counter_i0_i2_LC_17_19_6  (
            .in0(N__3227),
            .in1(N__4349),
            .in2(N__3213),
            .in3(N__4528),
            .lcout(\eeprom.delay_counter_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5121),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.mux_182_Mux_0_i1_4_lut_LC_17_20_2 .C_ON=1'b0;
    defparam \eeprom.mux_182_Mux_0_i1_4_lut_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.mux_182_Mux_0_i1_4_lut_LC_17_20_2 .LUT_INIT=16'b0100010001001110;
    LogicCell40 \eeprom.mux_182_Mux_0_i1_4_lut_LC_17_20_2  (
            .in0(N__4473),
            .in1(N__4220),
            .in2(N__5946),
            .in3(N__3606),
            .lcout(),
            .ltout(n693_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.rw_43_LC_17_20_3 .C_ON=1'b0;
    defparam \eeprom.rw_43_LC_17_20_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.rw_43_LC_17_20_3 .LUT_INIT=16'b1011101010001010;
    LogicCell40 \eeprom.rw_43_LC_17_20_3  (
            .in0(N__4763),
            .in1(N__3952),
            .in2(N__3111),
            .in3(N__4474),
            .lcout(rw),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5123),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_3_lut_adj_13_LC_17_20_5 .C_ON=1'b0;
    defparam \eeprom.i1_3_lut_adj_13_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_3_lut_adj_13_LC_17_20_5 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \eeprom.i1_3_lut_adj_13_LC_17_20_5  (
            .in0(N__4219),
            .in1(N__3951),
            .in2(_gnd_net_),
            .in3(N__4472),
            .lcout(\eeprom.n1601 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_counter_362__i0_LC_17_21_0.C_ON=1'b1;
    defparam delay_counter_362__i0_LC_17_21_0.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i0_LC_17_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i0_LC_17_21_0 (
            .in0(_gnd_net_),
            .in1(N__3726),
            .in2(_gnd_net_),
            .in3(N__3108),
            .lcout(delay_counter_0),
            .ltout(),
            .carryin(bfn_17_21_0_),
            .carryout(n2263),
            .clk(N__5127),
            .ce(),
            .sr(N__4116));
    defparam delay_counter_362__i1_LC_17_21_1.C_ON=1'b1;
    defparam delay_counter_362__i1_LC_17_21_1.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i1_LC_17_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i1_LC_17_21_1 (
            .in0(_gnd_net_),
            .in1(N__3884),
            .in2(_gnd_net_),
            .in3(N__3138),
            .lcout(delay_counter_1),
            .ltout(),
            .carryin(n2263),
            .carryout(n2264),
            .clk(N__5127),
            .ce(),
            .sr(N__4116));
    defparam delay_counter_362__i2_LC_17_21_2.C_ON=1'b1;
    defparam delay_counter_362__i2_LC_17_21_2.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i2_LC_17_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i2_LC_17_21_2 (
            .in0(_gnd_net_),
            .in1(N__4247),
            .in2(_gnd_net_),
            .in3(N__3135),
            .lcout(delay_counter_2),
            .ltout(),
            .carryin(n2264),
            .carryout(n2265),
            .clk(N__5127),
            .ce(),
            .sr(N__4116));
    defparam delay_counter_362__i3_LC_17_21_3.C_ON=1'b1;
    defparam delay_counter_362__i3_LC_17_21_3.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i3_LC_17_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i3_LC_17_21_3 (
            .in0(_gnd_net_),
            .in1(N__3740),
            .in2(_gnd_net_),
            .in3(N__3132),
            .lcout(delay_counter_3),
            .ltout(),
            .carryin(n2265),
            .carryout(n2266),
            .clk(N__5127),
            .ce(),
            .sr(N__4116));
    defparam delay_counter_362__i4_LC_17_21_4.C_ON=1'b1;
    defparam delay_counter_362__i4_LC_17_21_4.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i4_LC_17_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i4_LC_17_21_4 (
            .in0(_gnd_net_),
            .in1(N__3870),
            .in2(_gnd_net_),
            .in3(N__3129),
            .lcout(delay_counter_4),
            .ltout(),
            .carryin(n2266),
            .carryout(n2267),
            .clk(N__5127),
            .ce(),
            .sr(N__4116));
    defparam delay_counter_362__i5_LC_17_21_5.C_ON=1'b1;
    defparam delay_counter_362__i5_LC_17_21_5.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i5_LC_17_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i5_LC_17_21_5 (
            .in0(_gnd_net_),
            .in1(N__4271),
            .in2(_gnd_net_),
            .in3(N__3126),
            .lcout(delay_counter_5),
            .ltout(),
            .carryin(n2267),
            .carryout(n2268),
            .clk(N__5127),
            .ce(),
            .sr(N__4116));
    defparam delay_counter_362__i6_LC_17_21_6.C_ON=1'b1;
    defparam delay_counter_362__i6_LC_17_21_6.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i6_LC_17_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i6_LC_17_21_6 (
            .in0(_gnd_net_),
            .in1(N__3753),
            .in2(_gnd_net_),
            .in3(N__3123),
            .lcout(delay_counter_6),
            .ltout(),
            .carryin(n2268),
            .carryout(n2269),
            .clk(N__5127),
            .ce(),
            .sr(N__4116));
    defparam delay_counter_362__i7_LC_17_21_7.C_ON=1'b1;
    defparam delay_counter_362__i7_LC_17_21_7.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i7_LC_17_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i7_LC_17_21_7 (
            .in0(_gnd_net_),
            .in1(N__3909),
            .in2(_gnd_net_),
            .in3(N__3120),
            .lcout(delay_counter_7),
            .ltout(),
            .carryin(n2269),
            .carryout(n2270),
            .clk(N__5127),
            .ce(),
            .sr(N__4116));
    defparam delay_counter_362__i8_LC_17_22_0.C_ON=1'b1;
    defparam delay_counter_362__i8_LC_17_22_0.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i8_LC_17_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i8_LC_17_22_0 (
            .in0(_gnd_net_),
            .in1(N__3897),
            .in2(_gnd_net_),
            .in3(N__3117),
            .lcout(delay_counter_8),
            .ltout(),
            .carryin(bfn_17_22_0_),
            .carryout(n2271),
            .clk(N__5130),
            .ce(),
            .sr(N__4111));
    defparam delay_counter_362__i9_LC_17_22_1.C_ON=1'b1;
    defparam delay_counter_362__i9_LC_17_22_1.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i9_LC_17_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i9_LC_17_22_1 (
            .in0(_gnd_net_),
            .in1(N__3765),
            .in2(_gnd_net_),
            .in3(N__3114),
            .lcout(delay_counter_9),
            .ltout(),
            .carryin(n2271),
            .carryout(n2272),
            .clk(N__5130),
            .ce(),
            .sr(N__4111));
    defparam delay_counter_362__i10_LC_17_22_2.C_ON=1'b1;
    defparam delay_counter_362__i10_LC_17_22_2.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i10_LC_17_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i10_LC_17_22_2 (
            .in0(_gnd_net_),
            .in1(N__3858),
            .in2(_gnd_net_),
            .in3(N__3165),
            .lcout(delay_counter_10),
            .ltout(),
            .carryin(n2272),
            .carryout(n2273),
            .clk(N__5130),
            .ce(),
            .sr(N__4111));
    defparam delay_counter_362__i11_LC_17_22_3.C_ON=1'b1;
    defparam delay_counter_362__i11_LC_17_22_3.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i11_LC_17_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i11_LC_17_22_3 (
            .in0(_gnd_net_),
            .in1(N__3833),
            .in2(_gnd_net_),
            .in3(N__3162),
            .lcout(delay_counter_11),
            .ltout(),
            .carryin(n2273),
            .carryout(n2274),
            .clk(N__5130),
            .ce(),
            .sr(N__4111));
    defparam delay_counter_362__i12_LC_17_22_4.C_ON=1'b1;
    defparam delay_counter_362__i12_LC_17_22_4.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i12_LC_17_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i12_LC_17_22_4 (
            .in0(_gnd_net_),
            .in1(N__3846),
            .in2(_gnd_net_),
            .in3(N__3159),
            .lcout(delay_counter_12),
            .ltout(),
            .carryin(n2274),
            .carryout(n2275),
            .clk(N__5130),
            .ce(),
            .sr(N__4111));
    defparam delay_counter_362__i13_LC_17_22_5.C_ON=1'b1;
    defparam delay_counter_362__i13_LC_17_22_5.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i13_LC_17_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i13_LC_17_22_5 (
            .in0(_gnd_net_),
            .in1(N__3819),
            .in2(_gnd_net_),
            .in3(N__3156),
            .lcout(delay_counter_13),
            .ltout(),
            .carryin(n2275),
            .carryout(n2276),
            .clk(N__5130),
            .ce(),
            .sr(N__4111));
    defparam delay_counter_362__i14_LC_17_22_6.C_ON=1'b1;
    defparam delay_counter_362__i14_LC_17_22_6.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i14_LC_17_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i14_LC_17_22_6 (
            .in0(_gnd_net_),
            .in1(N__3690),
            .in2(_gnd_net_),
            .in3(N__3153),
            .lcout(delay_counter_14),
            .ltout(),
            .carryin(n2276),
            .carryout(n2277),
            .clk(N__5130),
            .ce(),
            .sr(N__4111));
    defparam delay_counter_362__i15_LC_17_22_7.C_ON=1'b1;
    defparam delay_counter_362__i15_LC_17_22_7.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i15_LC_17_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i15_LC_17_22_7 (
            .in0(_gnd_net_),
            .in1(N__3702),
            .in2(_gnd_net_),
            .in3(N__3150),
            .lcout(delay_counter_15),
            .ltout(),
            .carryin(n2277),
            .carryout(n2278),
            .clk(N__5130),
            .ce(),
            .sr(N__4111));
    defparam delay_counter_362__i16_LC_17_23_0.C_ON=1'b1;
    defparam delay_counter_362__i16_LC_17_23_0.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i16_LC_17_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i16_LC_17_23_0 (
            .in0(_gnd_net_),
            .in1(N__3804),
            .in2(_gnd_net_),
            .in3(N__3147),
            .lcout(delay_counter_16),
            .ltout(),
            .carryin(bfn_17_23_0_),
            .carryout(n2279),
            .clk(N__5134),
            .ce(),
            .sr(N__4101));
    defparam delay_counter_362__i17_LC_17_23_1.C_ON=1'b1;
    defparam delay_counter_362__i17_LC_17_23_1.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i17_LC_17_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i17_LC_17_23_1 (
            .in0(_gnd_net_),
            .in1(N__3714),
            .in2(_gnd_net_),
            .in3(N__3144),
            .lcout(delay_counter_17),
            .ltout(),
            .carryin(n2279),
            .carryout(n2280),
            .clk(N__5134),
            .ce(),
            .sr(N__4101));
    defparam delay_counter_362__i18_LC_17_23_2.C_ON=1'b1;
    defparam delay_counter_362__i18_LC_17_23_2.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i18_LC_17_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i18_LC_17_23_2 (
            .in0(_gnd_net_),
            .in1(N__3792),
            .in2(_gnd_net_),
            .in3(N__3141),
            .lcout(delay_counter_18),
            .ltout(),
            .carryin(n2280),
            .carryout(n2281),
            .clk(N__5134),
            .ce(),
            .sr(N__4101));
    defparam delay_counter_362__i19_LC_17_23_3.C_ON=1'b1;
    defparam delay_counter_362__i19_LC_17_23_3.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i19_LC_17_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i19_LC_17_23_3 (
            .in0(_gnd_net_),
            .in1(N__3777),
            .in2(_gnd_net_),
            .in3(N__3192),
            .lcout(delay_counter_19),
            .ltout(),
            .carryin(n2281),
            .carryout(n2282),
            .clk(N__5134),
            .ce(),
            .sr(N__4101));
    defparam delay_counter_362__i20_LC_17_23_4.C_ON=1'b1;
    defparam delay_counter_362__i20_LC_17_23_4.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i20_LC_17_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i20_LC_17_23_4 (
            .in0(_gnd_net_),
            .in1(N__4163),
            .in2(_gnd_net_),
            .in3(N__3189),
            .lcout(delay_counter_20),
            .ltout(),
            .carryin(n2282),
            .carryout(n2283),
            .clk(N__5134),
            .ce(),
            .sr(N__4101));
    defparam delay_counter_362__i21_LC_17_23_5.C_ON=1'b1;
    defparam delay_counter_362__i21_LC_17_23_5.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i21_LC_17_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i21_LC_17_23_5 (
            .in0(_gnd_net_),
            .in1(N__3672),
            .in2(_gnd_net_),
            .in3(N__3186),
            .lcout(delay_counter_21),
            .ltout(),
            .carryin(n2283),
            .carryout(n2284),
            .clk(N__5134),
            .ce(),
            .sr(N__4101));
    defparam delay_counter_362__i22_LC_17_23_6.C_ON=1'b1;
    defparam delay_counter_362__i22_LC_17_23_6.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i22_LC_17_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i22_LC_17_23_6 (
            .in0(_gnd_net_),
            .in1(N__4188),
            .in2(_gnd_net_),
            .in3(N__3183),
            .lcout(delay_counter_22),
            .ltout(),
            .carryin(n2284),
            .carryout(n2285),
            .clk(N__5134),
            .ce(),
            .sr(N__4101));
    defparam delay_counter_362__i23_LC_17_23_7.C_ON=1'b1;
    defparam delay_counter_362__i23_LC_17_23_7.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i23_LC_17_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i23_LC_17_23_7 (
            .in0(_gnd_net_),
            .in1(N__3660),
            .in2(_gnd_net_),
            .in3(N__3180),
            .lcout(delay_counter_23),
            .ltout(),
            .carryin(n2285),
            .carryout(n2286),
            .clk(N__5134),
            .ce(),
            .sr(N__4101));
    defparam delay_counter_362__i24_LC_17_24_0.C_ON=1'b1;
    defparam delay_counter_362__i24_LC_17_24_0.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i24_LC_17_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i24_LC_17_24_0 (
            .in0(_gnd_net_),
            .in1(N__3999),
            .in2(_gnd_net_),
            .in3(N__3177),
            .lcout(delay_counter_24),
            .ltout(),
            .carryin(bfn_17_24_0_),
            .carryout(n2287),
            .clk(N__5135),
            .ce(),
            .sr(N__4112));
    defparam delay_counter_362__i25_LC_17_24_1.C_ON=1'b1;
    defparam delay_counter_362__i25_LC_17_24_1.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i25_LC_17_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i25_LC_17_24_1 (
            .in0(_gnd_net_),
            .in1(N__4176),
            .in2(_gnd_net_),
            .in3(N__3174),
            .lcout(delay_counter_25),
            .ltout(),
            .carryin(n2287),
            .carryout(n2288),
            .clk(N__5135),
            .ce(),
            .sr(N__4112));
    defparam delay_counter_362__i26_LC_17_24_2.C_ON=1'b1;
    defparam delay_counter_362__i26_LC_17_24_2.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i26_LC_17_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i26_LC_17_24_2 (
            .in0(_gnd_net_),
            .in1(N__4038),
            .in2(_gnd_net_),
            .in3(N__3171),
            .lcout(delay_counter_26),
            .ltout(),
            .carryin(n2288),
            .carryout(n2289),
            .clk(N__5135),
            .ce(),
            .sr(N__4112));
    defparam delay_counter_362__i27_LC_17_24_3.C_ON=1'b1;
    defparam delay_counter_362__i27_LC_17_24_3.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i27_LC_17_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i27_LC_17_24_3 (
            .in0(_gnd_net_),
            .in1(N__4013),
            .in2(_gnd_net_),
            .in3(N__3168),
            .lcout(delay_counter_27),
            .ltout(),
            .carryin(n2289),
            .carryout(n2290),
            .clk(N__5135),
            .ce(),
            .sr(N__4112));
    defparam delay_counter_362__i28_LC_17_24_4.C_ON=1'b1;
    defparam delay_counter_362__i28_LC_17_24_4.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i28_LC_17_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i28_LC_17_24_4 (
            .in0(_gnd_net_),
            .in1(N__4062),
            .in2(_gnd_net_),
            .in3(N__3249),
            .lcout(delay_counter_28),
            .ltout(),
            .carryin(n2290),
            .carryout(n2291),
            .clk(N__5135),
            .ce(),
            .sr(N__4112));
    defparam delay_counter_362__i29_LC_17_24_5.C_ON=1'b1;
    defparam delay_counter_362__i29_LC_17_24_5.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i29_LC_17_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i29_LC_17_24_5 (
            .in0(_gnd_net_),
            .in1(N__4074),
            .in2(_gnd_net_),
            .in3(N__3246),
            .lcout(delay_counter_29),
            .ltout(),
            .carryin(n2291),
            .carryout(n2292),
            .clk(N__5135),
            .ce(),
            .sr(N__4112));
    defparam delay_counter_362__i30_LC_17_24_6.C_ON=1'b1;
    defparam delay_counter_362__i30_LC_17_24_6.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i30_LC_17_24_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i30_LC_17_24_6 (
            .in0(_gnd_net_),
            .in1(N__4026),
            .in2(_gnd_net_),
            .in3(N__3243),
            .lcout(delay_counter_30),
            .ltout(),
            .carryin(n2292),
            .carryout(n2293),
            .clk(N__5135),
            .ce(),
            .sr(N__4112));
    defparam delay_counter_362__i31_LC_17_24_7.C_ON=1'b0;
    defparam delay_counter_362__i31_LC_17_24_7.SEQ_MODE=4'b1000;
    defparam delay_counter_362__i31_LC_17_24_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 delay_counter_362__i31_LC_17_24_7 (
            .in0(_gnd_net_),
            .in1(N__4135),
            .in2(_gnd_net_),
            .in3(N__3240),
            .lcout(delay_counter_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5135),
            .ce(),
            .sr(N__4112));
    defparam \eeprom.add_158_2_lut_LC_18_17_0 .C_ON=1'b1;
    defparam \eeprom.add_158_2_lut_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_158_2_lut_LC_18_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_158_2_lut_LC_18_17_0  (
            .in0(_gnd_net_),
            .in1(N__3516),
            .in2(N__3426),
            .in3(_gnd_net_),
            .lcout(\eeprom.delay_counter_15_N_171_0 ),
            .ltout(),
            .carryin(bfn_18_17_0_),
            .carryout(\eeprom.n2241 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_158_3_lut_LC_18_17_1 .C_ON=1'b1;
    defparam \eeprom.add_158_3_lut_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_158_3_lut_LC_18_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_158_3_lut_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(N__3453),
            .in2(N__3548),
            .in3(N__3237),
            .lcout(\eeprom.delay_counter_15_N_171_1 ),
            .ltout(),
            .carryin(\eeprom.n2241 ),
            .carryout(\eeprom.n2242 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_158_4_lut_LC_18_17_2 .C_ON=1'b1;
    defparam \eeprom.add_158_4_lut_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_158_4_lut_LC_18_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_158_4_lut_LC_18_17_2  (
            .in0(_gnd_net_),
            .in1(N__3520),
            .in2(N__3234),
            .in3(N__3201),
            .lcout(\eeprom.delay_counter_15_N_171_2 ),
            .ltout(),
            .carryin(\eeprom.n2242 ),
            .carryout(\eeprom.n2243 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_158_5_lut_LC_18_17_3 .C_ON=1'b1;
    defparam \eeprom.add_158_5_lut_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_158_5_lut_LC_18_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_158_5_lut_LC_18_17_3  (
            .in0(_gnd_net_),
            .in1(N__4699),
            .in2(N__3549),
            .in3(N__3198),
            .lcout(\eeprom.delay_counter_15_N_171_3 ),
            .ltout(),
            .carryin(\eeprom.n2243 ),
            .carryout(\eeprom.n2244 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_158_6_lut_LC_18_17_4 .C_ON=1'b1;
    defparam \eeprom.add_158_6_lut_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_158_6_lut_LC_18_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_158_6_lut_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(N__3524),
            .in2(N__3633),
            .in3(N__3195),
            .lcout(\eeprom.delay_counter_15_N_171_4 ),
            .ltout(),
            .carryin(\eeprom.n2244 ),
            .carryout(\eeprom.n2245 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_158_7_lut_LC_18_17_5 .C_ON=1'b1;
    defparam \eeprom.add_158_7_lut_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_158_7_lut_LC_18_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_158_7_lut_LC_18_17_5  (
            .in0(_gnd_net_),
            .in1(N__3396),
            .in2(N__3550),
            .in3(N__3354),
            .lcout(\eeprom.delay_counter_15_N_171_5 ),
            .ltout(),
            .carryin(\eeprom.n2245 ),
            .carryout(\eeprom.n2246 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_158_8_lut_LC_18_17_6 .C_ON=1'b1;
    defparam \eeprom.add_158_8_lut_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_158_8_lut_LC_18_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_158_8_lut_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(N__3528),
            .in2(N__3351),
            .in3(N__3318),
            .lcout(\eeprom.delay_counter_15_N_171_6 ),
            .ltout(),
            .carryin(\eeprom.n2246 ),
            .carryout(\eeprom.n2247 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_158_9_lut_LC_18_17_7 .C_ON=1'b1;
    defparam \eeprom.add_158_9_lut_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_158_9_lut_LC_18_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_158_9_lut_LC_18_17_7  (
            .in0(_gnd_net_),
            .in1(N__4649),
            .in2(N__3551),
            .in3(N__3315),
            .lcout(\eeprom.delay_counter_15_N_171_7 ),
            .ltout(),
            .carryin(\eeprom.n2247 ),
            .carryout(\eeprom.n2248 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_158_10_lut_LC_18_18_0 .C_ON=1'b1;
    defparam \eeprom.add_158_10_lut_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_158_10_lut_LC_18_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_158_10_lut_LC_18_18_0  (
            .in0(_gnd_net_),
            .in1(N__3312),
            .in2(N__3552),
            .in3(N__3291),
            .lcout(\eeprom.delay_counter_15_N_171_8 ),
            .ltout(),
            .carryin(bfn_18_18_0_),
            .carryout(\eeprom.n2249 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_158_11_lut_LC_18_18_1 .C_ON=1'b1;
    defparam \eeprom.add_158_11_lut_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_158_11_lut_LC_18_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_158_11_lut_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(N__3535),
            .in2(N__4622),
            .in3(N__3288),
            .lcout(\eeprom.delay_counter_15_N_171_9 ),
            .ltout(),
            .carryin(\eeprom.n2249 ),
            .carryout(\eeprom.n2250 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_158_12_lut_LC_18_18_2 .C_ON=1'b1;
    defparam \eeprom.add_158_12_lut_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_158_12_lut_LC_18_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_158_12_lut_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(N__3371),
            .in2(N__3553),
            .in3(N__3285),
            .lcout(\eeprom.delay_counter_15_N_171_10 ),
            .ltout(),
            .carryin(\eeprom.n2250 ),
            .carryout(\eeprom.n2251 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_158_13_lut_LC_18_18_3 .C_ON=1'b1;
    defparam \eeprom.add_158_13_lut_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_158_13_lut_LC_18_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_158_13_lut_LC_18_18_3  (
            .in0(_gnd_net_),
            .in1(N__3539),
            .in2(N__4668),
            .in3(N__3282),
            .lcout(\eeprom.delay_counter_15_N_171_11 ),
            .ltout(),
            .carryin(\eeprom.n2251 ),
            .carryout(\eeprom.n2252 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_158_14_lut_LC_18_18_4 .C_ON=1'b1;
    defparam \eeprom.add_158_14_lut_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_158_14_lut_LC_18_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_158_14_lut_LC_18_18_4  (
            .in0(_gnd_net_),
            .in1(N__3279),
            .in2(N__3554),
            .in3(N__3255),
            .lcout(\eeprom.delay_counter_15_N_171_12 ),
            .ltout(),
            .carryin(\eeprom.n2252 ),
            .carryout(\eeprom.n2253 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_158_15_lut_LC_18_18_5 .C_ON=1'b1;
    defparam \eeprom.add_158_15_lut_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_158_15_lut_LC_18_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_158_15_lut_LC_18_18_5  (
            .in0(_gnd_net_),
            .in1(N__3543),
            .in2(N__4293),
            .in3(N__3252),
            .lcout(\eeprom.delay_counter_15_N_171_13 ),
            .ltout(),
            .carryin(\eeprom.n2253 ),
            .carryout(\eeprom.n2254 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_158_16_lut_LC_18_18_6 .C_ON=1'b1;
    defparam \eeprom.add_158_16_lut_LC_18_18_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_158_16_lut_LC_18_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.add_158_16_lut_LC_18_18_6  (
            .in0(_gnd_net_),
            .in1(N__4563),
            .in2(N__3555),
            .in3(N__3558),
            .lcout(\eeprom.delay_counter_15_N_171_14 ),
            .ltout(),
            .carryin(\eeprom.n2254 ),
            .carryout(\eeprom.n2255 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.add_158_17_lut_LC_18_18_7 .C_ON=1'b0;
    defparam \eeprom.add_158_17_lut_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.add_158_17_lut_LC_18_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \eeprom.add_158_17_lut_LC_18_18_7  (
            .in0(N__4584),
            .in1(N__3547),
            .in2(_gnd_net_),
            .in3(N__3477),
            .lcout(\eeprom.delay_counter_15_N_171_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i5_4_lut_adj_15_LC_18_19_0 .C_ON=1'b0;
    defparam \eeprom.i5_4_lut_adj_15_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i5_4_lut_adj_15_LC_18_19_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i5_4_lut_adj_15_LC_18_19_0  (
            .in0(N__3418),
            .in1(N__3391),
            .in2(N__3372),
            .in3(N__3625),
            .lcout(),
            .ltout(\eeprom.n13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1_3_lut_LC_18_19_1 .C_ON=1'b0;
    defparam \eeprom.i1_3_lut_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1_3_lut_LC_18_19_1 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \eeprom.i1_3_lut_LC_18_19_1  (
            .in0(_gnd_net_),
            .in1(N__3474),
            .in2(N__3468),
            .in3(N__4288),
            .lcout(),
            .ltout(\eeprom.n7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i5_4_lut_LC_18_19_2 .C_ON=1'b0;
    defparam \eeprom.i5_4_lut_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i5_4_lut_LC_18_19_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i5_4_lut_LC_18_19_2  (
            .in0(N__3448),
            .in1(N__4704),
            .in2(N__3465),
            .in3(N__4596),
            .lcout(\eeprom.n1500 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_i0_i1_LC_18_19_3 .C_ON=1'b0;
    defparam \eeprom.delay_counter_i0_i1_LC_18_19_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i1_LC_18_19_3 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \eeprom.delay_counter_i0_i1_LC_18_19_3  (
            .in0(N__3462),
            .in1(N__4356),
            .in2(N__4544),
            .in3(N__3449),
            .lcout(\eeprom.delay_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5124),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_i0_i0_LC_18_19_4 .C_ON=1'b0;
    defparam \eeprom.delay_counter_i0_i0_LC_18_19_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i0_LC_18_19_4 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \eeprom.delay_counter_i0_i0_LC_18_19_4  (
            .in0(N__3419),
            .in1(N__4517),
            .in2(N__4372),
            .in3(N__3435),
            .lcout(\eeprom.delay_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5124),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_i0_i5_LC_18_19_5 .C_ON=1'b0;
    defparam \eeprom.delay_counter_i0_i5_LC_18_19_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i5_LC_18_19_5 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \eeprom.delay_counter_i0_i5_LC_18_19_5  (
            .in0(N__3392),
            .in1(N__4358),
            .in2(N__4546),
            .in3(N__3405),
            .lcout(\eeprom.delay_counter_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5124),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_i0_i10_LC_18_19_6 .C_ON=1'b0;
    defparam \eeprom.delay_counter_i0_i10_LC_18_19_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i10_LC_18_19_6 .LUT_INIT=16'b1111101000111010;
    LogicCell40 \eeprom.delay_counter_i0_i10_LC_18_19_6  (
            .in0(N__3370),
            .in1(N__4518),
            .in2(N__4373),
            .in3(N__3378),
            .lcout(\eeprom.delay_counter_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5124),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_i0_i4_LC_18_19_7 .C_ON=1'b0;
    defparam \eeprom.delay_counter_i0_i4_LC_18_19_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i4_LC_18_19_7 .LUT_INIT=16'b1110111000101110;
    LogicCell40 \eeprom.delay_counter_i0_i4_LC_18_19_7  (
            .in0(N__3626),
            .in1(N__4357),
            .in2(N__4545),
            .in3(N__3642),
            .lcout(\eeprom.delay_counter_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5124),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i1682_2_lut_3_lut_LC_18_20_0 .C_ON=1'b0;
    defparam \eeprom.i1682_2_lut_3_lut_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i1682_2_lut_3_lut_LC_18_20_0 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \eeprom.i1682_2_lut_3_lut_LC_18_20_0  (
            .in0(N__4469),
            .in1(N__5929),
            .in2(_gnd_net_),
            .in3(N__3947),
            .lcout(\eeprom.n2453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.data_ready_42_LC_18_20_1 .C_ON=1'b0;
    defparam \eeprom.data_ready_42_LC_18_20_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.data_ready_42_LC_18_20_1 .LUT_INIT=16'b1110111000000010;
    LogicCell40 \eeprom.data_ready_42_LC_18_20_1  (
            .in0(N__3949),
            .in1(N__4471),
            .in2(N__5944),
            .in3(N__3612),
            .lcout(n324),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5128),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_2_lut_adj_10_LC_18_20_2 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_2_lut_adj_10_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_2_lut_adj_10_LC_18_20_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \eeprom.i2c.i1_2_lut_adj_10_LC_18_20_2  (
            .in0(N__5877),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5661),
            .lcout(n41),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i525_3_lut_LC_18_20_3 .C_ON=1'b0;
    defparam \eeprom.i525_3_lut_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i525_3_lut_LC_18_20_3 .LUT_INIT=16'b1010100010101000;
    LogicCell40 \eeprom.i525_3_lut_LC_18_20_3  (
            .in0(N__3948),
            .in1(N__4468),
            .in2(N__5945),
            .in3(_gnd_net_),
            .lcout(\eeprom.n1018 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2_2_lut_adj_14_LC_18_20_4 .C_ON=1'b0;
    defparam \eeprom.i2_2_lut_adj_14_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2_2_lut_adj_14_LC_18_20_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \eeprom.i2_2_lut_adj_14_LC_18_20_4  (
            .in0(_gnd_net_),
            .in1(N__3605),
            .in2(_gnd_net_),
            .in3(N__5550),
            .lcout(),
            .ltout(n6_adj_405_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1566_4_lut_LC_18_20_5.C_ON=1'b0;
    defparam i1566_4_lut_LC_18_20_5.SEQ_MODE=4'b0000;
    defparam i1566_4_lut_LC_18_20_5.LUT_INIT=16'b1100110011001000;
    LogicCell40 i1566_4_lut_LC_18_20_5 (
            .in0(N__5777),
            .in1(N__4467),
            .in2(N__3585),
            .in3(N__3582),
            .lcout(),
            .ltout(n2483_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2_4_lut_LC_18_20_6 .C_ON=1'b0;
    defparam \eeprom.i2_4_lut_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2_4_lut_LC_18_20_6 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \eeprom.i2_4_lut_LC_18_20_6  (
            .in0(N__4218),
            .in1(N__3576),
            .in2(N__3570),
            .in3(N__3567),
            .lcout(n1568),
            .ltout(n1568_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.state__i1_LC_18_20_7 .C_ON=1'b0;
    defparam \eeprom.state__i1_LC_18_20_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.state__i1_LC_18_20_7 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \eeprom.state__i1_LC_18_20_7  (
            .in0(N__3950),
            .in1(N__4470),
            .in2(N__3561),
            .in3(_gnd_net_),
            .lcout(state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5128),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.state__i0_LC_18_21_0 .C_ON=1'b0;
    defparam \eeprom.state__i0_LC_18_21_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.state__i0_LC_18_21_0 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \eeprom.state__i0_LC_18_21_0  (
            .in0(N__5947),
            .in1(N__3953),
            .in2(_gnd_net_),
            .in3(N__4516),
            .lcout(state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5131),
            .ce(N__3918),
            .sr(_gnd_net_));
    defparam i7_4_lut_LC_18_22_0.C_ON=1'b0;
    defparam i7_4_lut_LC_18_22_0.SEQ_MODE=4'b0000;
    defparam i7_4_lut_LC_18_22_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i7_4_lut_LC_18_22_0 (
            .in0(N__3908),
            .in1(N__3896),
            .in2(N__3885),
            .in3(N__3869),
            .lcout(n17_adj_406),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_LC_18_22_2.C_ON=1'b0;
    defparam i2_4_lut_LC_18_22_2.SEQ_MODE=4'b0000;
    defparam i2_4_lut_LC_18_22_2.LUT_INIT=16'b1111111011111100;
    LogicCell40 i2_4_lut_LC_18_22_2 (
            .in0(N__3857),
            .in1(N__3845),
            .in2(N__3834),
            .in3(N__4227),
            .lcout(),
            .ltout(n2512_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_LC_18_22_3.C_ON=1'b0;
    defparam i4_4_lut_LC_18_22_3.SEQ_MODE=4'b0000;
    defparam i4_4_lut_LC_18_22_3.LUT_INIT=16'b1111111111101100;
    LogicCell40 i4_4_lut_LC_18_22_3 (
            .in0(N__3818),
            .in1(N__3678),
            .in2(N__3807),
            .in3(N__3803),
            .lcout(),
            .ltout(n2495_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_LC_18_22_4.C_ON=1'b0;
    defparam i3_4_lut_LC_18_22_4.SEQ_MODE=4'b0000;
    defparam i3_4_lut_LC_18_22_4.LUT_INIT=16'b1100110010000000;
    LogicCell40 i3_4_lut_LC_18_22_4 (
            .in0(N__3791),
            .in1(N__3648),
            .in2(N__3780),
            .in3(N__3776),
            .lcout(n8_adj_412),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_LC_18_22_6.C_ON=1'b0;
    defparam i6_4_lut_LC_18_22_6.SEQ_MODE=4'b0000;
    defparam i6_4_lut_LC_18_22_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_LC_18_22_6 (
            .in0(N__3764),
            .in1(N__3752),
            .in2(N__3741),
            .in3(N__3725),
            .lcout(n16_adj_407),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_3_lut_LC_18_23_0.C_ON=1'b0;
    defparam i3_3_lut_LC_18_23_0.SEQ_MODE=4'b0000;
    defparam i3_3_lut_LC_18_23_0.LUT_INIT=16'b1111111111101110;
    LogicCell40 i3_3_lut_LC_18_23_0 (
            .in0(N__3713),
            .in1(N__3701),
            .in2(_gnd_net_),
            .in3(N__3689),
            .lcout(n8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_18_23_1.C_ON=1'b0;
    defparam i1_2_lut_LC_18_23_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_18_23_1.LUT_INIT=16'b1010101000000000;
    LogicCell40 i1_2_lut_LC_18_23_1 (
            .in0(N__3671),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3659),
            .lcout(n6_adj_413),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9_4_lut_LC_18_23_2.C_ON=1'b0;
    defparam i9_4_lut_LC_18_23_2.SEQ_MODE=4'b0000;
    defparam i9_4_lut_LC_18_23_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i9_4_lut_LC_18_23_2 (
            .in0(N__4272),
            .in1(N__4257),
            .in2(N__4251),
            .in3(N__4233),
            .lcout(n2536),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam read_15_LC_18_23_3.C_ON=1'b0;
    defparam read_15_LC_18_23_3.SEQ_MODE=4'b1000;
    defparam read_15_LC_18_23_3.LUT_INIT=16'b0101010101010100;
    LogicCell40 read_15_LC_18_23_3 (
            .in0(N__4137),
            .in1(N__4050),
            .in2(N__3987),
            .in3(N__4143),
            .lcout(read_N),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5136),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_19_LC_18_23_6.C_ON=1'b0;
    defparam i1_4_lut_adj_19_LC_18_23_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_19_LC_18_23_6.LUT_INIT=16'b1110110011001100;
    LogicCell40 i1_4_lut_adj_19_LC_18_23_6 (
            .in0(N__4187),
            .in1(N__4175),
            .in2(N__4164),
            .in3(N__4149),
            .lcout(n9_adj_404),
            .ltout(n9_adj_404_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1011_4_lut_LC_18_23_7.C_ON=1'b0;
    defparam i1011_4_lut_LC_18_23_7.SEQ_MODE=4'b0000;
    defparam i1011_4_lut_LC_18_23_7.LUT_INIT=16'b0101010101010100;
    LogicCell40 i1011_4_lut_LC_18_23_7 (
            .in0(N__4136),
            .in1(N__4049),
            .in2(N__4119),
            .in3(N__3983),
            .lcout(addr_10__N_70),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_LC_18_24_5.C_ON=1'b0;
    defparam i2_2_lut_LC_18_24_5.SEQ_MODE=4'b0000;
    defparam i2_2_lut_LC_18_24_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 i2_2_lut_LC_18_24_5 (
            .in0(_gnd_net_),
            .in1(N__4073),
            .in2(_gnd_net_),
            .in3(N__4061),
            .lcout(n10_adj_403),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_18_LC_18_24_6.C_ON=1'b0;
    defparam i6_4_lut_adj_18_LC_18_24_6.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_18_LC_18_24_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_adj_18_LC_18_24_6 (
            .in0(N__4037),
            .in1(N__4025),
            .in2(N__4014),
            .in3(N__3998),
            .lcout(n14_adj_401),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_i0_i7_LC_19_17_2 .C_ON=1'b0;
    defparam \eeprom.delay_counter_i0_i7_LC_19_17_2 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i7_LC_19_17_2 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \eeprom.delay_counter_i0_i7_LC_19_17_2  (
            .in0(N__4548),
            .in1(N__4408),
            .in2(N__4650),
            .in3(N__3966),
            .lcout(\eeprom.delay_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5119),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_i0_i3_LC_19_17_3 .C_ON=1'b0;
    defparam \eeprom.delay_counter_i0_i3_LC_19_17_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i3_LC_19_17_3 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \eeprom.delay_counter_i0_i3_LC_19_17_3  (
            .in0(N__4547),
            .in1(N__4700),
            .in2(N__4413),
            .in3(N__4710),
            .lcout(\eeprom.delay_counter_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5119),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_i0_i11_LC_19_18_0 .C_ON=1'b0;
    defparam \eeprom.delay_counter_i0_i11_LC_19_18_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i11_LC_19_18_0 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \eeprom.delay_counter_i0_i11_LC_19_18_0  (
            .in0(N__4540),
            .in1(N__4664),
            .in2(N__4410),
            .in3(N__4680),
            .lcout(\eeprom.delay_counter_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5125),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_i0_i9_LC_19_18_1 .C_ON=1'b0;
    defparam \eeprom.delay_counter_i0_i9_LC_19_18_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i9_LC_19_18_1 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \eeprom.delay_counter_i0_i9_LC_19_18_1  (
            .in0(N__4404),
            .in1(N__4543),
            .in2(N__4623),
            .in3(N__4674),
            .lcout(\eeprom.delay_counter_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5125),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2_2_lut_LC_19_18_2 .C_ON=1'b0;
    defparam \eeprom.i2_2_lut_LC_19_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2_2_lut_LC_19_18_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \eeprom.i2_2_lut_LC_19_18_2  (
            .in0(_gnd_net_),
            .in1(N__4561),
            .in2(_gnd_net_),
            .in3(N__4582),
            .lcout(),
            .ltout(\eeprom.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2_4_lut_adj_16_LC_19_18_3 .C_ON=1'b0;
    defparam \eeprom.i2_4_lut_adj_16_LC_19_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2_4_lut_adj_16_LC_19_18_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i2_4_lut_adj_16_LC_19_18_3  (
            .in0(N__4663),
            .in1(N__4642),
            .in2(N__4626),
            .in3(N__4609),
            .lcout(\eeprom.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_i0_i15_LC_19_18_4 .C_ON=1'b0;
    defparam \eeprom.delay_counter_i0_i15_LC_19_18_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i15_LC_19_18_4 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \eeprom.delay_counter_i0_i15_LC_19_18_4  (
            .in0(N__4542),
            .in1(N__4583),
            .in2(N__4412),
            .in3(N__4590),
            .lcout(\eeprom.delay_counter_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5125),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_i0_i14_LC_19_18_6 .C_ON=1'b0;
    defparam \eeprom.delay_counter_i0_i14_LC_19_18_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i14_LC_19_18_6 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \eeprom.delay_counter_i0_i14_LC_19_18_6  (
            .in0(N__4541),
            .in1(N__4569),
            .in2(N__4411),
            .in3(N__4562),
            .lcout(\eeprom.delay_counter_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5125),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i2c_clk_122_LC_19_19_2 .C_ON=1'b0;
    defparam \eeprom.i2c.i2c_clk_122_LC_19_19_2 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.i2c_clk_122_LC_19_19_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \eeprom.i2c.i2c_clk_122_LC_19_19_2  (
            .in0(N__6106),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5066),
            .lcout(\eeprom.i2c.i2c_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5129),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.delay_counter_i0_i13_LC_19_19_7 .C_ON=1'b0;
    defparam \eeprom.delay_counter_i0_i13_LC_19_19_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.delay_counter_i0_i13_LC_19_19_7 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \eeprom.delay_counter_i0_i13_LC_19_19_7  (
            .in0(N__4539),
            .in1(N__4292),
            .in2(N__4409),
            .in3(N__4299),
            .lcout(\eeprom.delay_counter_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5129),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.write_enable_132_LC_19_20_6 .C_ON=1'b0;
    defparam \eeprom.i2c.write_enable_132_LC_19_20_6 .SEQ_MODE=4'b1001;
    defparam \eeprom.i2c.write_enable_132_LC_19_20_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \eeprom.i2c.write_enable_132_LC_19_20_6  (
            .in0(N__4799),
            .in1(N__5761),
            .in2(_gnd_net_),
            .in3(N__5861),
            .lcout(sda_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVeeprom.i2c.write_enable_132C_net ),
            .ce(N__4719),
            .sr(N__4740));
    defparam \eeprom.i2c.i22_3_lut_3_lut_LC_19_21_0 .C_ON=1'b0;
    defparam \eeprom.i2c.i22_3_lut_3_lut_LC_19_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i22_3_lut_3_lut_LC_19_21_0 .LUT_INIT=16'b0101010100100010;
    LogicCell40 \eeprom.i2c.i22_3_lut_3_lut_LC_19_21_0  (
            .in0(N__5517),
            .in1(N__5616),
            .in2(_gnd_net_),
            .in3(N__5726),
            .lcout(\eeprom.i2c.n11_adj_379 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i56_3_lut_LC_19_21_1 .C_ON=1'b0;
    defparam \eeprom.i2c.i56_3_lut_LC_19_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i56_3_lut_LC_19_21_1 .LUT_INIT=16'b0010001001100110;
    LogicCell40 \eeprom.i2c.i56_3_lut_LC_19_21_1  (
            .in0(N__5724),
            .in1(N__5516),
            .in2(_gnd_net_),
            .in3(N__5837),
            .lcout(\eeprom.i2c.n33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_7__I_0_140_i11_2_lut_3_lut_4_lut_LC_19_21_2 .C_ON=1'b0;
    defparam \eeprom.i2c.state_7__I_0_140_i11_2_lut_3_lut_4_lut_LC_19_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.state_7__I_0_140_i11_2_lut_3_lut_4_lut_LC_19_21_2 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \eeprom.i2c.state_7__I_0_140_i11_2_lut_3_lut_4_lut_LC_19_21_2  (
            .in0(N__5840),
            .in1(N__5618),
            .in2(N__5539),
            .in3(N__5727),
            .lcout(n11_adj_399),
            .ltout(n11_adj_399_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1673_2_lut_3_lut_LC_19_21_3.C_ON=1'b0;
    defparam i1673_2_lut_3_lut_LC_19_21_3.SEQ_MODE=4'b0000;
    defparam i1673_2_lut_3_lut_LC_19_21_3.LUT_INIT=16'b1111110011110000;
    LogicCell40 i1673_2_lut_3_lut_LC_19_21_3 (
            .in0(_gnd_net_),
            .in1(N__4924),
            .in2(N__4743),
            .in3(N__4958),
            .lcout(n2569),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_3_lut_adj_9_LC_19_21_4 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_3_lut_adj_9_LC_19_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_3_lut_adj_9_LC_19_21_4 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \eeprom.i2c.i1_3_lut_adj_9_LC_19_21_4  (
            .in0(N__4986),
            .in1(N__5617),
            .in2(_gnd_net_),
            .in3(N__4731),
            .lcout(\eeprom.i2c.n1669 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_4_lut_4_lut_LC_19_21_5 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_4_lut_4_lut_LC_19_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_4_lut_4_lut_LC_19_21_5 .LUT_INIT=16'b0001000100110010;
    LogicCell40 \eeprom.i2c.i1_4_lut_4_lut_LC_19_21_5  (
            .in0(N__5725),
            .in1(N__5515),
            .in2(N__5648),
            .in3(N__5838),
            .lcout(\eeprom.i2c.n37 ),
            .ltout(\eeprom.i2c.n37_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_3_lut_adj_8_LC_19_21_6 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_3_lut_adj_8_LC_19_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_3_lut_adj_8_LC_19_21_6 .LUT_INIT=16'b1111001111110000;
    LogicCell40 \eeprom.i2c.i1_3_lut_adj_8_LC_19_21_6  (
            .in0(_gnd_net_),
            .in1(N__5615),
            .in2(N__4734),
            .in3(N__4730),
            .lcout(\eeprom.i2c.n39 ),
            .ltout(\eeprom.i2c.n39_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1692_4_lut_4_lut_LC_19_21_7 .C_ON=1'b0;
    defparam \eeprom.i2c.i1692_4_lut_4_lut_LC_19_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1692_4_lut_4_lut_LC_19_21_7 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \eeprom.i2c.i1692_4_lut_4_lut_LC_19_21_7  (
            .in0(N__5619),
            .in1(N__4798),
            .in2(N__4722),
            .in3(N__5839),
            .lcout(\eeprom.i2c.n1027 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.sda_out_133_LC_19_22_3 .C_ON=1'b0;
    defparam \eeprom.i2c.sda_out_133_LC_19_22_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.sda_out_133_LC_19_22_3 .LUT_INIT=16'b0000010001010100;
    LogicCell40 \eeprom.i2c.sda_out_133_LC_19_22_3  (
            .in0(N__5874),
            .in1(N__4866),
            .in2(N__4803),
            .in3(N__5768),
            .lcout(sda_out),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVeeprom.i2c.sda_out_133C_net ),
            .ce(N__4998),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_2_lut_LC_20_18_1 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_2_lut_LC_20_18_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_2_lut_LC_20_18_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \eeprom.i2c.i1_2_lut_LC_20_18_1  (
            .in0(_gnd_net_),
            .in1(N__5147),
            .in2(_gnd_net_),
            .in3(N__5195),
            .lcout(),
            .ltout(\eeprom.i2c.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i4_4_lut_LC_20_18_2 .C_ON=1'b0;
    defparam \eeprom.i2c.i4_4_lut_LC_20_18_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i4_4_lut_LC_20_18_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \eeprom.i2c.i4_4_lut_LC_20_18_2  (
            .in0(N__5210),
            .in1(N__5180),
            .in2(N__4782),
            .in3(N__5165),
            .lcout(\eeprom.i2c.counter2_7__N_256 ),
            .ltout(\eeprom.i2c.counter2_7__N_256_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_2_lut_3_lut_adj_11_LC_20_18_3 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_2_lut_3_lut_adj_11_LC_20_18_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_2_lut_3_lut_adj_11_LC_20_18_3 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \eeprom.i2c.i1_2_lut_3_lut_adj_11_LC_20_18_3  (
            .in0(_gnd_net_),
            .in1(N__6117),
            .in2(N__4779),
            .in3(N__4849),
            .lcout(\eeprom.i2c.n1580 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.enable_slow_121_LC_20_19_6 .C_ON=1'b0;
    defparam \eeprom.i2c.enable_slow_121_LC_20_19_6 .SEQ_MODE=4'b1001;
    defparam \eeprom.i2c.enable_slow_121_LC_20_19_6 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \eeprom.i2c.enable_slow_121_LC_20_19_6  (
            .in0(N__6110),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5065),
            .lcout(state_7_N_269_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5132),
            .ce(N__4776),
            .sr(N__4856));
    defparam \eeprom.i2c.state_i0_i0_LC_20_20_0 .C_ON=1'b0;
    defparam \eeprom.i2c.state_i0_i0_LC_20_20_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.state_i0_i0_LC_20_20_0 .LUT_INIT=16'b1010101000111111;
    LogicCell40 \eeprom.i2c.state_i0_i0_LC_20_20_0  (
            .in0(N__5776),
            .in1(N__5250),
            .in2(N__5457),
            .in3(N__4884),
            .lcout(state_0_adj_397),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6130),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.saved_addr__i1_LC_20_20_1 .C_ON=1'b0;
    defparam \eeprom.i2c.saved_addr__i1_LC_20_20_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.saved_addr__i1_LC_20_20_1 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \eeprom.i2c.saved_addr__i1_LC_20_20_1  (
            .in0(N__5909),
            .in1(N__5264),
            .in2(N__4770),
            .in3(N__5040),
            .lcout(saved_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6130),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1004_2_lut_3_lut_LC_20_20_3 .C_ON=1'b0;
    defparam \eeprom.i2c.i1004_2_lut_3_lut_LC_20_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1004_2_lut_3_lut_LC_20_20_3 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \eeprom.i2c.i1004_2_lut_3_lut_LC_20_20_3  (
            .in0(N__5637),
            .in1(N__5772),
            .in2(_gnd_net_),
            .in3(N__5857),
            .lcout(n1835),
            .ltout(n1835_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_3_lut_LC_20_20_4 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_3_lut_LC_20_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_3_lut_LC_20_20_4 .LUT_INIT=16'b1111101010101010;
    LogicCell40 \eeprom.i2c.i1_3_lut_LC_20_20_4  (
            .in0(N__5354),
            .in1(_gnd_net_),
            .in2(N__4752),
            .in3(N__5537),
            .lcout(n949),
            .ltout(n949_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_i0_i2_LC_20_20_5 .C_ON=1'b0;
    defparam \eeprom.i2c.state_i0_i2_LC_20_20_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.state_i0_i2_LC_20_20_5 .LUT_INIT=16'b1111011100000111;
    LogicCell40 \eeprom.i2c.state_i0_i2_LC_20_20_5  (
            .in0(N__5456),
            .in1(N__4749),
            .in2(N__4887),
            .in3(N__5859),
            .lcout(state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6130),
            .ce(),
            .sr(_gnd_net_));
    defparam i1630_4_lut_4_lut_LC_20_20_6.C_ON=1'b0;
    defparam i1630_4_lut_4_lut_LC_20_20_6.SEQ_MODE=4'b0000;
    defparam i1630_4_lut_4_lut_LC_20_20_6.LUT_INIT=16'b1110111111001011;
    LogicCell40 i1630_4_lut_4_lut_LC_20_20_6 (
            .in0(N__5858),
            .in1(N__5638),
            .in2(N__5778),
            .in3(N__5538),
            .lcout(),
            .ltout(n2547_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_i0_i1_LC_20_20_7 .C_ON=1'b0;
    defparam \eeprom.i2c.state_i0_i1_LC_20_20_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.state_i0_i1_LC_20_20_7 .LUT_INIT=16'b1011101110001011;
    LogicCell40 \eeprom.i2c.state_i0_i1_LC_20_20_7  (
            .in0(N__5639),
            .in1(N__4883),
            .in2(N__4872),
            .in3(N__5010),
            .lcout(state_1_adj_396),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6130),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1667_2_lut_LC_20_21_0 .C_ON=1'b0;
    defparam \eeprom.i2c.i1667_2_lut_LC_20_21_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1667_2_lut_LC_20_21_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \eeprom.i2c.i1667_2_lut_LC_20_21_0  (
            .in0(_gnd_net_),
            .in1(N__5038),
            .in2(_gnd_net_),
            .in3(N__6379),
            .lcout(),
            .ltout(\eeprom.i2c.n2574_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1666_4_lut_LC_20_21_1 .C_ON=1'b0;
    defparam \eeprom.i2c.i1666_4_lut_LC_20_21_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1666_4_lut_LC_20_21_1 .LUT_INIT=16'b1001100000000000;
    LogicCell40 \eeprom.i2c.i1666_4_lut_LC_20_21_1  (
            .in0(N__6347),
            .in1(N__5335),
            .in2(N__4869),
            .in3(N__5623),
            .lcout(\eeprom.i2c.n2557 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i2_4_lut_4_lut_LC_20_21_2 .C_ON=1'b0;
    defparam \eeprom.i2c.i2_4_lut_4_lut_LC_20_21_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i2_4_lut_4_lut_LC_20_21_2 .LUT_INIT=16'b1101110101011101;
    LogicCell40 \eeprom.i2c.i2_4_lut_4_lut_LC_20_21_2  (
            .in0(N__5624),
            .in1(N__5758),
            .in2(N__4860),
            .in3(N__6245),
            .lcout(),
            .ltout(n2538_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_20_21_3.C_ON=1'b0;
    defparam i1_4_lut_LC_20_21_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_20_21_3.LUT_INIT=16'b0010001011110010;
    LogicCell40 i1_4_lut_LC_20_21_3 (
            .in0(N__6246),
            .in1(N__5021),
            .in2(N__4824),
            .in3(N__5392),
            .lcout(),
            .ltout(n4_adj_411_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_LC_20_21_4.C_ON=1'b0;
    defparam i2_3_lut_4_lut_LC_20_21_4.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_LC_20_21_4.LUT_INIT=16'b1111000011110010;
    LogicCell40 i2_3_lut_4_lut_LC_20_21_4 (
            .in0(N__5625),
            .in1(N__4809),
            .in2(N__4821),
            .in3(N__5759),
            .lcout(),
            .ltout(n2507_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_i0_i3_LC_20_21_5 .C_ON=1'b0;
    defparam \eeprom.i2c.state_i0_i3_LC_20_21_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.state_i0_i3_LC_20_21_5 .LUT_INIT=16'b1010101011111000;
    LogicCell40 \eeprom.i2c.state_i0_i3_LC_20_21_5  (
            .in0(N__5536),
            .in1(N__4818),
            .in2(N__4812),
            .in3(N__5355),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6170),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_7__I_0_142_i10_2_lut_LC_20_21_6 .C_ON=1'b0;
    defparam \eeprom.i2c.state_7__I_0_142_i10_2_lut_LC_20_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.state_7__I_0_142_i10_2_lut_LC_20_21_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \eeprom.i2c.state_7__I_0_142_i10_2_lut_LC_20_21_6  (
            .in0(_gnd_net_),
            .in1(N__5535),
            .in2(_gnd_net_),
            .in3(N__5860),
            .lcout(n10_adj_394),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1674_3_lut_4_lut_LC_20_21_7.C_ON=1'b0;
    defparam i1674_3_lut_4_lut_LC_20_21_7.SEQ_MODE=4'b0000;
    defparam i1674_3_lut_4_lut_LC_20_21_7.LUT_INIT=16'b0000001000001010;
    LogicCell40 i1674_3_lut_4_lut_LC_20_21_7 (
            .in0(N__5039),
            .in1(N__4923),
            .in2(N__5025),
            .in3(N__4959),
            .lcout(n2566),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1686_4_lut_LC_20_22_0 .C_ON=1'b0;
    defparam \eeprom.i2c.i1686_4_lut_LC_20_22_0 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1686_4_lut_LC_20_22_0 .LUT_INIT=16'b0100010001001100;
    LogicCell40 \eeprom.i2c.i1686_4_lut_LC_20_22_0  (
            .in0(N__5651),
            .in1(N__5004),
            .in2(N__4968),
            .in3(N__5870),
            .lcout(\eeprom.i2c.n2406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_2_lut_3_lut_LC_20_22_1 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_2_lut_3_lut_LC_20_22_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_2_lut_3_lut_LC_20_22_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \eeprom.i2c.i1_2_lut_3_lut_LC_20_22_1  (
            .in0(N__5872),
            .in1(N__5767),
            .in2(_gnd_net_),
            .in3(N__5523),
            .lcout(),
            .ltout(\eeprom.i2c.n1051_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i17_4_lut_LC_20_22_2 .C_ON=1'b0;
    defparam \eeprom.i2c.i17_4_lut_LC_20_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i17_4_lut_LC_20_22_2 .LUT_INIT=16'b0000100011111000;
    LogicCell40 \eeprom.i2c.i17_4_lut_LC_20_22_2  (
            .in0(N__4985),
            .in1(N__5403),
            .in2(N__4971),
            .in3(N__4896),
            .lcout(\eeprom.i2c.n1548 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_3_lut_2_lut_LC_20_22_3 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_3_lut_2_lut_LC_20_22_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_3_lut_2_lut_LC_20_22_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \eeprom.i2c.i1_3_lut_2_lut_LC_20_22_3  (
            .in0(_gnd_net_),
            .in1(N__5765),
            .in2(_gnd_net_),
            .in3(N__5521),
            .lcout(\eeprom.i2c.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i463_2_lut_LC_20_22_4 .C_ON=1'b0;
    defparam \eeprom.i2c.i463_2_lut_LC_20_22_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i463_2_lut_LC_20_22_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \eeprom.i2c.i463_2_lut_LC_20_22_4  (
            .in0(_gnd_net_),
            .in1(N__4957),
            .in2(_gnd_net_),
            .in3(N__4928),
            .lcout(state_7_N_285_3),
            .ltout(state_7_N_285_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1558_3_lut_4_lut_LC_20_22_5 .C_ON=1'b0;
    defparam \eeprom.i2c.i1558_3_lut_4_lut_LC_20_22_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1558_3_lut_4_lut_LC_20_22_5 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \eeprom.i2c.i1558_3_lut_4_lut_LC_20_22_5  (
            .in0(N__5871),
            .in1(N__5217),
            .in2(N__4899),
            .in3(N__5522),
            .lcout(\eeprom.i2c.n2475 ),
            .ltout(\eeprom.i2c.n2475_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1545_2_lut_4_lut_LC_20_22_6 .C_ON=1'b0;
    defparam \eeprom.i2c.i1545_2_lut_4_lut_LC_20_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1545_2_lut_4_lut_LC_20_22_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \eeprom.i2c.i1545_2_lut_4_lut_LC_20_22_6  (
            .in0(N__5524),
            .in1(N__5769),
            .in2(N__4890),
            .in3(N__5873),
            .lcout(\eeprom.i2c.n1655 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_7__I_0_142_i9_2_lut_LC_20_22_7 .C_ON=1'b0;
    defparam \eeprom.i2c.state_7__I_0_142_i9_2_lut_LC_20_22_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.state_7__I_0_142_i9_2_lut_LC_20_22_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \eeprom.i2c.state_7__I_0_142_i9_2_lut_LC_20_22_7  (
            .in0(_gnd_net_),
            .in1(N__5766),
            .in2(_gnd_net_),
            .in3(N__5652),
            .lcout(\eeprom.i2c.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.counter2_364_365__i1_LC_21_18_0 .C_ON=1'b1;
    defparam \eeprom.i2c.counter2_364_365__i1_LC_21_18_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter2_364_365__i1_LC_21_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter2_364_365__i1_LC_21_18_0  (
            .in0(_gnd_net_),
            .in1(N__5211),
            .in2(_gnd_net_),
            .in3(N__5199),
            .lcout(\eeprom.i2c.counter2_0 ),
            .ltout(),
            .carryin(bfn_21_18_0_),
            .carryout(\eeprom.i2c.n2319 ),
            .clk(N__5133),
            .ce(),
            .sr(N__5070));
    defparam \eeprom.i2c.counter2_364_365__i2_LC_21_18_1 .C_ON=1'b1;
    defparam \eeprom.i2c.counter2_364_365__i2_LC_21_18_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter2_364_365__i2_LC_21_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter2_364_365__i2_LC_21_18_1  (
            .in0(_gnd_net_),
            .in1(N__5196),
            .in2(_gnd_net_),
            .in3(N__5184),
            .lcout(\eeprom.i2c.counter2_1 ),
            .ltout(),
            .carryin(\eeprom.i2c.n2319 ),
            .carryout(\eeprom.i2c.n2320 ),
            .clk(N__5133),
            .ce(),
            .sr(N__5070));
    defparam \eeprom.i2c.counter2_364_365__i3_LC_21_18_2 .C_ON=1'b1;
    defparam \eeprom.i2c.counter2_364_365__i3_LC_21_18_2 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter2_364_365__i3_LC_21_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter2_364_365__i3_LC_21_18_2  (
            .in0(_gnd_net_),
            .in1(N__5181),
            .in2(_gnd_net_),
            .in3(N__5169),
            .lcout(\eeprom.i2c.counter2_2 ),
            .ltout(),
            .carryin(\eeprom.i2c.n2320 ),
            .carryout(\eeprom.i2c.n2321 ),
            .clk(N__5133),
            .ce(),
            .sr(N__5070));
    defparam \eeprom.i2c.counter2_364_365__i4_LC_21_18_3 .C_ON=1'b1;
    defparam \eeprom.i2c.counter2_364_365__i4_LC_21_18_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter2_364_365__i4_LC_21_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter2_364_365__i4_LC_21_18_3  (
            .in0(_gnd_net_),
            .in1(N__5166),
            .in2(_gnd_net_),
            .in3(N__5154),
            .lcout(\eeprom.i2c.counter2_3 ),
            .ltout(),
            .carryin(\eeprom.i2c.n2321 ),
            .carryout(\eeprom.i2c.n2322 ),
            .clk(N__5133),
            .ce(),
            .sr(N__5070));
    defparam \eeprom.i2c.counter2_364_365__i5_LC_21_18_4 .C_ON=1'b0;
    defparam \eeprom.i2c.counter2_364_365__i5_LC_21_18_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter2_364_365__i5_LC_21_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter2_364_365__i5_LC_21_18_4  (
            .in0(_gnd_net_),
            .in1(N__5148),
            .in2(_gnd_net_),
            .in3(N__5151),
            .lcout(\eeprom.i2c.counter2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5133),
            .ce(),
            .sr(N__5070));
    defparam \eeprom.i2c.data_out_i0_i7_LC_21_20_0 .C_ON=1'b0;
    defparam \eeprom.i2c.data_out_i0_i7_LC_21_20_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.data_out_i0_i7_LC_21_20_0 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \eeprom.i2c.data_out_i0_i7_LC_21_20_0  (
            .in0(N__5430),
            .in1(N__6424),
            .in2(N__5049),
            .in3(N__6269),
            .lcout(n306),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6165),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.equal_25_i11_2_lut_3_lut_4_lut_LC_21_20_1 .C_ON=1'b0;
    defparam \eeprom.i2c.equal_25_i11_2_lut_3_lut_4_lut_LC_21_20_1 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.equal_25_i11_2_lut_3_lut_4_lut_LC_21_20_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i2c.equal_25_i11_2_lut_3_lut_4_lut_LC_21_20_1  (
            .in0(N__5741),
            .in1(N__5525),
            .in2(N__5649),
            .in3(N__5841),
            .lcout(n15_adj_393),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_7__I_0_139_i11_2_lut_4_lut_LC_21_20_2 .C_ON=1'b0;
    defparam \eeprom.i2c.state_7__I_0_139_i11_2_lut_4_lut_LC_21_20_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.state_7__I_0_139_i11_2_lut_4_lut_LC_21_20_2 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \eeprom.i2c.state_7__I_0_139_i11_2_lut_4_lut_LC_21_20_2  (
            .in0(N__5843),
            .in1(N__5742),
            .in2(N__5650),
            .in3(N__5533),
            .lcout(n11_adj_400),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_2_lut_3_lut_4_lut_adj_12_LC_21_20_3 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_2_lut_3_lut_4_lut_adj_12_LC_21_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_2_lut_3_lut_4_lut_adj_12_LC_21_20_3 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \eeprom.i2c.i1_2_lut_3_lut_4_lut_adj_12_LC_21_20_3  (
            .in0(N__5745),
            .in1(N__5343),
            .in2(N__5397),
            .in3(N__5631),
            .lcout(n1518),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.state_7__I_0_143_i10_2_lut_LC_21_20_4 .C_ON=1'b0;
    defparam \eeprom.i2c.state_7__I_0_143_i10_2_lut_LC_21_20_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.state_7__I_0_143_i10_2_lut_LC_21_20_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \eeprom.i2c.state_7__I_0_143_i10_2_lut_LC_21_20_4  (
            .in0(N__5842),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5532),
            .lcout(n10_adj_398),
            .ltout(n10_adj_398_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_2_lut_3_lut_4_lut_LC_21_20_5 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_2_lut_3_lut_4_lut_LC_21_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_2_lut_3_lut_4_lut_LC_21_20_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \eeprom.i2c.i1_2_lut_3_lut_4_lut_LC_21_20_5  (
            .in0(N__5744),
            .in1(N__5342),
            .in2(N__5268),
            .in3(N__5630),
            .lcout(n1523),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_3_lut_LC_21_20_6.C_ON=1'b0;
    defparam i1_3_lut_3_lut_LC_21_20_6.SEQ_MODE=4'b0000;
    defparam i1_3_lut_3_lut_LC_21_20_6.LUT_INIT=16'b1111111100010001;
    LogicCell40 i1_3_lut_3_lut_LC_21_20_6 (
            .in0(N__5844),
            .in1(N__5265),
            .in2(_gnd_net_),
            .in3(N__5534),
            .lcout(),
            .ltout(n2460_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1676_4_lut_LC_21_20_7.C_ON=1'b0;
    defparam i1676_4_lut_LC_21_20_7.SEQ_MODE=4'b0000;
    defparam i1676_4_lut_LC_21_20_7.LUT_INIT=16'b1100110011001000;
    LogicCell40 i1676_4_lut_LC_21_20_7 (
            .in0(N__5743),
            .in1(N__5372),
            .in2(N__5253),
            .in3(N__5629),
            .lcout(n2560),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.data_out_i0_i6_LC_21_21_0 .C_ON=1'b0;
    defparam \eeprom.i2c.data_out_i0_i6_LC_21_21_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.data_out_i0_i6_LC_21_21_0 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \eeprom.i2c.data_out_i0_i6_LC_21_21_0  (
            .in0(N__6258),
            .in1(N__5241),
            .in2(N__6312),
            .in3(N__5429),
            .lcout(n308),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6180),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.data_out_i0_i0_LC_21_21_1 .C_ON=1'b0;
    defparam \eeprom.i2c.data_out_i0_i0_LC_21_21_1 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.data_out_i0_i0_LC_21_21_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \eeprom.i2c.data_out_i0_i0_LC_21_21_1  (
            .in0(N__5414),
            .in1(N__6306),
            .in2(N__5235),
            .in3(N__6256),
            .lcout(n320),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6180),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.data_out_i0_i1_LC_21_21_2 .C_ON=1'b0;
    defparam \eeprom.i2c.data_out_i0_i1_LC_21_21_2 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.data_out_i0_i1_LC_21_21_2 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \eeprom.i2c.data_out_i0_i1_LC_21_21_2  (
            .in0(N__6257),
            .in1(N__6433),
            .in2(N__5226),
            .in3(N__5415),
            .lcout(n318),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6180),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.equal_50_i4_2_lut_LC_21_21_3 .C_ON=1'b0;
    defparam \eeprom.i2c.equal_50_i4_2_lut_LC_21_21_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.equal_50_i4_2_lut_LC_21_21_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \eeprom.i2c.equal_50_i4_2_lut_LC_21_21_3  (
            .in0(_gnd_net_),
            .in1(N__6346),
            .in2(_gnd_net_),
            .in3(N__6380),
            .lcout(n4_adj_408),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i986_2_lut_LC_21_21_4 .C_ON=1'b0;
    defparam \eeprom.i2c.i986_2_lut_LC_21_21_4 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i986_2_lut_LC_21_21_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \eeprom.i2c.i986_2_lut_LC_21_21_4  (
            .in0(N__6381),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6348),
            .lcout(n1817),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i5_4_lut_LC_21_21_5 .C_ON=1'b0;
    defparam \eeprom.i2c.i5_4_lut_LC_21_21_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i5_4_lut_LC_21_21_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i2c.i5_4_lut_LC_21_21_5  (
            .in0(N__5334),
            .in1(N__6050),
            .in2(N__5288),
            .in3(N__5303),
            .lcout(),
            .ltout(\eeprom.i2c.n12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i6_4_lut_LC_21_21_6 .C_ON=1'b0;
    defparam \eeprom.i2c.i6_4_lut_LC_21_21_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i6_4_lut_LC_21_21_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \eeprom.i2c.i6_4_lut_LC_21_21_6  (
            .in0(N__6014),
            .in1(N__6032),
            .in2(N__5418),
            .in3(N__5413),
            .lcout(\eeprom.i2c.n942 ),
            .ltout(\eeprom.i2c.n942_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i1_4_lut_LC_21_21_7 .C_ON=1'b0;
    defparam \eeprom.i2c.i1_4_lut_LC_21_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i1_4_lut_LC_21_21_7 .LUT_INIT=16'b0011000001110000;
    LogicCell40 \eeprom.i2c.i1_4_lut_LC_21_21_7  (
            .in0(N__5396),
            .in1(N__5373),
            .in2(N__5358),
            .in3(N__5760),
            .lcout(n1532),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.counter_i0_LC_21_22_0 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i0_LC_21_22_0 .SEQ_MODE=4'b1001;
    defparam \eeprom.i2c.counter_i0_LC_21_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i0_LC_21_22_0  (
            .in0(_gnd_net_),
            .in1(N__5336),
            .in2(_gnd_net_),
            .in3(N__5313),
            .lcout(\eeprom.i2c.counter_0 ),
            .ltout(),
            .carryin(bfn_21_22_0_),
            .carryout(\eeprom.i2c.n2256 ),
            .clk(N__6169),
            .ce(N__6003),
            .sr(N__5997));
    defparam \eeprom.i2c.counter_i1_LC_21_22_1 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i1_LC_21_22_1 .SEQ_MODE=4'b1001;
    defparam \eeprom.i2c.counter_i1_LC_21_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i1_LC_21_22_1  (
            .in0(_gnd_net_),
            .in1(N__6382),
            .in2(N__5986),
            .in3(N__5310),
            .lcout(\eeprom.i2c.counter_1 ),
            .ltout(),
            .carryin(\eeprom.i2c.n2256 ),
            .carryout(\eeprom.i2c.n2257 ),
            .clk(N__6169),
            .ce(N__6003),
            .sr(N__5997));
    defparam \eeprom.i2c.counter_i2_LC_21_22_2 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i2_LC_21_22_2 .SEQ_MODE=4'b1001;
    defparam \eeprom.i2c.counter_i2_LC_21_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i2_LC_21_22_2  (
            .in0(_gnd_net_),
            .in1(N__5976),
            .in2(N__6354),
            .in3(N__5307),
            .lcout(\eeprom.i2c.counter_2 ),
            .ltout(),
            .carryin(\eeprom.i2c.n2257 ),
            .carryout(\eeprom.i2c.n2258 ),
            .clk(N__6169),
            .ce(N__6003),
            .sr(N__5997));
    defparam \eeprom.i2c.counter_i3_LC_21_22_3 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i3_LC_21_22_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter_i3_LC_21_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i3_LC_21_22_3  (
            .in0(_gnd_net_),
            .in1(N__5304),
            .in2(N__5987),
            .in3(N__5292),
            .lcout(\eeprom.i2c.counter_3 ),
            .ltout(),
            .carryin(\eeprom.i2c.n2258 ),
            .carryout(\eeprom.i2c.n2259 ),
            .clk(N__6169),
            .ce(N__6003),
            .sr(N__5997));
    defparam \eeprom.i2c.counter_i4_LC_21_22_4 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i4_LC_21_22_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter_i4_LC_21_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i4_LC_21_22_4  (
            .in0(_gnd_net_),
            .in1(N__5980),
            .in2(N__5289),
            .in3(N__5271),
            .lcout(\eeprom.i2c.counter_4 ),
            .ltout(),
            .carryin(\eeprom.i2c.n2259 ),
            .carryout(\eeprom.i2c.n2260 ),
            .clk(N__6169),
            .ce(N__6003),
            .sr(N__5997));
    defparam \eeprom.i2c.counter_i5_LC_21_22_5 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i5_LC_21_22_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter_i5_LC_21_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i5_LC_21_22_5  (
            .in0(_gnd_net_),
            .in1(N__6051),
            .in2(N__5988),
            .in3(N__6039),
            .lcout(\eeprom.i2c.counter_5 ),
            .ltout(),
            .carryin(\eeprom.i2c.n2260 ),
            .carryout(\eeprom.i2c.n2261 ),
            .clk(N__6169),
            .ce(N__6003),
            .sr(N__5997));
    defparam \eeprom.i2c.counter_i6_LC_21_22_6 .C_ON=1'b1;
    defparam \eeprom.i2c.counter_i6_LC_21_22_6 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter_i6_LC_21_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \eeprom.i2c.counter_i6_LC_21_22_6  (
            .in0(_gnd_net_),
            .in1(N__5984),
            .in2(N__6036),
            .in3(N__6021),
            .lcout(\eeprom.i2c.counter_6 ),
            .ltout(),
            .carryin(\eeprom.i2c.n2261 ),
            .carryout(\eeprom.i2c.n2262 ),
            .clk(N__6169),
            .ce(N__6003),
            .sr(N__5997));
    defparam \eeprom.i2c.counter_i7_LC_21_22_7 .C_ON=1'b0;
    defparam \eeprom.i2c.counter_i7_LC_21_22_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.counter_i7_LC_21_22_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \eeprom.i2c.counter_i7_LC_21_22_7  (
            .in0(N__5985),
            .in1(N__6015),
            .in2(_gnd_net_),
            .in3(N__6018),
            .lcout(\eeprom.i2c.counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6169),
            .ce(N__6003),
            .sr(N__5997));
    defparam CONSTANT_ONE_LUT4_LC_21_24_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_21_24_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_21_24_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_21_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i26_2_lut_LC_22_20_3 .C_ON=1'b0;
    defparam \eeprom.i2c.i26_2_lut_LC_22_20_3 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i26_2_lut_LC_22_20_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \eeprom.i2c.i26_2_lut_LC_22_20_3  (
            .in0(_gnd_net_),
            .in1(N__5770),
            .in2(_gnd_net_),
            .in3(N__5548),
            .lcout(),
            .ltout(\eeprom.i2c.n10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i2c_scl_enable_124_LC_22_20_4 .C_ON=1'b0;
    defparam \eeprom.i2c.i2c_scl_enable_124_LC_22_20_4 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.i2c_scl_enable_124_LC_22_20_4 .LUT_INIT=16'b1010101010001010;
    LogicCell40 \eeprom.i2c.i2c_scl_enable_124_LC_22_20_4  (
            .in0(N__5908),
            .in1(N__5653),
            .in2(N__5880),
            .in3(N__5875),
            .lcout(scl_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVeeprom.i2c.i2c_scl_enable_124C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i995_3_lut_4_lut_4_lut_LC_22_20_5 .C_ON=1'b0;
    defparam \eeprom.i2c.i995_3_lut_4_lut_4_lut_LC_22_20_5 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i995_3_lut_4_lut_4_lut_LC_22_20_5 .LUT_INIT=16'b1111101111011111;
    LogicCell40 \eeprom.i2c.i995_3_lut_4_lut_4_lut_LC_22_20_5  (
            .in0(N__5876),
            .in1(N__5771),
            .in2(N__5660),
            .in3(N__5549),
            .lcout(n1826),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.data_out_i0_i3_LC_22_22_0 .C_ON=1'b0;
    defparam \eeprom.i2c.data_out_i0_i3_LC_22_22_0 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.data_out_i0_i3_LC_22_22_0 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \eeprom.i2c.data_out_i0_i3_LC_22_22_0  (
            .in0(N__6266),
            .in1(N__6318),
            .in2(N__5439),
            .in3(N__6434),
            .lcout(n314),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6183),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.equal_45_i4_2_lut_LC_22_22_2 .C_ON=1'b0;
    defparam \eeprom.i2c.equal_45_i4_2_lut_LC_22_22_2 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.equal_45_i4_2_lut_LC_22_22_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \eeprom.i2c.equal_45_i4_2_lut_LC_22_22_2  (
            .in0(_gnd_net_),
            .in1(N__6383),
            .in2(_gnd_net_),
            .in3(N__6352),
            .lcout(n4_adj_395),
            .ltout(n4_adj_395_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.data_out_i0_i5_LC_22_22_3 .C_ON=1'b0;
    defparam \eeprom.i2c.data_out_i0_i5_LC_22_22_3 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.data_out_i0_i5_LC_22_22_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \eeprom.i2c.data_out_i0_i5_LC_22_22_3  (
            .in0(N__6435),
            .in1(N__6405),
            .in2(N__6408),
            .in3(N__6268),
            .lcout(n310),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6183),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.data_out_i0_i4_LC_22_22_5 .C_ON=1'b0;
    defparam \eeprom.i2c.data_out_i0_i4_LC_22_22_5 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.data_out_i0_i4_LC_22_22_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \eeprom.i2c.data_out_i0_i4_LC_22_22_5  (
            .in0(N__6399),
            .in1(N__6311),
            .in2(N__6393),
            .in3(N__6267),
            .lcout(n312),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6183),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.equal_48_i4_2_lut_LC_22_22_6 .C_ON=1'b0;
    defparam \eeprom.i2c.equal_48_i4_2_lut_LC_22_22_6 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.equal_48_i4_2_lut_LC_22_22_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \eeprom.i2c.equal_48_i4_2_lut_LC_22_22_6  (
            .in0(_gnd_net_),
            .in1(N__6384),
            .in2(_gnd_net_),
            .in3(N__6353),
            .lcout(n4),
            .ltout(n4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.data_out_i0_i2_LC_22_22_7 .C_ON=1'b0;
    defparam \eeprom.i2c.data_out_i0_i2_LC_22_22_7 .SEQ_MODE=4'b1000;
    defparam \eeprom.i2c.data_out_i0_i2_LC_22_22_7 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \eeprom.i2c.data_out_i0_i2_LC_22_22_7  (
            .in0(N__6213),
            .in1(N__6310),
            .in2(N__6285),
            .in3(N__6265),
            .lcout(n316),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6183),
            .ce(),
            .sr(_gnd_net_));
    defparam \eeprom.i2c.i989_2_lut_LC_23_21_7 .C_ON=1'b0;
    defparam \eeprom.i2c.i989_2_lut_LC_23_21_7 .SEQ_MODE=4'b0000;
    defparam \eeprom.i2c.i989_2_lut_LC_23_21_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \eeprom.i2c.i989_2_lut_LC_23_21_7  (
            .in0(N__6194),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6182),
            .lcout(scl_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
