-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Jan 30 2020 23:28:46

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    TX : out std_logic;
    SDA : inout std_logic;
    SCL : inout std_logic;
    RX : in std_logic;
    NEOPXL : out std_logic;
    LED : out std_logic;
    INLC : out std_logic;
    INLB : out std_logic;
    INLA : out std_logic;
    INHC : out std_logic;
    INHB : out std_logic;
    INHA : out std_logic;
    HALL3 : in std_logic;
    HALL2 : in std_logic;
    HALL1 : in std_logic;
    FAULT_N : in std_logic;
    ENCODER1_B : in std_logic;
    ENCODER1_A : in std_logic;
    ENCODER0_B : in std_logic;
    ENCODER0_A : in std_logic;
    DE : out std_logic;
    CS_MISO : in std_logic;
    CS_CLK : out std_logic;
    CS : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__6680\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3859\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3433\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3219\ : std_logic;
signal \N__3216\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3201\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3144\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3126\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3087\ : std_logic;
signal \N__3084\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3018\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3009\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2845\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2824\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2809\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2788\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2725\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \n2955_cascade_\ : std_logic;
signal \LED_c\ : std_logic;
signal n2954 : std_logic;
signal \bfn_19_13_0_\ : std_logic;
signal \eeprom.n2671\ : std_logic;
signal \eeprom.n2672\ : std_logic;
signal \eeprom.n2673\ : std_logic;
signal \eeprom.n2674\ : std_logic;
signal \eeprom.n2675\ : std_logic;
signal \eeprom.n2676\ : std_logic;
signal \eeprom.n2677\ : std_logic;
signal \eeprom.n2678\ : std_logic;
signal \bfn_19_14_0_\ : std_logic;
signal \eeprom.n2679\ : std_logic;
signal \eeprom.n2680\ : std_logic;
signal \eeprom.n2681\ : std_logic;
signal \eeprom.n2682\ : std_logic;
signal \eeprom.n2683\ : std_logic;
signal \eeprom.n2684\ : std_logic;
signal \eeprom.n2685\ : std_logic;
signal n26 : std_logic;
signal \bfn_19_17_0_\ : std_logic;
signal n25_adj_407 : std_logic;
signal n2691 : std_logic;
signal n24_adj_406 : std_logic;
signal n2692 : std_logic;
signal n23_adj_405 : std_logic;
signal n2693 : std_logic;
signal n22_adj_404 : std_logic;
signal n2694 : std_logic;
signal n21 : std_logic;
signal n2695 : std_logic;
signal n20_adj_403 : std_logic;
signal n2696 : std_logic;
signal n19 : std_logic;
signal n2697 : std_logic;
signal n2698 : std_logic;
signal n18_adj_402 : std_logic;
signal \bfn_19_18_0_\ : std_logic;
signal n17 : std_logic;
signal n2699 : std_logic;
signal n16 : std_logic;
signal n2700 : std_logic;
signal n15_adj_401 : std_logic;
signal n2701 : std_logic;
signal n14_adj_400 : std_logic;
signal n2702 : std_logic;
signal n13_adj_399 : std_logic;
signal n2703 : std_logic;
signal n12 : std_logic;
signal n2704 : std_logic;
signal n11 : std_logic;
signal n2705 : std_logic;
signal n2706 : std_logic;
signal n10_adj_398 : std_logic;
signal \bfn_19_19_0_\ : std_logic;
signal n9 : std_logic;
signal n2707 : std_logic;
signal n8_adj_397 : std_logic;
signal n2708 : std_logic;
signal n7 : std_logic;
signal n2709 : std_logic;
signal n6_adj_396 : std_logic;
signal n2710 : std_logic;
signal blink_counter_21 : std_logic;
signal n2711 : std_logic;
signal blink_counter_22 : std_logic;
signal n2712 : std_logic;
signal blink_counter_23 : std_logic;
signal n2713 : std_logic;
signal n2714 : std_logic;
signal blink_counter_24 : std_logic;
signal \bfn_19_20_0_\ : std_logic;
signal n2715 : std_logic;
signal blink_counter_25 : std_logic;
signal \eeprom.delay_counter_7\ : std_logic;
signal \eeprom.delay_counter_2\ : std_logic;
signal \eeprom.delay_counter_5\ : std_logic;
signal \eeprom.delay_counter_11\ : std_logic;
signal \eeprom.n1934\ : std_logic;
signal \eeprom.delay_counter_13\ : std_logic;
signal \eeprom.delay_counter_9\ : std_logic;
signal \eeprom.delay_counter_0\ : std_logic;
signal \eeprom.delay_counter_4\ : std_logic;
signal \eeprom.delay_counter_14\ : std_logic;
signal \eeprom.delay_counter_3\ : std_logic;
signal \eeprom.delay_counter_1\ : std_logic;
signal \eeprom.delay_counter_15\ : std_logic;
signal \eeprom.n1799\ : std_logic;
signal \eeprom.delay_counter_12\ : std_logic;
signal \eeprom.delay_counter_10\ : std_logic;
signal \eeprom.delay_counter_8\ : std_logic;
signal \eeprom.delay_counter_6\ : std_logic;
signal \eeprom.n26_adj_388\ : std_logic;
signal \eeprom.n27\ : std_logic;
signal \eeprom.n28_cascade_\ : std_logic;
signal \eeprom.n25\ : std_logic;
signal \eeprom.n1703_cascade_\ : std_logic;
signal \eeprom.n730\ : std_logic;
signal \bfn_21_8_0_\ : std_logic;
signal \eeprom.i2c.n2686\ : std_logic;
signal \eeprom.i2c.n2687\ : std_logic;
signal \eeprom.i2c.n2688\ : std_logic;
signal \eeprom.i2c.n2689\ : std_logic;
signal \eeprom.i2c.n2690\ : std_logic;
signal \eeprom.i2c.n10_adj_384_cascade_\ : std_logic;
signal \eeprom.i2c.n10_adj_377\ : std_logic;
signal \eeprom.i2c.n2972\ : std_logic;
signal \INVeeprom.i2c.data_out_i0_i1C_net\ : std_logic;
signal \INVeeprom.i2c.data_out_i0_i3C_net\ : std_logic;
signal data_2 : std_logic;
signal data_1 : std_logic;
signal data_3 : std_logic;
signal data_0 : std_logic;
signal \n10_cascade_\ : std_logic;
signal \eeprom.n4\ : std_logic;
signal \eeprom.n22\ : std_logic;
signal \eeprom.n26\ : std_logic;
signal \eeprom.n2727\ : std_logic;
signal \eeprom.n2727_cascade_\ : std_logic;
signal \eeprom.i2c.n2881\ : std_logic;
signal read : std_logic;
signal \eeprom.n1703\ : std_logic;
signal \n805_cascade_\ : std_logic;
signal state_1 : std_logic;
signal state_0 : std_logic;
signal data_ready : std_logic;
signal n2476 : std_logic;
signal \n2476_cascade_\ : std_logic;
signal n15 : std_logic;
signal \ID_READOUT_FSM_state_1\ : std_logic;
signal n20 : std_logic;
signal \ID_READOUT_FSM_state_0\ : std_logic;
signal \n20_cascade_\ : std_logic;
signal n6 : std_logic;
signal n1841 : std_logic;
signal \eeprom.i2c.n9_cascade_\ : std_logic;
signal \eeprom.i2c.n2873\ : std_logic;
signal \eeprom.i2c.counter2_2\ : std_logic;
signal \eeprom.i2c.counter2_5\ : std_logic;
signal \eeprom.i2c.counter2_4\ : std_logic;
signal \eeprom.i2c.counter2_3\ : std_logic;
signal \eeprom.i2c.counter2_1\ : std_logic;
signal \eeprom.i2c.n10_adj_379_cascade_\ : std_logic;
signal \eeprom.i2c.counter2_0\ : std_logic;
signal \eeprom.i2c.n1171\ : std_logic;
signal \eeprom.i2c.n2927\ : std_logic;
signal n4 : std_logic;
signal \n4_cascade_\ : std_logic;
signal \eeprom.i2c.n2951_cascade_\ : std_logic;
signal \eeprom.i2c.n37_cascade_\ : std_logic;
signal \eeprom.i2c.n1935\ : std_logic;
signal \eeprom.i2c.n15_cascade_\ : std_logic;
signal \eeprom.i2c.n2454\ : std_logic;
signal \eeprom.i2c.n15\ : std_logic;
signal \bfn_22_11_0_\ : std_logic;
signal \eeprom.i2c.n2664\ : std_logic;
signal \eeprom.i2c.n2665\ : std_logic;
signal \eeprom.i2c.counter_3\ : std_logic;
signal \eeprom.i2c.n2666\ : std_logic;
signal \eeprom.i2c.counter_4\ : std_logic;
signal \eeprom.i2c.n2667\ : std_logic;
signal \eeprom.i2c.counter_5\ : std_logic;
signal \eeprom.i2c.n2668\ : std_logic;
signal \eeprom.i2c.counter_6\ : std_logic;
signal \eeprom.i2c.n2669\ : std_logic;
signal \eeprom.i2c.n2670\ : std_logic;
signal \eeprom.i2c.counter_7\ : std_logic;
signal n14_adj_395 : std_logic;
signal \n4_adj_394_cascade_\ : std_logic;
signal data_4 : std_logic;
signal n1717 : std_logic;
signal data_6 : std_logic;
signal n2424 : std_logic;
signal \n2424_cascade_\ : std_logic;
signal data_7 : std_logic;
signal n4_adj_394 : std_logic;
signal n1722 : std_logic;
signal data_5 : std_logic;
signal \INVeeprom.i2c.data_out_i0_i4C_net\ : std_logic;
signal n4_adj_393 : std_logic;
signal n14 : std_logic;
signal \n13_cascade_\ : std_logic;
signal \n18_cascade_\ : std_logic;
signal \n2935_cascade_\ : std_logic;
signal n2939 : std_logic;
signal \n36_cascade_\ : std_logic;
signal \n22_cascade_\ : std_logic;
signal \n25_cascade_\ : std_logic;
signal n104 : std_logic;
signal n24 : std_logic;
signal n23 : std_logic;
signal \eeprom.i2c.n1837\ : std_logic;
signal \eeprom.i2c.n1928\ : std_logic;
signal \eeprom.i2c.n37\ : std_logic;
signal \eeprom.i2c.n33\ : std_logic;
signal \eeprom.i2c.n9\ : std_logic;
signal \eeprom.i2c.n10_adj_384\ : std_logic;
signal \eeprom.i2c.n1739_cascade_\ : std_logic;
signal \eeprom.i2c.n1054\ : std_logic;
signal n2414 : std_logic;
signal \n1061_cascade_\ : std_logic;
signal \eeprom.i2c.n2869\ : std_logic;
signal \state_7_N_289_3\ : std_logic;
signal n1061 : std_logic;
signal \eeprom.i2c.n2479\ : std_logic;
signal \eeprom.i2c.n10\ : std_logic;
signal \eeprom.i2c.n7\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal n2434 : std_logic;
signal \n2434_cascade_\ : std_logic;
signal n2958 : std_logic;
signal \eeprom.i2c.counter_1\ : std_logic;
signal \eeprom.i2c.counter_0\ : std_logic;
signal \eeprom.i2c.counter_2\ : std_logic;
signal \eeprom.i2c.n2967_cascade_\ : std_logic;
signal rw : std_logic;
signal saved_addr_0 : std_logic;
signal \eeprom.enable\ : std_logic;
signal delay_counter_0 : std_logic;
signal \bfn_23_13_0_\ : std_logic;
signal delay_counter_1 : std_logic;
signal n2633 : std_logic;
signal delay_counter_2 : std_logic;
signal n2634 : std_logic;
signal delay_counter_3 : std_logic;
signal n2635 : std_logic;
signal delay_counter_4 : std_logic;
signal n2636 : std_logic;
signal delay_counter_5 : std_logic;
signal n2637 : std_logic;
signal delay_counter_6 : std_logic;
signal n2638 : std_logic;
signal delay_counter_7 : std_logic;
signal n2639 : std_logic;
signal n2640 : std_logic;
signal delay_counter_8 : std_logic;
signal \bfn_23_14_0_\ : std_logic;
signal delay_counter_9 : std_logic;
signal n2641 : std_logic;
signal delay_counter_10 : std_logic;
signal n2642 : std_logic;
signal delay_counter_11 : std_logic;
signal n2643 : std_logic;
signal delay_counter_12 : std_logic;
signal n2644 : std_logic;
signal delay_counter_13 : std_logic;
signal n2645 : std_logic;
signal delay_counter_14 : std_logic;
signal n2646 : std_logic;
signal delay_counter_15 : std_logic;
signal n2647 : std_logic;
signal n2648 : std_logic;
signal delay_counter_16 : std_logic;
signal \bfn_23_15_0_\ : std_logic;
signal delay_counter_17 : std_logic;
signal n2649 : std_logic;
signal delay_counter_18 : std_logic;
signal n2650 : std_logic;
signal delay_counter_19 : std_logic;
signal n2651 : std_logic;
signal delay_counter_20 : std_logic;
signal n2652 : std_logic;
signal delay_counter_21 : std_logic;
signal n2653 : std_logic;
signal delay_counter_22 : std_logic;
signal n2654 : std_logic;
signal delay_counter_23 : std_logic;
signal n2655 : std_logic;
signal n2656 : std_logic;
signal delay_counter_24 : std_logic;
signal \bfn_23_16_0_\ : std_logic;
signal delay_counter_25 : std_logic;
signal n2657 : std_logic;
signal delay_counter_26 : std_logic;
signal n2658 : std_logic;
signal delay_counter_27 : std_logic;
signal n2659 : std_logic;
signal delay_counter_28 : std_logic;
signal n2660 : std_logic;
signal delay_counter_29 : std_logic;
signal n2661 : std_logic;
signal delay_counter_30 : std_logic;
signal n2662 : std_logic;
signal n2663 : std_logic;
signal delay_counter_31 : std_logic;
signal n1740 : std_logic;
signal n1895 : std_logic;
signal sda_out : std_logic;
signal sda_enable : std_logic;
signal \INVeeprom.i2c.write_enable_130C_net\ : std_logic;
signal \eeprom.i2c.n1152\ : std_logic;
signal \eeprom.i2c.n1932\ : std_logic;
signal \eeprom.i2c.n11_adj_378\ : std_logic;
signal \eeprom.i2c.n13\ : std_logic;
signal \eeprom.i2c.n11_adj_381\ : std_logic;
signal \eeprom.i2c.n2963\ : std_logic;
signal \eeprom.i2c.n11\ : std_logic;
signal \eeprom.i2c.sda_out_adj_376\ : std_logic;
signal \INVeeprom.i2c.sda_out_131C_net\ : std_logic;
signal \eeprom.i2c.n2791\ : std_logic;
signal \eeprom.i2c.n11_adj_380\ : std_logic;
signal state_0_adj_392 : std_logic;
signal \eeprom.state_3\ : std_logic;
signal \eeprom.i2c.state_1_adj_375\ : std_logic;
signal \eeprom.i2c.state_2\ : std_logic;
signal \INVeeprom.i2c.i2c_scl_enable_123C_net\ : std_logic;
signal n47 : std_logic;
signal \state_7_N_273_0\ : std_logic;
signal \CLK_c\ : std_logic;
signal \eeprom.i2c.n1766\ : std_logic;
signal \eeprom.i2c.i2c_clk\ : std_logic;
signal scl_enable : std_logic;
signal scl_c : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CS_CLK_wire\ : std_logic;
signal \CS_wire\ : std_logic;
signal \DE_wire\ : std_logic;
signal \INHA_wire\ : std_logic;
signal \INHB_wire\ : std_logic;
signal \INHC_wire\ : std_logic;
signal \INLA_wire\ : std_logic;
signal \INLB_wire\ : std_logic;
signal \INLC_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \NEOPXL_wire\ : std_logic;
signal \TX_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    CS_CLK <= \CS_CLK_wire\;
    CS <= \CS_wire\;
    DE <= \DE_wire\;
    INHA <= \INHA_wire\;
    INHB <= \INHB_wire\;
    INHC <= \INHC_wire\;
    INLA <= \INLA_wire\;
    INLB <= \INLB_wire\;
    INLC <= \INLC_wire\;
    LED <= \LED_wire\;
    NEOPXL <= \NEOPXL_wire\;
    TX <= \TX_wire\;
    USBPU <= \USBPU_wire\;
    \CLK_wire\ <= CLK;

    \CS_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6680\,
            DIN => \N__6679\,
            DOUT => \N__6678\,
            PACKAGEPIN => \CS_CLK_wire\
        );

    \CS_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6680\,
            PADOUT => \N__6679\,
            PADIN => \N__6678\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \CS_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6671\,
            DIN => \N__6670\,
            DOUT => \N__6669\,
            PACKAGEPIN => \CS_wire\
        );

    \CS_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6671\,
            PADOUT => \N__6670\,
            PADIN => \N__6669\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \DE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6662\,
            DIN => \N__6661\,
            DOUT => \N__6660\,
            PACKAGEPIN => \DE_wire\
        );

    \DE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6662\,
            PADOUT => \N__6661\,
            PADIN => \N__6660\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHA_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6653\,
            DIN => \N__6652\,
            DOUT => \N__6651\,
            PACKAGEPIN => \INHA_wire\
        );

    \INHA_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6653\,
            PADOUT => \N__6652\,
            PADIN => \N__6651\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHB_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6644\,
            DIN => \N__6643\,
            DOUT => \N__6642\,
            PACKAGEPIN => \INHB_wire\
        );

    \INHB_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6644\,
            PADOUT => \N__6643\,
            PADIN => \N__6642\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6635\,
            DIN => \N__6634\,
            DOUT => \N__6633\,
            PACKAGEPIN => \INHC_wire\
        );

    \INHC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6635\,
            PADOUT => \N__6634\,
            PADIN => \N__6633\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLA_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6626\,
            DIN => \N__6625\,
            DOUT => \N__6624\,
            PACKAGEPIN => \INLA_wire\
        );

    \INLA_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6626\,
            PADOUT => \N__6625\,
            PADIN => \N__6624\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLB_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6617\,
            DIN => \N__6616\,
            DOUT => \N__6615\,
            PACKAGEPIN => \INLB_wire\
        );

    \INLB_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6617\,
            PADOUT => \N__6616\,
            PADIN => \N__6615\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6608\,
            DIN => \N__6607\,
            DOUT => \N__6606\,
            PACKAGEPIN => \INLC_wire\
        );

    \INLC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6608\,
            PADOUT => \N__6607\,
            PADIN => \N__6606\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6599\,
            DIN => \N__6598\,
            DOUT => \N__6597\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6599\,
            PADOUT => \N__6598\,
            PADIN => \N__6597\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__2782\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \NEOPXL_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6590\,
            DIN => \N__6589\,
            DOUT => \N__6588\,
            PACKAGEPIN => \NEOPXL_wire\
        );

    \NEOPXL_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6590\,
            PADOUT => \N__6589\,
            PADIN => \N__6588\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \TX_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6581\,
            DIN => \N__6580\,
            DOUT => \N__6579\,
            PACKAGEPIN => \TX_wire\
        );

    \TX_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6581\,
            PADOUT => \N__6580\,
            PADIN => \N__6579\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6572\,
            DIN => \N__6571\,
            DOUT => \N__6570\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6572\,
            PADOUT => \N__6571\,
            PADIN => \N__6570\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \scl_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__6563\,
            DIN => \N__6562\,
            DOUT => \N__6561\,
            PACKAGEPIN => SCL
        );

    \scl_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6563\,
            PADOUT => \N__6562\,
            PADIN => \N__6561\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__5605\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__5638\
        );

    \sda_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__6554\,
            DIN => \N__6553\,
            DOUT => \N__6552\,
            PACKAGEPIN => SDA
        );

    \sda_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6554\,
            PADOUT => \N__6553\,
            PADIN => \N__6552\,
            CLOCKENABLE => 'H',
            DIN0 => \state_7_N_289_3\,
            DIN1 => OPEN,
            DOUT0 => \N__5428\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__5410\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6545\,
            DIN => \N__6544\,
            DOUT => \N__6543\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6545\,
            PADOUT => \N__6544\,
            PADIN => \N__6543\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__1503\ : InMux
    port map (
            O => \N__6526\,
            I => \N__6523\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__6523\,
            I => \eeprom.i2c.n2963\
        );

    \I__1501\ : CascadeMux
    port map (
            O => \N__6520\,
            I => \N__6517\
        );

    \I__1500\ : InMux
    port map (
            O => \N__6517\,
            I => \N__6514\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__6514\,
            I => \N__6509\
        );

    \I__1498\ : InMux
    port map (
            O => \N__6513\,
            I => \N__6506\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__6512\,
            I => \N__6503\
        );

    \I__1496\ : Span4Mux_v
    port map (
            O => \N__6509\,
            I => \N__6500\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__6506\,
            I => \N__6497\
        );

    \I__1494\ : InMux
    port map (
            O => \N__6503\,
            I => \N__6494\
        );

    \I__1493\ : Odrv4
    port map (
            O => \N__6500\,
            I => \eeprom.i2c.n11\
        );

    \I__1492\ : Odrv12
    port map (
            O => \N__6497\,
            I => \eeprom.i2c.n11\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__6494\,
            I => \eeprom.i2c.n11\
        );

    \I__1490\ : InMux
    port map (
            O => \N__6487\,
            I => \N__6484\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__6484\,
            I => \N__6481\
        );

    \I__1488\ : Odrv12
    port map (
            O => \N__6481\,
            I => \eeprom.i2c.sda_out_adj_376\
        );

    \I__1487\ : CEMux
    port map (
            O => \N__6478\,
            I => \N__6475\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__6475\,
            I => \N__6472\
        );

    \I__1485\ : Odrv4
    port map (
            O => \N__6472\,
            I => \eeprom.i2c.n2791\
        );

    \I__1484\ : InMux
    port map (
            O => \N__6469\,
            I => \N__6466\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__6466\,
            I => \N__6463\
        );

    \I__1482\ : Odrv4
    port map (
            O => \N__6463\,
            I => \eeprom.i2c.n11_adj_380\
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__6460\,
            I => \N__6456\
        );

    \I__1480\ : InMux
    port map (
            O => \N__6459\,
            I => \N__6453\
        );

    \I__1479\ : InMux
    port map (
            O => \N__6456\,
            I => \N__6450\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__6453\,
            I => \N__6441\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__6450\,
            I => \N__6438\
        );

    \I__1476\ : InMux
    port map (
            O => \N__6449\,
            I => \N__6434\
        );

    \I__1475\ : InMux
    port map (
            O => \N__6448\,
            I => \N__6431\
        );

    \I__1474\ : InMux
    port map (
            O => \N__6447\,
            I => \N__6423\
        );

    \I__1473\ : InMux
    port map (
            O => \N__6446\,
            I => \N__6423\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__6445\,
            I => \N__6414\
        );

    \I__1471\ : CascadeMux
    port map (
            O => \N__6444\,
            I => \N__6411\
        );

    \I__1470\ : Span4Mux_v
    port map (
            O => \N__6441\,
            I => \N__6405\
        );

    \I__1469\ : Span4Mux_h
    port map (
            O => \N__6438\,
            I => \N__6402\
        );

    \I__1468\ : InMux
    port map (
            O => \N__6437\,
            I => \N__6399\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__6434\,
            I => \N__6394\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__6431\,
            I => \N__6394\
        );

    \I__1465\ : InMux
    port map (
            O => \N__6430\,
            I => \N__6391\
        );

    \I__1464\ : InMux
    port map (
            O => \N__6429\,
            I => \N__6386\
        );

    \I__1463\ : InMux
    port map (
            O => \N__6428\,
            I => \N__6386\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__6423\,
            I => \N__6383\
        );

    \I__1461\ : InMux
    port map (
            O => \N__6422\,
            I => \N__6376\
        );

    \I__1460\ : InMux
    port map (
            O => \N__6421\,
            I => \N__6376\
        );

    \I__1459\ : InMux
    port map (
            O => \N__6420\,
            I => \N__6376\
        );

    \I__1458\ : InMux
    port map (
            O => \N__6419\,
            I => \N__6371\
        );

    \I__1457\ : InMux
    port map (
            O => \N__6418\,
            I => \N__6371\
        );

    \I__1456\ : InMux
    port map (
            O => \N__6417\,
            I => \N__6368\
        );

    \I__1455\ : InMux
    port map (
            O => \N__6414\,
            I => \N__6361\
        );

    \I__1454\ : InMux
    port map (
            O => \N__6411\,
            I => \N__6361\
        );

    \I__1453\ : InMux
    port map (
            O => \N__6410\,
            I => \N__6361\
        );

    \I__1452\ : InMux
    port map (
            O => \N__6409\,
            I => \N__6356\
        );

    \I__1451\ : InMux
    port map (
            O => \N__6408\,
            I => \N__6356\
        );

    \I__1450\ : Odrv4
    port map (
            O => \N__6405\,
            I => state_0_adj_392
        );

    \I__1449\ : Odrv4
    port map (
            O => \N__6402\,
            I => state_0_adj_392
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__6399\,
            I => state_0_adj_392
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__6394\,
            I => state_0_adj_392
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__6391\,
            I => state_0_adj_392
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__6386\,
            I => state_0_adj_392
        );

    \I__1444\ : Odrv4
    port map (
            O => \N__6383\,
            I => state_0_adj_392
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__6376\,
            I => state_0_adj_392
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__6371\,
            I => state_0_adj_392
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__6368\,
            I => state_0_adj_392
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__6361\,
            I => state_0_adj_392
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__6356\,
            I => state_0_adj_392
        );

    \I__1438\ : CascadeMux
    port map (
            O => \N__6331\,
            I => \N__6324\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__6330\,
            I => \N__6321\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__6329\,
            I => \N__6313\
        );

    \I__1435\ : InMux
    port map (
            O => \N__6328\,
            I => \N__6309\
        );

    \I__1434\ : InMux
    port map (
            O => \N__6327\,
            I => \N__6306\
        );

    \I__1433\ : InMux
    port map (
            O => \N__6324\,
            I => \N__6302\
        );

    \I__1432\ : InMux
    port map (
            O => \N__6321\,
            I => \N__6299\
        );

    \I__1431\ : InMux
    port map (
            O => \N__6320\,
            I => \N__6292\
        );

    \I__1430\ : InMux
    port map (
            O => \N__6319\,
            I => \N__6292\
        );

    \I__1429\ : InMux
    port map (
            O => \N__6318\,
            I => \N__6285\
        );

    \I__1428\ : InMux
    port map (
            O => \N__6317\,
            I => \N__6285\
        );

    \I__1427\ : InMux
    port map (
            O => \N__6316\,
            I => \N__6285\
        );

    \I__1426\ : InMux
    port map (
            O => \N__6313\,
            I => \N__6282\
        );

    \I__1425\ : InMux
    port map (
            O => \N__6312\,
            I => \N__6277\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__6309\,
            I => \N__6274\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__6306\,
            I => \N__6271\
        );

    \I__1422\ : InMux
    port map (
            O => \N__6305\,
            I => \N__6268\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__6302\,
            I => \N__6264\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__6299\,
            I => \N__6261\
        );

    \I__1419\ : InMux
    port map (
            O => \N__6298\,
            I => \N__6256\
        );

    \I__1418\ : InMux
    port map (
            O => \N__6297\,
            I => \N__6256\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__6292\,
            I => \N__6250\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__6285\,
            I => \N__6250\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__6282\,
            I => \N__6245\
        );

    \I__1414\ : InMux
    port map (
            O => \N__6281\,
            I => \N__6242\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6280\,
            I => \N__6239\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__6277\,
            I => \N__6230\
        );

    \I__1411\ : Span4Mux_v
    port map (
            O => \N__6274\,
            I => \N__6230\
        );

    \I__1410\ : Span4Mux_h
    port map (
            O => \N__6271\,
            I => \N__6230\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__6268\,
            I => \N__6230\
        );

    \I__1408\ : InMux
    port map (
            O => \N__6267\,
            I => \N__6227\
        );

    \I__1407\ : Span4Mux_h
    port map (
            O => \N__6264\,
            I => \N__6220\
        );

    \I__1406\ : Span4Mux_h
    port map (
            O => \N__6261\,
            I => \N__6220\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__6256\,
            I => \N__6220\
        );

    \I__1404\ : InMux
    port map (
            O => \N__6255\,
            I => \N__6217\
        );

    \I__1403\ : Span4Mux_h
    port map (
            O => \N__6250\,
            I => \N__6214\
        );

    \I__1402\ : InMux
    port map (
            O => \N__6249\,
            I => \N__6209\
        );

    \I__1401\ : InMux
    port map (
            O => \N__6248\,
            I => \N__6209\
        );

    \I__1400\ : Odrv12
    port map (
            O => \N__6245\,
            I => \eeprom.state_3\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__6242\,
            I => \eeprom.state_3\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__6239\,
            I => \eeprom.state_3\
        );

    \I__1397\ : Odrv4
    port map (
            O => \N__6230\,
            I => \eeprom.state_3\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__6227\,
            I => \eeprom.state_3\
        );

    \I__1395\ : Odrv4
    port map (
            O => \N__6220\,
            I => \eeprom.state_3\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__6217\,
            I => \eeprom.state_3\
        );

    \I__1393\ : Odrv4
    port map (
            O => \N__6214\,
            I => \eeprom.state_3\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__6209\,
            I => \eeprom.state_3\
        );

    \I__1391\ : InMux
    port map (
            O => \N__6190\,
            I => \N__6185\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__6189\,
            I => \N__6181\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__6188\,
            I => \N__6175\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__6185\,
            I => \N__6167\
        );

    \I__1387\ : InMux
    port map (
            O => \N__6184\,
            I => \N__6164\
        );

    \I__1386\ : InMux
    port map (
            O => \N__6181\,
            I => \N__6161\
        );

    \I__1385\ : CascadeMux
    port map (
            O => \N__6180\,
            I => \N__6158\
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__6179\,
            I => \N__6150\
        );

    \I__1383\ : InMux
    port map (
            O => \N__6178\,
            I => \N__6141\
        );

    \I__1382\ : InMux
    port map (
            O => \N__6175\,
            I => \N__6141\
        );

    \I__1381\ : InMux
    port map (
            O => \N__6174\,
            I => \N__6141\
        );

    \I__1380\ : InMux
    port map (
            O => \N__6173\,
            I => \N__6141\
        );

    \I__1379\ : InMux
    port map (
            O => \N__6172\,
            I => \N__6136\
        );

    \I__1378\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6136\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__6170\,
            I => \N__6131\
        );

    \I__1376\ : Span4Mux_v
    port map (
            O => \N__6167\,
            I => \N__6126\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__6164\,
            I => \N__6126\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__6161\,
            I => \N__6123\
        );

    \I__1373\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6120\
        );

    \I__1372\ : InMux
    port map (
            O => \N__6157\,
            I => \N__6117\
        );

    \I__1371\ : InMux
    port map (
            O => \N__6156\,
            I => \N__6112\
        );

    \I__1370\ : InMux
    port map (
            O => \N__6155\,
            I => \N__6112\
        );

    \I__1369\ : InMux
    port map (
            O => \N__6154\,
            I => \N__6107\
        );

    \I__1368\ : InMux
    port map (
            O => \N__6153\,
            I => \N__6107\
        );

    \I__1367\ : InMux
    port map (
            O => \N__6150\,
            I => \N__6104\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__6141\,
            I => \N__6099\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__6136\,
            I => \N__6099\
        );

    \I__1364\ : InMux
    port map (
            O => \N__6135\,
            I => \N__6092\
        );

    \I__1363\ : InMux
    port map (
            O => \N__6134\,
            I => \N__6092\
        );

    \I__1362\ : InMux
    port map (
            O => \N__6131\,
            I => \N__6092\
        );

    \I__1361\ : Odrv4
    port map (
            O => \N__6126\,
            I => \eeprom.i2c.state_1_adj_375\
        );

    \I__1360\ : Odrv4
    port map (
            O => \N__6123\,
            I => \eeprom.i2c.state_1_adj_375\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__6120\,
            I => \eeprom.i2c.state_1_adj_375\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__6117\,
            I => \eeprom.i2c.state_1_adj_375\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__6112\,
            I => \eeprom.i2c.state_1_adj_375\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__6107\,
            I => \eeprom.i2c.state_1_adj_375\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__6104\,
            I => \eeprom.i2c.state_1_adj_375\
        );

    \I__1354\ : Odrv4
    port map (
            O => \N__6099\,
            I => \eeprom.i2c.state_1_adj_375\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__6092\,
            I => \eeprom.i2c.state_1_adj_375\
        );

    \I__1352\ : CascadeMux
    port map (
            O => \N__6073\,
            I => \N__6064\
        );

    \I__1351\ : InMux
    port map (
            O => \N__6072\,
            I => \N__6061\
        );

    \I__1350\ : InMux
    port map (
            O => \N__6071\,
            I => \N__6058\
        );

    \I__1349\ : InMux
    port map (
            O => \N__6070\,
            I => \N__6051\
        );

    \I__1348\ : InMux
    port map (
            O => \N__6069\,
            I => \N__6046\
        );

    \I__1347\ : InMux
    port map (
            O => \N__6068\,
            I => \N__6046\
        );

    \I__1346\ : InMux
    port map (
            O => \N__6067\,
            I => \N__6043\
        );

    \I__1345\ : InMux
    port map (
            O => \N__6064\,
            I => \N__6033\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__6061\,
            I => \N__6030\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__6058\,
            I => \N__6027\
        );

    \I__1342\ : InMux
    port map (
            O => \N__6057\,
            I => \N__6022\
        );

    \I__1341\ : InMux
    port map (
            O => \N__6056\,
            I => \N__6022\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6055\,
            I => \N__6017\
        );

    \I__1339\ : InMux
    port map (
            O => \N__6054\,
            I => \N__6017\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__6051\,
            I => \N__6012\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__6046\,
            I => \N__6012\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__6043\,
            I => \N__6005\
        );

    \I__1335\ : InMux
    port map (
            O => \N__6042\,
            I => \N__6000\
        );

    \I__1334\ : InMux
    port map (
            O => \N__6041\,
            I => \N__6000\
        );

    \I__1333\ : InMux
    port map (
            O => \N__6040\,
            I => \N__5995\
        );

    \I__1332\ : InMux
    port map (
            O => \N__6039\,
            I => \N__5995\
        );

    \I__1331\ : InMux
    port map (
            O => \N__6038\,
            I => \N__5988\
        );

    \I__1330\ : InMux
    port map (
            O => \N__6037\,
            I => \N__5988\
        );

    \I__1329\ : InMux
    port map (
            O => \N__6036\,
            I => \N__5988\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__6033\,
            I => \N__5985\
        );

    \I__1327\ : Span4Mux_v
    port map (
            O => \N__6030\,
            I => \N__5974\
        );

    \I__1326\ : Span4Mux_v
    port map (
            O => \N__6027\,
            I => \N__5974\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__6022\,
            I => \N__5974\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__6017\,
            I => \N__5974\
        );

    \I__1323\ : Span4Mux_v
    port map (
            O => \N__6012\,
            I => \N__5974\
        );

    \I__1322\ : InMux
    port map (
            O => \N__6011\,
            I => \N__5971\
        );

    \I__1321\ : InMux
    port map (
            O => \N__6010\,
            I => \N__5964\
        );

    \I__1320\ : InMux
    port map (
            O => \N__6009\,
            I => \N__5964\
        );

    \I__1319\ : InMux
    port map (
            O => \N__6008\,
            I => \N__5964\
        );

    \I__1318\ : Odrv4
    port map (
            O => \N__6005\,
            I => \eeprom.i2c.state_2\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__6000\,
            I => \eeprom.i2c.state_2\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__5995\,
            I => \eeprom.i2c.state_2\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__5988\,
            I => \eeprom.i2c.state_2\
        );

    \I__1314\ : Odrv4
    port map (
            O => \N__5985\,
            I => \eeprom.i2c.state_2\
        );

    \I__1313\ : Odrv4
    port map (
            O => \N__5974\,
            I => \eeprom.i2c.state_2\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__5971\,
            I => \eeprom.i2c.state_2\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__5964\,
            I => \eeprom.i2c.state_2\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__5947\,
            I => \N__5943\
        );

    \I__1309\ : InMux
    port map (
            O => \N__5946\,
            I => \N__5935\
        );

    \I__1308\ : InMux
    port map (
            O => \N__5943\,
            I => \N__5935\
        );

    \I__1307\ : InMux
    port map (
            O => \N__5942\,
            I => \N__5932\
        );

    \I__1306\ : InMux
    port map (
            O => \N__5941\,
            I => \N__5929\
        );

    \I__1305\ : InMux
    port map (
            O => \N__5940\,
            I => \N__5926\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__5935\,
            I => \N__5920\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__5932\,
            I => \N__5920\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__5929\,
            I => \N__5915\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__5926\,
            I => \N__5915\
        );

    \I__1300\ : InMux
    port map (
            O => \N__5925\,
            I => \N__5912\
        );

    \I__1299\ : Span4Mux_v
    port map (
            O => \N__5920\,
            I => \N__5906\
        );

    \I__1298\ : Span4Mux_v
    port map (
            O => \N__5915\,
            I => \N__5903\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__5912\,
            I => \N__5900\
        );

    \I__1296\ : InMux
    port map (
            O => \N__5911\,
            I => \N__5897\
        );

    \I__1295\ : InMux
    port map (
            O => \N__5910\,
            I => \N__5892\
        );

    \I__1294\ : InMux
    port map (
            O => \N__5909\,
            I => \N__5892\
        );

    \I__1293\ : Odrv4
    port map (
            O => \N__5906\,
            I => n47
        );

    \I__1292\ : Odrv4
    port map (
            O => \N__5903\,
            I => n47
        );

    \I__1291\ : Odrv4
    port map (
            O => \N__5900\,
            I => n47
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__5897\,
            I => n47
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5892\,
            I => n47
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__5881\,
            I => \N__5877\
        );

    \I__1287\ : InMux
    port map (
            O => \N__5880\,
            I => \N__5872\
        );

    \I__1286\ : InMux
    port map (
            O => \N__5877\,
            I => \N__5872\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__5872\,
            I => \N__5869\
        );

    \I__1284\ : Span4Mux_v
    port map (
            O => \N__5869\,
            I => \N__5864\
        );

    \I__1283\ : InMux
    port map (
            O => \N__5868\,
            I => \N__5861\
        );

    \I__1282\ : InMux
    port map (
            O => \N__5867\,
            I => \N__5858\
        );

    \I__1281\ : Odrv4
    port map (
            O => \N__5864\,
            I => \state_7_N_273_0\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__5861\,
            I => \state_7_N_273_0\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__5858\,
            I => \state_7_N_273_0\
        );

    \I__1278\ : ClkMux
    port map (
            O => \N__5851\,
            I => \N__5800\
        );

    \I__1277\ : ClkMux
    port map (
            O => \N__5850\,
            I => \N__5800\
        );

    \I__1276\ : ClkMux
    port map (
            O => \N__5849\,
            I => \N__5800\
        );

    \I__1275\ : ClkMux
    port map (
            O => \N__5848\,
            I => \N__5800\
        );

    \I__1274\ : ClkMux
    port map (
            O => \N__5847\,
            I => \N__5800\
        );

    \I__1273\ : ClkMux
    port map (
            O => \N__5846\,
            I => \N__5800\
        );

    \I__1272\ : ClkMux
    port map (
            O => \N__5845\,
            I => \N__5800\
        );

    \I__1271\ : ClkMux
    port map (
            O => \N__5844\,
            I => \N__5800\
        );

    \I__1270\ : ClkMux
    port map (
            O => \N__5843\,
            I => \N__5800\
        );

    \I__1269\ : ClkMux
    port map (
            O => \N__5842\,
            I => \N__5800\
        );

    \I__1268\ : ClkMux
    port map (
            O => \N__5841\,
            I => \N__5800\
        );

    \I__1267\ : ClkMux
    port map (
            O => \N__5840\,
            I => \N__5800\
        );

    \I__1266\ : ClkMux
    port map (
            O => \N__5839\,
            I => \N__5800\
        );

    \I__1265\ : ClkMux
    port map (
            O => \N__5838\,
            I => \N__5800\
        );

    \I__1264\ : ClkMux
    port map (
            O => \N__5837\,
            I => \N__5800\
        );

    \I__1263\ : ClkMux
    port map (
            O => \N__5836\,
            I => \N__5800\
        );

    \I__1262\ : ClkMux
    port map (
            O => \N__5835\,
            I => \N__5800\
        );

    \I__1261\ : GlobalMux
    port map (
            O => \N__5800\,
            I => \N__5797\
        );

    \I__1260\ : gio2CtrlBuf
    port map (
            O => \N__5797\,
            I => \CLK_c\
        );

    \I__1259\ : CEMux
    port map (
            O => \N__5794\,
            I => \N__5791\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__5791\,
            I => \N__5788\
        );

    \I__1257\ : Span4Mux_h
    port map (
            O => \N__5788\,
            I => \N__5785\
        );

    \I__1256\ : Odrv4
    port map (
            O => \N__5785\,
            I => \eeprom.i2c.n1766\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5782\,
            I => \N__5779\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__5779\,
            I => \N__5776\
        );

    \I__1253\ : Span4Mux_v
    port map (
            O => \N__5776\,
            I => \N__5772\
        );

    \I__1252\ : ClkMux
    port map (
            O => \N__5775\,
            I => \N__5768\
        );

    \I__1251\ : Span4Mux_h
    port map (
            O => \N__5772\,
            I => \N__5761\
        );

    \I__1250\ : ClkMux
    port map (
            O => \N__5771\,
            I => \N__5758\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__5768\,
            I => \N__5753\
        );

    \I__1248\ : ClkMux
    port map (
            O => \N__5767\,
            I => \N__5750\
        );

    \I__1247\ : ClkMux
    port map (
            O => \N__5766\,
            I => \N__5746\
        );

    \I__1246\ : ClkMux
    port map (
            O => \N__5765\,
            I => \N__5743\
        );

    \I__1245\ : ClkMux
    port map (
            O => \N__5764\,
            I => \N__5738\
        );

    \I__1244\ : Span4Mux_v
    port map (
            O => \N__5761\,
            I => \N__5732\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__5758\,
            I => \N__5732\
        );

    \I__1242\ : ClkMux
    port map (
            O => \N__5757\,
            I => \N__5729\
        );

    \I__1241\ : ClkMux
    port map (
            O => \N__5756\,
            I => \N__5725\
        );

    \I__1240\ : Span4Mux_v
    port map (
            O => \N__5753\,
            I => \N__5720\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__5750\,
            I => \N__5720\
        );

    \I__1238\ : ClkMux
    port map (
            O => \N__5749\,
            I => \N__5717\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__5746\,
            I => \N__5712\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__5743\,
            I => \N__5712\
        );

    \I__1235\ : ClkMux
    port map (
            O => \N__5742\,
            I => \N__5709\
        );

    \I__1234\ : ClkMux
    port map (
            O => \N__5741\,
            I => \N__5706\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__5738\,
            I => \N__5703\
        );

    \I__1232\ : ClkMux
    port map (
            O => \N__5737\,
            I => \N__5700\
        );

    \I__1231\ : Span4Mux_v
    port map (
            O => \N__5732\,
            I => \N__5695\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__5729\,
            I => \N__5695\
        );

    \I__1229\ : ClkMux
    port map (
            O => \N__5728\,
            I => \N__5692\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__5725\,
            I => \N__5689\
        );

    \I__1227\ : Span4Mux_v
    port map (
            O => \N__5720\,
            I => \N__5686\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__5717\,
            I => \N__5683\
        );

    \I__1225\ : Span4Mux_v
    port map (
            O => \N__5712\,
            I => \N__5680\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__5709\,
            I => \N__5677\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__5706\,
            I => \N__5666\
        );

    \I__1222\ : Span4Mux_v
    port map (
            O => \N__5703\,
            I => \N__5666\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__5700\,
            I => \N__5666\
        );

    \I__1220\ : Span4Mux_v
    port map (
            O => \N__5695\,
            I => \N__5666\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5692\,
            I => \N__5666\
        );

    \I__1218\ : Span4Mux_h
    port map (
            O => \N__5689\,
            I => \N__5662\
        );

    \I__1217\ : Span4Mux_v
    port map (
            O => \N__5686\,
            I => \N__5655\
        );

    \I__1216\ : Span4Mux_v
    port map (
            O => \N__5683\,
            I => \N__5655\
        );

    \I__1215\ : Span4Mux_h
    port map (
            O => \N__5680\,
            I => \N__5655\
        );

    \I__1214\ : Span4Mux_v
    port map (
            O => \N__5677\,
            I => \N__5650\
        );

    \I__1213\ : Span4Mux_v
    port map (
            O => \N__5666\,
            I => \N__5650\
        );

    \I__1212\ : InMux
    port map (
            O => \N__5665\,
            I => \N__5647\
        );

    \I__1211\ : Odrv4
    port map (
            O => \N__5662\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1210\ : Odrv4
    port map (
            O => \N__5655\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1209\ : Odrv4
    port map (
            O => \N__5650\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__5647\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__1207\ : IoInMux
    port map (
            O => \N__5638\,
            I => \N__5635\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__5635\,
            I => \N__5632\
        );

    \I__1205\ : IoSpan4Mux
    port map (
            O => \N__5632\,
            I => \N__5629\
        );

    \I__1204\ : Span4Mux_s1_h
    port map (
            O => \N__5629\,
            I => \N__5625\
        );

    \I__1203\ : InMux
    port map (
            O => \N__5628\,
            I => \N__5622\
        );

    \I__1202\ : Span4Mux_h
    port map (
            O => \N__5625\,
            I => \N__5619\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__5622\,
            I => \N__5616\
        );

    \I__1200\ : Span4Mux_v
    port map (
            O => \N__5619\,
            I => \N__5611\
        );

    \I__1199\ : Span4Mux_v
    port map (
            O => \N__5616\,
            I => \N__5611\
        );

    \I__1198\ : Span4Mux_v
    port map (
            O => \N__5611\,
            I => \N__5608\
        );

    \I__1197\ : Odrv4
    port map (
            O => \N__5608\,
            I => scl_enable
        );

    \I__1196\ : IoInMux
    port map (
            O => \N__5605\,
            I => \N__5602\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__5602\,
            I => \N__5599\
        );

    \I__1194\ : IoSpan4Mux
    port map (
            O => \N__5599\,
            I => \N__5596\
        );

    \I__1193\ : Span4Mux_s2_h
    port map (
            O => \N__5596\,
            I => \N__5593\
        );

    \I__1192\ : Odrv4
    port map (
            O => \N__5593\,
            I => scl_c
        );

    \I__1191\ : InMux
    port map (
            O => \N__5590\,
            I => \N__5586\
        );

    \I__1190\ : InMux
    port map (
            O => \N__5589\,
            I => \N__5583\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5586\,
            I => delay_counter_28
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__5583\,
            I => delay_counter_28
        );

    \I__1187\ : InMux
    port map (
            O => \N__5578\,
            I => n2660
        );

    \I__1186\ : CascadeMux
    port map (
            O => \N__5575\,
            I => \N__5571\
        );

    \I__1185\ : InMux
    port map (
            O => \N__5574\,
            I => \N__5568\
        );

    \I__1184\ : InMux
    port map (
            O => \N__5571\,
            I => \N__5565\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__5568\,
            I => delay_counter_29
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__5565\,
            I => delay_counter_29
        );

    \I__1181\ : InMux
    port map (
            O => \N__5560\,
            I => n2661
        );

    \I__1180\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5553\
        );

    \I__1179\ : InMux
    port map (
            O => \N__5556\,
            I => \N__5550\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__5553\,
            I => delay_counter_30
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__5550\,
            I => delay_counter_30
        );

    \I__1176\ : InMux
    port map (
            O => \N__5545\,
            I => n2662
        );

    \I__1175\ : InMux
    port map (
            O => \N__5542\,
            I => n2663
        );

    \I__1174\ : InMux
    port map (
            O => \N__5539\,
            I => \N__5536\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__5536\,
            I => \N__5532\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5535\,
            I => \N__5529\
        );

    \I__1171\ : Span4Mux_h
    port map (
            O => \N__5532\,
            I => \N__5526\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__5529\,
            I => delay_counter_31
        );

    \I__1169\ : Odrv4
    port map (
            O => \N__5526\,
            I => delay_counter_31
        );

    \I__1168\ : CEMux
    port map (
            O => \N__5521\,
            I => \N__5518\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__5518\,
            I => \N__5513\
        );

    \I__1166\ : CEMux
    port map (
            O => \N__5517\,
            I => \N__5510\
        );

    \I__1165\ : CEMux
    port map (
            O => \N__5516\,
            I => \N__5506\
        );

    \I__1164\ : Span4Mux_v
    port map (
            O => \N__5513\,
            I => \N__5501\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__5510\,
            I => \N__5501\
        );

    \I__1162\ : CEMux
    port map (
            O => \N__5509\,
            I => \N__5498\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__5506\,
            I => \N__5493\
        );

    \I__1160\ : Span4Mux_v
    port map (
            O => \N__5501\,
            I => \N__5493\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__5498\,
            I => \N__5490\
        );

    \I__1158\ : Span4Mux_v
    port map (
            O => \N__5493\,
            I => \N__5486\
        );

    \I__1157\ : Span4Mux_h
    port map (
            O => \N__5490\,
            I => \N__5483\
        );

    \I__1156\ : InMux
    port map (
            O => \N__5489\,
            I => \N__5480\
        );

    \I__1155\ : Odrv4
    port map (
            O => \N__5486\,
            I => n1740
        );

    \I__1154\ : Odrv4
    port map (
            O => \N__5483\,
            I => n1740
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__5480\,
            I => n1740
        );

    \I__1152\ : SRMux
    port map (
            O => \N__5473\,
            I => \N__5468\
        );

    \I__1151\ : SRMux
    port map (
            O => \N__5472\,
            I => \N__5465\
        );

    \I__1150\ : SRMux
    port map (
            O => \N__5471\,
            I => \N__5462\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__5468\,
            I => \N__5459\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__5465\,
            I => \N__5456\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__5462\,
            I => \N__5452\
        );

    \I__1146\ : Span4Mux_v
    port map (
            O => \N__5459\,
            I => \N__5447\
        );

    \I__1145\ : Span4Mux_v
    port map (
            O => \N__5456\,
            I => \N__5447\
        );

    \I__1144\ : SRMux
    port map (
            O => \N__5455\,
            I => \N__5444\
        );

    \I__1143\ : Span4Mux_h
    port map (
            O => \N__5452\,
            I => \N__5441\
        );

    \I__1142\ : Span4Mux_h
    port map (
            O => \N__5447\,
            I => \N__5438\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__5444\,
            I => \N__5435\
        );

    \I__1140\ : Odrv4
    port map (
            O => \N__5441\,
            I => n1895
        );

    \I__1139\ : Odrv4
    port map (
            O => \N__5438\,
            I => n1895
        );

    \I__1138\ : Odrv12
    port map (
            O => \N__5435\,
            I => n1895
        );

    \I__1137\ : IoInMux
    port map (
            O => \N__5428\,
            I => \N__5425\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__5425\,
            I => \N__5422\
        );

    \I__1135\ : IoSpan4Mux
    port map (
            O => \N__5422\,
            I => \N__5419\
        );

    \I__1134\ : Span4Mux_s3_h
    port map (
            O => \N__5419\,
            I => \N__5416\
        );

    \I__1133\ : Sp12to4
    port map (
            O => \N__5416\,
            I => \N__5413\
        );

    \I__1132\ : Odrv12
    port map (
            O => \N__5413\,
            I => sda_out
        );

    \I__1131\ : IoInMux
    port map (
            O => \N__5410\,
            I => \N__5407\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__5407\,
            I => \N__5404\
        );

    \I__1129\ : Span4Mux_s3_h
    port map (
            O => \N__5404\,
            I => \N__5401\
        );

    \I__1128\ : Span4Mux_h
    port map (
            O => \N__5401\,
            I => \N__5397\
        );

    \I__1127\ : InMux
    port map (
            O => \N__5400\,
            I => \N__5394\
        );

    \I__1126\ : Odrv4
    port map (
            O => \N__5397\,
            I => sda_enable
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__5394\,
            I => sda_enable
        );

    \I__1124\ : CEMux
    port map (
            O => \N__5389\,
            I => \N__5386\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__5386\,
            I => \eeprom.i2c.n1152\
        );

    \I__1122\ : SRMux
    port map (
            O => \N__5383\,
            I => \N__5380\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__5380\,
            I => \N__5377\
        );

    \I__1120\ : Span4Mux_v
    port map (
            O => \N__5377\,
            I => \N__5374\
        );

    \I__1119\ : Span4Mux_h
    port map (
            O => \N__5374\,
            I => \N__5371\
        );

    \I__1118\ : Odrv4
    port map (
            O => \N__5371\,
            I => \eeprom.i2c.n1932\
        );

    \I__1117\ : InMux
    port map (
            O => \N__5368\,
            I => \N__5365\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__5365\,
            I => \N__5362\
        );

    \I__1115\ : Span4Mux_h
    port map (
            O => \N__5362\,
            I => \N__5358\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5361\,
            I => \N__5355\
        );

    \I__1113\ : Odrv4
    port map (
            O => \N__5358\,
            I => \eeprom.i2c.n11_adj_378\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__5355\,
            I => \eeprom.i2c.n11_adj_378\
        );

    \I__1111\ : InMux
    port map (
            O => \N__5350\,
            I => \N__5347\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__5347\,
            I => \eeprom.i2c.n13\
        );

    \I__1109\ : InMux
    port map (
            O => \N__5344\,
            I => \N__5341\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__5341\,
            I => \eeprom.i2c.n11_adj_381\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5338\,
            I => \N__5334\
        );

    \I__1106\ : InMux
    port map (
            O => \N__5337\,
            I => \N__5331\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__5334\,
            I => delay_counter_20
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__5331\,
            I => delay_counter_20
        );

    \I__1103\ : InMux
    port map (
            O => \N__5326\,
            I => n2652
        );

    \I__1102\ : InMux
    port map (
            O => \N__5323\,
            I => \N__5319\
        );

    \I__1101\ : InMux
    port map (
            O => \N__5322\,
            I => \N__5316\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__5319\,
            I => delay_counter_21
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__5316\,
            I => delay_counter_21
        );

    \I__1098\ : InMux
    port map (
            O => \N__5311\,
            I => n2653
        );

    \I__1097\ : InMux
    port map (
            O => \N__5308\,
            I => \N__5304\
        );

    \I__1096\ : InMux
    port map (
            O => \N__5307\,
            I => \N__5301\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__5304\,
            I => delay_counter_22
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__5301\,
            I => delay_counter_22
        );

    \I__1093\ : InMux
    port map (
            O => \N__5296\,
            I => n2654
        );

    \I__1092\ : InMux
    port map (
            O => \N__5293\,
            I => \N__5289\
        );

    \I__1091\ : InMux
    port map (
            O => \N__5292\,
            I => \N__5286\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__5289\,
            I => delay_counter_23
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__5286\,
            I => delay_counter_23
        );

    \I__1088\ : InMux
    port map (
            O => \N__5281\,
            I => n2655
        );

    \I__1087\ : InMux
    port map (
            O => \N__5278\,
            I => \N__5274\
        );

    \I__1086\ : InMux
    port map (
            O => \N__5277\,
            I => \N__5271\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__5274\,
            I => \N__5268\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__5271\,
            I => delay_counter_24
        );

    \I__1083\ : Odrv4
    port map (
            O => \N__5268\,
            I => delay_counter_24
        );

    \I__1082\ : InMux
    port map (
            O => \N__5263\,
            I => \bfn_23_16_0_\
        );

    \I__1081\ : CascadeMux
    port map (
            O => \N__5260\,
            I => \N__5256\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5259\,
            I => \N__5253\
        );

    \I__1079\ : InMux
    port map (
            O => \N__5256\,
            I => \N__5250\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__5253\,
            I => delay_counter_25
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__5250\,
            I => delay_counter_25
        );

    \I__1076\ : InMux
    port map (
            O => \N__5245\,
            I => n2657
        );

    \I__1075\ : InMux
    port map (
            O => \N__5242\,
            I => \N__5238\
        );

    \I__1074\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5235\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__5238\,
            I => \N__5232\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__5235\,
            I => delay_counter_26
        );

    \I__1071\ : Odrv4
    port map (
            O => \N__5232\,
            I => delay_counter_26
        );

    \I__1070\ : InMux
    port map (
            O => \N__5227\,
            I => n2658
        );

    \I__1069\ : InMux
    port map (
            O => \N__5224\,
            I => \N__5220\
        );

    \I__1068\ : InMux
    port map (
            O => \N__5223\,
            I => \N__5217\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__5220\,
            I => delay_counter_27
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__5217\,
            I => delay_counter_27
        );

    \I__1065\ : InMux
    port map (
            O => \N__5212\,
            I => n2659
        );

    \I__1064\ : InMux
    port map (
            O => \N__5209\,
            I => \N__5205\
        );

    \I__1063\ : InMux
    port map (
            O => \N__5208\,
            I => \N__5202\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__5205\,
            I => delay_counter_11
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__5202\,
            I => delay_counter_11
        );

    \I__1060\ : InMux
    port map (
            O => \N__5197\,
            I => n2643
        );

    \I__1059\ : InMux
    port map (
            O => \N__5194\,
            I => \N__5190\
        );

    \I__1058\ : InMux
    port map (
            O => \N__5193\,
            I => \N__5187\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__5190\,
            I => delay_counter_12
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__5187\,
            I => delay_counter_12
        );

    \I__1055\ : InMux
    port map (
            O => \N__5182\,
            I => n2644
        );

    \I__1054\ : InMux
    port map (
            O => \N__5179\,
            I => \N__5175\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5178\,
            I => \N__5172\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__5175\,
            I => delay_counter_13
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__5172\,
            I => delay_counter_13
        );

    \I__1050\ : InMux
    port map (
            O => \N__5167\,
            I => n2645
        );

    \I__1049\ : InMux
    port map (
            O => \N__5164\,
            I => \N__5160\
        );

    \I__1048\ : InMux
    port map (
            O => \N__5163\,
            I => \N__5157\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__5160\,
            I => delay_counter_14
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__5157\,
            I => delay_counter_14
        );

    \I__1045\ : InMux
    port map (
            O => \N__5152\,
            I => n2646
        );

    \I__1044\ : CascadeMux
    port map (
            O => \N__5149\,
            I => \N__5145\
        );

    \I__1043\ : InMux
    port map (
            O => \N__5148\,
            I => \N__5142\
        );

    \I__1042\ : InMux
    port map (
            O => \N__5145\,
            I => \N__5139\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__5142\,
            I => delay_counter_15
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__5139\,
            I => delay_counter_15
        );

    \I__1039\ : InMux
    port map (
            O => \N__5134\,
            I => n2647
        );

    \I__1038\ : InMux
    port map (
            O => \N__5131\,
            I => \N__5127\
        );

    \I__1037\ : InMux
    port map (
            O => \N__5130\,
            I => \N__5124\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__5127\,
            I => delay_counter_16
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__5124\,
            I => delay_counter_16
        );

    \I__1034\ : InMux
    port map (
            O => \N__5119\,
            I => \bfn_23_15_0_\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5116\,
            I => \N__5112\
        );

    \I__1032\ : InMux
    port map (
            O => \N__5115\,
            I => \N__5109\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__5112\,
            I => delay_counter_17
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__5109\,
            I => delay_counter_17
        );

    \I__1029\ : InMux
    port map (
            O => \N__5104\,
            I => n2649
        );

    \I__1028\ : InMux
    port map (
            O => \N__5101\,
            I => \N__5097\
        );

    \I__1027\ : InMux
    port map (
            O => \N__5100\,
            I => \N__5094\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__5097\,
            I => delay_counter_18
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__5094\,
            I => delay_counter_18
        );

    \I__1024\ : InMux
    port map (
            O => \N__5089\,
            I => n2650
        );

    \I__1023\ : InMux
    port map (
            O => \N__5086\,
            I => \N__5082\
        );

    \I__1022\ : InMux
    port map (
            O => \N__5085\,
            I => \N__5079\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__5082\,
            I => delay_counter_19
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__5079\,
            I => delay_counter_19
        );

    \I__1019\ : InMux
    port map (
            O => \N__5074\,
            I => n2651
        );

    \I__1018\ : CascadeMux
    port map (
            O => \N__5071\,
            I => \N__5067\
        );

    \I__1017\ : InMux
    port map (
            O => \N__5070\,
            I => \N__5064\
        );

    \I__1016\ : InMux
    port map (
            O => \N__5067\,
            I => \N__5061\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__5064\,
            I => delay_counter_3
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__5061\,
            I => delay_counter_3
        );

    \I__1013\ : InMux
    port map (
            O => \N__5056\,
            I => n2635
        );

    \I__1012\ : CascadeMux
    port map (
            O => \N__5053\,
            I => \N__5049\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5052\,
            I => \N__5046\
        );

    \I__1010\ : InMux
    port map (
            O => \N__5049\,
            I => \N__5043\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__5046\,
            I => delay_counter_4
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5043\,
            I => delay_counter_4
        );

    \I__1007\ : InMux
    port map (
            O => \N__5038\,
            I => n2636
        );

    \I__1006\ : InMux
    port map (
            O => \N__5035\,
            I => \N__5031\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5034\,
            I => \N__5028\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__5031\,
            I => \N__5025\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5028\,
            I => delay_counter_5
        );

    \I__1002\ : Odrv4
    port map (
            O => \N__5025\,
            I => delay_counter_5
        );

    \I__1001\ : InMux
    port map (
            O => \N__5020\,
            I => n2637
        );

    \I__1000\ : InMux
    port map (
            O => \N__5017\,
            I => \N__5013\
        );

    \I__999\ : InMux
    port map (
            O => \N__5016\,
            I => \N__5010\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__5013\,
            I => delay_counter_6
        );

    \I__997\ : LocalMux
    port map (
            O => \N__5010\,
            I => delay_counter_6
        );

    \I__996\ : InMux
    port map (
            O => \N__5005\,
            I => n2638
        );

    \I__995\ : InMux
    port map (
            O => \N__5002\,
            I => \N__4998\
        );

    \I__994\ : InMux
    port map (
            O => \N__5001\,
            I => \N__4995\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__4998\,
            I => delay_counter_7
        );

    \I__992\ : LocalMux
    port map (
            O => \N__4995\,
            I => delay_counter_7
        );

    \I__991\ : InMux
    port map (
            O => \N__4990\,
            I => n2639
        );

    \I__990\ : InMux
    port map (
            O => \N__4987\,
            I => \N__4983\
        );

    \I__989\ : InMux
    port map (
            O => \N__4986\,
            I => \N__4980\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__4983\,
            I => delay_counter_8
        );

    \I__987\ : LocalMux
    port map (
            O => \N__4980\,
            I => delay_counter_8
        );

    \I__986\ : InMux
    port map (
            O => \N__4975\,
            I => \bfn_23_14_0_\
        );

    \I__985\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4968\
        );

    \I__984\ : InMux
    port map (
            O => \N__4971\,
            I => \N__4965\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__4968\,
            I => delay_counter_9
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4965\,
            I => delay_counter_9
        );

    \I__981\ : InMux
    port map (
            O => \N__4960\,
            I => n2641
        );

    \I__980\ : InMux
    port map (
            O => \N__4957\,
            I => \N__4953\
        );

    \I__979\ : InMux
    port map (
            O => \N__4956\,
            I => \N__4950\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__4953\,
            I => delay_counter_10
        );

    \I__977\ : LocalMux
    port map (
            O => \N__4950\,
            I => delay_counter_10
        );

    \I__976\ : InMux
    port map (
            O => \N__4945\,
            I => n2642
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__4942\,
            I => \N__4939\
        );

    \I__974\ : InMux
    port map (
            O => \N__4939\,
            I => \N__4936\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__4936\,
            I => \N__4933\
        );

    \I__972\ : Odrv4
    port map (
            O => \N__4933\,
            I => n2434
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__4930\,
            I => \n2434_cascade_\
        );

    \I__970\ : InMux
    port map (
            O => \N__4927\,
            I => \N__4924\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__4924\,
            I => \N__4921\
        );

    \I__968\ : Odrv4
    port map (
            O => \N__4921\,
            I => n2958
        );

    \I__967\ : InMux
    port map (
            O => \N__4918\,
            I => \N__4911\
        );

    \I__966\ : InMux
    port map (
            O => \N__4917\,
            I => \N__4907\
        );

    \I__965\ : InMux
    port map (
            O => \N__4916\,
            I => \N__4900\
        );

    \I__964\ : InMux
    port map (
            O => \N__4915\,
            I => \N__4900\
        );

    \I__963\ : InMux
    port map (
            O => \N__4914\,
            I => \N__4900\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__4911\,
            I => \N__4897\
        );

    \I__961\ : InMux
    port map (
            O => \N__4910\,
            I => \N__4894\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4907\,
            I => \eeprom.i2c.counter_1\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4900\,
            I => \eeprom.i2c.counter_1\
        );

    \I__958\ : Odrv4
    port map (
            O => \N__4897\,
            I => \eeprom.i2c.counter_1\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__4894\,
            I => \eeprom.i2c.counter_1\
        );

    \I__956\ : InMux
    port map (
            O => \N__4885\,
            I => \N__4881\
        );

    \I__955\ : InMux
    port map (
            O => \N__4884\,
            I => \N__4878\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4881\,
            I => \N__4872\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4878\,
            I => \N__4869\
        );

    \I__952\ : InMux
    port map (
            O => \N__4877\,
            I => \N__4866\
        );

    \I__951\ : InMux
    port map (
            O => \N__4876\,
            I => \N__4863\
        );

    \I__950\ : InMux
    port map (
            O => \N__4875\,
            I => \N__4860\
        );

    \I__949\ : Sp12to4
    port map (
            O => \N__4872\,
            I => \N__4853\
        );

    \I__948\ : Sp12to4
    port map (
            O => \N__4869\,
            I => \N__4853\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4866\,
            I => \N__4853\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4863\,
            I => \eeprom.i2c.counter_0\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4860\,
            I => \eeprom.i2c.counter_0\
        );

    \I__944\ : Odrv12
    port map (
            O => \N__4853\,
            I => \eeprom.i2c.counter_0\
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__4846\,
            I => \N__4841\
        );

    \I__942\ : CascadeMux
    port map (
            O => \N__4845\,
            I => \N__4837\
        );

    \I__941\ : InMux
    port map (
            O => \N__4844\,
            I => \N__4832\
        );

    \I__940\ : InMux
    port map (
            O => \N__4841\,
            I => \N__4829\
        );

    \I__939\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4822\
        );

    \I__938\ : InMux
    port map (
            O => \N__4837\,
            I => \N__4822\
        );

    \I__937\ : InMux
    port map (
            O => \N__4836\,
            I => \N__4822\
        );

    \I__936\ : InMux
    port map (
            O => \N__4835\,
            I => \N__4819\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__4832\,
            I => \N__4816\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__4829\,
            I => \eeprom.i2c.counter_2\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4822\,
            I => \eeprom.i2c.counter_2\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4819\,
            I => \eeprom.i2c.counter_2\
        );

    \I__931\ : Odrv4
    port map (
            O => \N__4816\,
            I => \eeprom.i2c.counter_2\
        );

    \I__930\ : CascadeMux
    port map (
            O => \N__4807\,
            I => \eeprom.i2c.n2967_cascade_\
        );

    \I__929\ : InMux
    port map (
            O => \N__4804\,
            I => \N__4801\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__4801\,
            I => \N__4798\
        );

    \I__927\ : Span4Mux_v
    port map (
            O => \N__4798\,
            I => \N__4794\
        );

    \I__926\ : InMux
    port map (
            O => \N__4797\,
            I => \N__4791\
        );

    \I__925\ : Odrv4
    port map (
            O => \N__4794\,
            I => rw
        );

    \I__924\ : LocalMux
    port map (
            O => \N__4791\,
            I => rw
        );

    \I__923\ : InMux
    port map (
            O => \N__4786\,
            I => \N__4781\
        );

    \I__922\ : InMux
    port map (
            O => \N__4785\,
            I => \N__4776\
        );

    \I__921\ : InMux
    port map (
            O => \N__4784\,
            I => \N__4776\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4781\,
            I => saved_addr_0
        );

    \I__919\ : LocalMux
    port map (
            O => \N__4776\,
            I => saved_addr_0
        );

    \I__918\ : InMux
    port map (
            O => \N__4771\,
            I => \N__4767\
        );

    \I__917\ : InMux
    port map (
            O => \N__4770\,
            I => \N__4764\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4767\,
            I => \N__4761\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__4764\,
            I => \N__4758\
        );

    \I__914\ : Odrv4
    port map (
            O => \N__4761\,
            I => \eeprom.enable\
        );

    \I__913\ : Odrv12
    port map (
            O => \N__4758\,
            I => \eeprom.enable\
        );

    \I__912\ : InMux
    port map (
            O => \N__4753\,
            I => \N__4749\
        );

    \I__911\ : InMux
    port map (
            O => \N__4752\,
            I => \N__4746\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__4749\,
            I => delay_counter_0
        );

    \I__909\ : LocalMux
    port map (
            O => \N__4746\,
            I => delay_counter_0
        );

    \I__908\ : InMux
    port map (
            O => \N__4741\,
            I => \bfn_23_13_0_\
        );

    \I__907\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4734\
        );

    \I__906\ : InMux
    port map (
            O => \N__4737\,
            I => \N__4731\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__4734\,
            I => delay_counter_1
        );

    \I__904\ : LocalMux
    port map (
            O => \N__4731\,
            I => delay_counter_1
        );

    \I__903\ : InMux
    port map (
            O => \N__4726\,
            I => n2633
        );

    \I__902\ : InMux
    port map (
            O => \N__4723\,
            I => \N__4719\
        );

    \I__901\ : InMux
    port map (
            O => \N__4722\,
            I => \N__4716\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4719\,
            I => \N__4713\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__4716\,
            I => delay_counter_2
        );

    \I__898\ : Odrv4
    port map (
            O => \N__4713\,
            I => delay_counter_2
        );

    \I__897\ : InMux
    port map (
            O => \N__4708\,
            I => n2634
        );

    \I__896\ : CascadeMux
    port map (
            O => \N__4705\,
            I => \eeprom.i2c.n1739_cascade_\
        );

    \I__895\ : InMux
    port map (
            O => \N__4702\,
            I => \N__4698\
        );

    \I__894\ : InMux
    port map (
            O => \N__4701\,
            I => \N__4695\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4698\,
            I => \eeprom.i2c.n1054\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4695\,
            I => \eeprom.i2c.n1054\
        );

    \I__891\ : InMux
    port map (
            O => \N__4690\,
            I => \N__4684\
        );

    \I__890\ : InMux
    port map (
            O => \N__4689\,
            I => \N__4684\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__4684\,
            I => n2414
        );

    \I__888\ : CascadeMux
    port map (
            O => \N__4681\,
            I => \n1061_cascade_\
        );

    \I__887\ : InMux
    port map (
            O => \N__4678\,
            I => \N__4672\
        );

    \I__886\ : InMux
    port map (
            O => \N__4677\,
            I => \N__4672\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4672\,
            I => \N__4669\
        );

    \I__884\ : Odrv12
    port map (
            O => \N__4669\,
            I => \eeprom.i2c.n2869\
        );

    \I__883\ : CascadeMux
    port map (
            O => \N__4666\,
            I => \N__4660\
        );

    \I__882\ : InMux
    port map (
            O => \N__4665\,
            I => \N__4653\
        );

    \I__881\ : InMux
    port map (
            O => \N__4664\,
            I => \N__4644\
        );

    \I__880\ : InMux
    port map (
            O => \N__4663\,
            I => \N__4644\
        );

    \I__879\ : InMux
    port map (
            O => \N__4660\,
            I => \N__4644\
        );

    \I__878\ : InMux
    port map (
            O => \N__4659\,
            I => \N__4644\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__4658\,
            I => \N__4640\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__4657\,
            I => \N__4636\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__4656\,
            I => \N__4632\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__4653\,
            I => \N__4626\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__4644\,
            I => \N__4626\
        );

    \I__872\ : InMux
    port map (
            O => \N__4643\,
            I => \N__4623\
        );

    \I__871\ : InMux
    port map (
            O => \N__4640\,
            I => \N__4620\
        );

    \I__870\ : CascadeMux
    port map (
            O => \N__4639\,
            I => \N__4616\
        );

    \I__869\ : InMux
    port map (
            O => \N__4636\,
            I => \N__4613\
        );

    \I__868\ : InMux
    port map (
            O => \N__4635\,
            I => \N__4608\
        );

    \I__867\ : InMux
    port map (
            O => \N__4632\,
            I => \N__4608\
        );

    \I__866\ : InMux
    port map (
            O => \N__4631\,
            I => \N__4605\
        );

    \I__865\ : Span4Mux_h
    port map (
            O => \N__4626\,
            I => \N__4598\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4623\,
            I => \N__4598\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__4620\,
            I => \N__4598\
        );

    \I__862\ : InMux
    port map (
            O => \N__4619\,
            I => \N__4593\
        );

    \I__861\ : InMux
    port map (
            O => \N__4616\,
            I => \N__4593\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4613\,
            I => \N__4586\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__4608\,
            I => \N__4586\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__4605\,
            I => \N__4586\
        );

    \I__857\ : Span4Mux_v
    port map (
            O => \N__4598\,
            I => \N__4581\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__4593\,
            I => \N__4581\
        );

    \I__855\ : Span4Mux_v
    port map (
            O => \N__4586\,
            I => \N__4578\
        );

    \I__854\ : Span4Mux_v
    port map (
            O => \N__4581\,
            I => \N__4575\
        );

    \I__853\ : Span4Mux_v
    port map (
            O => \N__4578\,
            I => \N__4572\
        );

    \I__852\ : Span4Mux_h
    port map (
            O => \N__4575\,
            I => \N__4569\
        );

    \I__851\ : Sp12to4
    port map (
            O => \N__4572\,
            I => \N__4566\
        );

    \I__850\ : Span4Mux_h
    port map (
            O => \N__4569\,
            I => \N__4563\
        );

    \I__849\ : Odrv12
    port map (
            O => \N__4566\,
            I => \state_7_N_289_3\
        );

    \I__848\ : Odrv4
    port map (
            O => \N__4563\,
            I => \state_7_N_289_3\
        );

    \I__847\ : CEMux
    port map (
            O => \N__4558\,
            I => \N__4555\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4555\,
            I => \N__4550\
        );

    \I__845\ : CEMux
    port map (
            O => \N__4554\,
            I => \N__4547\
        );

    \I__844\ : CEMux
    port map (
            O => \N__4553\,
            I => \N__4544\
        );

    \I__843\ : Span4Mux_v
    port map (
            O => \N__4550\,
            I => \N__4540\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4547\,
            I => \N__4535\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__4544\,
            I => \N__4535\
        );

    \I__840\ : CascadeMux
    port map (
            O => \N__4543\,
            I => \N__4531\
        );

    \I__839\ : Span4Mux_h
    port map (
            O => \N__4540\,
            I => \N__4527\
        );

    \I__838\ : Span4Mux_v
    port map (
            O => \N__4535\,
            I => \N__4524\
        );

    \I__837\ : InMux
    port map (
            O => \N__4534\,
            I => \N__4521\
        );

    \I__836\ : InMux
    port map (
            O => \N__4531\,
            I => \N__4518\
        );

    \I__835\ : InMux
    port map (
            O => \N__4530\,
            I => \N__4515\
        );

    \I__834\ : Odrv4
    port map (
            O => \N__4527\,
            I => n1061
        );

    \I__833\ : Odrv4
    port map (
            O => \N__4524\,
            I => n1061
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4521\,
            I => n1061
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4518\,
            I => n1061
        );

    \I__830\ : LocalMux
    port map (
            O => \N__4515\,
            I => n1061
        );

    \I__829\ : SRMux
    port map (
            O => \N__4504\,
            I => \N__4501\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__4501\,
            I => \N__4498\
        );

    \I__827\ : Span4Mux_h
    port map (
            O => \N__4498\,
            I => \N__4495\
        );

    \I__826\ : Odrv4
    port map (
            O => \N__4495\,
            I => \eeprom.i2c.n2479\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__4492\,
            I => \N__4489\
        );

    \I__824\ : InMux
    port map (
            O => \N__4489\,
            I => \N__4486\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__4486\,
            I => \eeprom.i2c.n10\
        );

    \I__822\ : InMux
    port map (
            O => \N__4483\,
            I => \N__4480\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4480\,
            I => \N__4477\
        );

    \I__820\ : Odrv4
    port map (
            O => \N__4477\,
            I => \eeprom.i2c.n7\
        );

    \I__819\ : InMux
    port map (
            O => \N__4474\,
            I => \N__4468\
        );

    \I__818\ : CascadeMux
    port map (
            O => \N__4473\,
            I => \N__4463\
        );

    \I__817\ : CascadeMux
    port map (
            O => \N__4472\,
            I => \N__4459\
        );

    \I__816\ : CascadeMux
    port map (
            O => \N__4471\,
            I => \N__4455\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4468\,
            I => \N__4452\
        );

    \I__814\ : InMux
    port map (
            O => \N__4467\,
            I => \N__4437\
        );

    \I__813\ : InMux
    port map (
            O => \N__4466\,
            I => \N__4437\
        );

    \I__812\ : InMux
    port map (
            O => \N__4463\,
            I => \N__4437\
        );

    \I__811\ : InMux
    port map (
            O => \N__4462\,
            I => \N__4437\
        );

    \I__810\ : InMux
    port map (
            O => \N__4459\,
            I => \N__4437\
        );

    \I__809\ : InMux
    port map (
            O => \N__4458\,
            I => \N__4437\
        );

    \I__808\ : InMux
    port map (
            O => \N__4455\,
            I => \N__4437\
        );

    \I__807\ : Odrv4
    port map (
            O => \N__4452\,
            I => \CONSTANT_ONE_NET\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4437\,
            I => \CONSTANT_ONE_NET\
        );

    \I__805\ : CascadeMux
    port map (
            O => \N__4432\,
            I => \n22_cascade_\
        );

    \I__804\ : CascadeMux
    port map (
            O => \N__4429\,
            I => \n25_cascade_\
        );

    \I__803\ : InMux
    port map (
            O => \N__4426\,
            I => \N__4421\
        );

    \I__802\ : InMux
    port map (
            O => \N__4425\,
            I => \N__4416\
        );

    \I__801\ : InMux
    port map (
            O => \N__4424\,
            I => \N__4416\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4421\,
            I => n104
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4416\,
            I => n104
        );

    \I__798\ : InMux
    port map (
            O => \N__4411\,
            I => \N__4408\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4408\,
            I => n24
        );

    \I__796\ : InMux
    port map (
            O => \N__4405\,
            I => \N__4402\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__4402\,
            I => \N__4399\
        );

    \I__794\ : Odrv4
    port map (
            O => \N__4399\,
            I => n23
        );

    \I__793\ : CEMux
    port map (
            O => \N__4396\,
            I => \N__4392\
        );

    \I__792\ : CEMux
    port map (
            O => \N__4395\,
            I => \N__4389\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__4392\,
            I => \N__4386\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__4389\,
            I => \N__4383\
        );

    \I__789\ : Odrv12
    port map (
            O => \N__4386\,
            I => \eeprom.i2c.n1837\
        );

    \I__788\ : Odrv12
    port map (
            O => \N__4383\,
            I => \eeprom.i2c.n1837\
        );

    \I__787\ : SRMux
    port map (
            O => \N__4378\,
            I => \N__4374\
        );

    \I__786\ : SRMux
    port map (
            O => \N__4377\,
            I => \N__4371\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__4374\,
            I => \N__4368\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__4371\,
            I => \N__4365\
        );

    \I__783\ : Odrv12
    port map (
            O => \N__4368\,
            I => \eeprom.i2c.n1928\
        );

    \I__782\ : Odrv12
    port map (
            O => \N__4365\,
            I => \eeprom.i2c.n1928\
        );

    \I__781\ : InMux
    port map (
            O => \N__4360\,
            I => \N__4356\
        );

    \I__780\ : InMux
    port map (
            O => \N__4359\,
            I => \N__4353\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__4356\,
            I => \eeprom.i2c.n37\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__4353\,
            I => \eeprom.i2c.n37\
        );

    \I__777\ : InMux
    port map (
            O => \N__4348\,
            I => \N__4344\
        );

    \I__776\ : InMux
    port map (
            O => \N__4347\,
            I => \N__4341\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4344\,
            I => \eeprom.i2c.n33\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__4341\,
            I => \eeprom.i2c.n33\
        );

    \I__773\ : InMux
    port map (
            O => \N__4336\,
            I => \N__4331\
        );

    \I__772\ : InMux
    port map (
            O => \N__4335\,
            I => \N__4328\
        );

    \I__771\ : InMux
    port map (
            O => \N__4334\,
            I => \N__4325\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__4331\,
            I => \N__4322\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__4328\,
            I => \eeprom.i2c.n9\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__4325\,
            I => \eeprom.i2c.n9\
        );

    \I__767\ : Odrv12
    port map (
            O => \N__4322\,
            I => \eeprom.i2c.n9\
        );

    \I__766\ : InMux
    port map (
            O => \N__4315\,
            I => \N__4312\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__4312\,
            I => \N__4307\
        );

    \I__764\ : InMux
    port map (
            O => \N__4311\,
            I => \N__4302\
        );

    \I__763\ : InMux
    port map (
            O => \N__4310\,
            I => \N__4302\
        );

    \I__762\ : Odrv4
    port map (
            O => \N__4307\,
            I => \eeprom.i2c.n10_adj_384\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__4302\,
            I => \eeprom.i2c.n10_adj_384\
        );

    \I__760\ : InMux
    port map (
            O => \N__4297\,
            I => \N__4291\
        );

    \I__759\ : InMux
    port map (
            O => \N__4296\,
            I => \N__4291\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__4291\,
            I => n4_adj_393
        );

    \I__757\ : InMux
    port map (
            O => \N__4288\,
            I => \N__4285\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__4285\,
            I => n14
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__4282\,
            I => \n13_cascade_\
        );

    \I__754\ : CascadeMux
    port map (
            O => \N__4279\,
            I => \n18_cascade_\
        );

    \I__753\ : CascadeMux
    port map (
            O => \N__4276\,
            I => \n2935_cascade_\
        );

    \I__752\ : InMux
    port map (
            O => \N__4273\,
            I => \N__4270\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4270\,
            I => n2939
        );

    \I__750\ : CascadeMux
    port map (
            O => \N__4267\,
            I => \n36_cascade_\
        );

    \I__749\ : InMux
    port map (
            O => \N__4264\,
            I => \eeprom.i2c.n2669\
        );

    \I__748\ : InMux
    port map (
            O => \N__4261\,
            I => \eeprom.i2c.n2670\
        );

    \I__747\ : InMux
    port map (
            O => \N__4258\,
            I => \N__4254\
        );

    \I__746\ : InMux
    port map (
            O => \N__4257\,
            I => \N__4251\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__4254\,
            I => \N__4248\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__4251\,
            I => \eeprom.i2c.counter_7\
        );

    \I__743\ : Odrv4
    port map (
            O => \N__4248\,
            I => \eeprom.i2c.counter_7\
        );

    \I__742\ : InMux
    port map (
            O => \N__4243\,
            I => \N__4240\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__4240\,
            I => n14_adj_395
        );

    \I__740\ : CascadeMux
    port map (
            O => \N__4237\,
            I => \n4_adj_394_cascade_\
        );

    \I__739\ : InMux
    port map (
            O => \N__4234\,
            I => \N__4228\
        );

    \I__738\ : InMux
    port map (
            O => \N__4233\,
            I => \N__4228\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__4228\,
            I => data_4
        );

    \I__736\ : InMux
    port map (
            O => \N__4225\,
            I => \N__4219\
        );

    \I__735\ : InMux
    port map (
            O => \N__4224\,
            I => \N__4214\
        );

    \I__734\ : InMux
    port map (
            O => \N__4223\,
            I => \N__4214\
        );

    \I__733\ : InMux
    port map (
            O => \N__4222\,
            I => \N__4211\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__4219\,
            I => \N__4206\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4214\,
            I => \N__4206\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__4211\,
            I => n1717
        );

    \I__729\ : Odrv4
    port map (
            O => \N__4206\,
            I => n1717
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__4201\,
            I => \N__4197\
        );

    \I__727\ : InMux
    port map (
            O => \N__4200\,
            I => \N__4192\
        );

    \I__726\ : InMux
    port map (
            O => \N__4197\,
            I => \N__4192\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__4192\,
            I => data_6
        );

    \I__724\ : InMux
    port map (
            O => \N__4189\,
            I => \N__4186\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__4186\,
            I => n2424
        );

    \I__722\ : CascadeMux
    port map (
            O => \N__4183\,
            I => \n2424_cascade_\
        );

    \I__721\ : InMux
    port map (
            O => \N__4180\,
            I => \N__4174\
        );

    \I__720\ : InMux
    port map (
            O => \N__4179\,
            I => \N__4174\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__4174\,
            I => data_7
        );

    \I__718\ : InMux
    port map (
            O => \N__4171\,
            I => \N__4168\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__4168\,
            I => n4_adj_394
        );

    \I__716\ : InMux
    port map (
            O => \N__4165\,
            I => \N__4159\
        );

    \I__715\ : InMux
    port map (
            O => \N__4164\,
            I => \N__4154\
        );

    \I__714\ : InMux
    port map (
            O => \N__4163\,
            I => \N__4154\
        );

    \I__713\ : InMux
    port map (
            O => \N__4162\,
            I => \N__4151\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__4159\,
            I => n1722
        );

    \I__711\ : LocalMux
    port map (
            O => \N__4154\,
            I => n1722
        );

    \I__710\ : LocalMux
    port map (
            O => \N__4151\,
            I => n1722
        );

    \I__709\ : CascadeMux
    port map (
            O => \N__4144\,
            I => \N__4141\
        );

    \I__708\ : InMux
    port map (
            O => \N__4141\,
            I => \N__4135\
        );

    \I__707\ : InMux
    port map (
            O => \N__4140\,
            I => \N__4135\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__4135\,
            I => data_5
        );

    \I__705\ : CascadeMux
    port map (
            O => \N__4132\,
            I => \eeprom.i2c.n15_cascade_\
        );

    \I__704\ : SRMux
    port map (
            O => \N__4129\,
            I => \N__4126\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__4126\,
            I => \N__4123\
        );

    \I__702\ : Span4Mux_v
    port map (
            O => \N__4123\,
            I => \N__4120\
        );

    \I__701\ : Odrv4
    port map (
            O => \N__4120\,
            I => \eeprom.i2c.n2454\
        );

    \I__700\ : InMux
    port map (
            O => \N__4117\,
            I => \N__4113\
        );

    \I__699\ : InMux
    port map (
            O => \N__4116\,
            I => \N__4110\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__4113\,
            I => \eeprom.i2c.n15\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__4110\,
            I => \eeprom.i2c.n15\
        );

    \I__696\ : InMux
    port map (
            O => \N__4105\,
            I => \eeprom.i2c.n2664\
        );

    \I__695\ : InMux
    port map (
            O => \N__4102\,
            I => \eeprom.i2c.n2665\
        );

    \I__694\ : InMux
    port map (
            O => \N__4099\,
            I => \N__4095\
        );

    \I__693\ : InMux
    port map (
            O => \N__4098\,
            I => \N__4092\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__4095\,
            I => \N__4089\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__4092\,
            I => \eeprom.i2c.counter_3\
        );

    \I__690\ : Odrv4
    port map (
            O => \N__4089\,
            I => \eeprom.i2c.counter_3\
        );

    \I__689\ : InMux
    port map (
            O => \N__4084\,
            I => \eeprom.i2c.n2666\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__4081\,
            I => \N__4077\
        );

    \I__687\ : InMux
    port map (
            O => \N__4080\,
            I => \N__4074\
        );

    \I__686\ : InMux
    port map (
            O => \N__4077\,
            I => \N__4071\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__4074\,
            I => \N__4068\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__4071\,
            I => \eeprom.i2c.counter_4\
        );

    \I__683\ : Odrv4
    port map (
            O => \N__4068\,
            I => \eeprom.i2c.counter_4\
        );

    \I__682\ : InMux
    port map (
            O => \N__4063\,
            I => \eeprom.i2c.n2667\
        );

    \I__681\ : InMux
    port map (
            O => \N__4060\,
            I => \N__4056\
        );

    \I__680\ : InMux
    port map (
            O => \N__4059\,
            I => \N__4053\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__4056\,
            I => \N__4050\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__4053\,
            I => \eeprom.i2c.counter_5\
        );

    \I__677\ : Odrv4
    port map (
            O => \N__4050\,
            I => \eeprom.i2c.counter_5\
        );

    \I__676\ : InMux
    port map (
            O => \N__4045\,
            I => \eeprom.i2c.n2668\
        );

    \I__675\ : CascadeMux
    port map (
            O => \N__4042\,
            I => \N__4038\
        );

    \I__674\ : InMux
    port map (
            O => \N__4041\,
            I => \N__4035\
        );

    \I__673\ : InMux
    port map (
            O => \N__4038\,
            I => \N__4032\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__4035\,
            I => \N__4029\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4032\,
            I => \eeprom.i2c.counter_6\
        );

    \I__670\ : Odrv12
    port map (
            O => \N__4029\,
            I => \eeprom.i2c.counter_6\
        );

    \I__669\ : SRMux
    port map (
            O => \N__4024\,
            I => \N__4021\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__4021\,
            I => \N__4018\
        );

    \I__667\ : Odrv4
    port map (
            O => \N__4018\,
            I => \eeprom.i2c.n2927\
        );

    \I__666\ : InMux
    port map (
            O => \N__4015\,
            I => \N__4009\
        );

    \I__665\ : InMux
    port map (
            O => \N__4014\,
            I => \N__4009\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__4009\,
            I => \N__4006\
        );

    \I__663\ : Odrv4
    port map (
            O => \N__4006\,
            I => n4
        );

    \I__662\ : CascadeMux
    port map (
            O => \N__4003\,
            I => \n4_cascade_\
        );

    \I__661\ : CascadeMux
    port map (
            O => \N__4000\,
            I => \eeprom.i2c.n2951_cascade_\
        );

    \I__660\ : CascadeMux
    port map (
            O => \N__3997\,
            I => \eeprom.i2c.n37_cascade_\
        );

    \I__659\ : SRMux
    port map (
            O => \N__3994\,
            I => \N__3991\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3991\,
            I => \N__3987\
        );

    \I__657\ : InMux
    port map (
            O => \N__3990\,
            I => \N__3984\
        );

    \I__656\ : Odrv4
    port map (
            O => \N__3987\,
            I => \eeprom.i2c.n1935\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__3984\,
            I => \eeprom.i2c.n1935\
        );

    \I__654\ : CascadeMux
    port map (
            O => \N__3979\,
            I => \N__3975\
        );

    \I__653\ : InMux
    port map (
            O => \N__3978\,
            I => \N__3962\
        );

    \I__652\ : InMux
    port map (
            O => \N__3975\,
            I => \N__3962\
        );

    \I__651\ : InMux
    port map (
            O => \N__3974\,
            I => \N__3962\
        );

    \I__650\ : InMux
    port map (
            O => \N__3973\,
            I => \N__3962\
        );

    \I__649\ : InMux
    port map (
            O => \N__3972\,
            I => \N__3957\
        );

    \I__648\ : InMux
    port map (
            O => \N__3971\,
            I => \N__3957\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3962\,
            I => \ID_READOUT_FSM_state_0\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3957\,
            I => \ID_READOUT_FSM_state_0\
        );

    \I__645\ : CascadeMux
    port map (
            O => \N__3952\,
            I => \n20_cascade_\
        );

    \I__644\ : InMux
    port map (
            O => \N__3949\,
            I => \N__3943\
        );

    \I__643\ : InMux
    port map (
            O => \N__3948\,
            I => \N__3943\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__3943\,
            I => n6
        );

    \I__641\ : InMux
    port map (
            O => \N__3940\,
            I => \N__3937\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__3937\,
            I => n1841
        );

    \I__639\ : CascadeMux
    port map (
            O => \N__3934\,
            I => \eeprom.i2c.n9_cascade_\
        );

    \I__638\ : InMux
    port map (
            O => \N__3931\,
            I => \N__3928\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__3928\,
            I => \eeprom.i2c.n2873\
        );

    \I__636\ : InMux
    port map (
            O => \N__3925\,
            I => \N__3921\
        );

    \I__635\ : InMux
    port map (
            O => \N__3924\,
            I => \N__3918\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3921\,
            I => \eeprom.i2c.counter2_2\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3918\,
            I => \eeprom.i2c.counter2_2\
        );

    \I__632\ : InMux
    port map (
            O => \N__3913\,
            I => \N__3909\
        );

    \I__631\ : InMux
    port map (
            O => \N__3912\,
            I => \N__3906\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__3909\,
            I => \eeprom.i2c.counter2_5\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__3906\,
            I => \eeprom.i2c.counter2_5\
        );

    \I__628\ : CascadeMux
    port map (
            O => \N__3901\,
            I => \N__3898\
        );

    \I__627\ : InMux
    port map (
            O => \N__3898\,
            I => \N__3894\
        );

    \I__626\ : InMux
    port map (
            O => \N__3897\,
            I => \N__3891\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3894\,
            I => \N__3888\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3891\,
            I => \eeprom.i2c.counter2_4\
        );

    \I__623\ : Odrv4
    port map (
            O => \N__3888\,
            I => \eeprom.i2c.counter2_4\
        );

    \I__622\ : InMux
    port map (
            O => \N__3883\,
            I => \N__3879\
        );

    \I__621\ : InMux
    port map (
            O => \N__3882\,
            I => \N__3876\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__3879\,
            I => \eeprom.i2c.counter2_3\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__3876\,
            I => \eeprom.i2c.counter2_3\
        );

    \I__618\ : InMux
    port map (
            O => \N__3871\,
            I => \N__3867\
        );

    \I__617\ : InMux
    port map (
            O => \N__3870\,
            I => \N__3864\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__3867\,
            I => \eeprom.i2c.counter2_1\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3864\,
            I => \eeprom.i2c.counter2_1\
        );

    \I__614\ : CascadeMux
    port map (
            O => \N__3859\,
            I => \eeprom.i2c.n10_adj_379_cascade_\
        );

    \I__613\ : InMux
    port map (
            O => \N__3856\,
            I => \N__3852\
        );

    \I__612\ : InMux
    port map (
            O => \N__3855\,
            I => \N__3849\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__3852\,
            I => \eeprom.i2c.counter2_0\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__3849\,
            I => \eeprom.i2c.counter2_0\
        );

    \I__609\ : CascadeMux
    port map (
            O => \N__3844\,
            I => \N__3841\
        );

    \I__608\ : InMux
    port map (
            O => \N__3841\,
            I => \N__3838\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__3838\,
            I => \eeprom.i2c.n1171\
        );

    \I__606\ : InMux
    port map (
            O => \N__3835\,
            I => \N__3832\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3832\,
            I => \N__3825\
        );

    \I__604\ : InMux
    port map (
            O => \N__3831\,
            I => \N__3820\
        );

    \I__603\ : InMux
    port map (
            O => \N__3830\,
            I => \N__3820\
        );

    \I__602\ : InMux
    port map (
            O => \N__3829\,
            I => \N__3817\
        );

    \I__601\ : InMux
    port map (
            O => \N__3828\,
            I => \N__3814\
        );

    \I__600\ : Odrv4
    port map (
            O => \N__3825\,
            I => read
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3820\,
            I => read
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3817\,
            I => read
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3814\,
            I => read
        );

    \I__596\ : InMux
    port map (
            O => \N__3805\,
            I => \N__3802\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3802\,
            I => \N__3797\
        );

    \I__594\ : InMux
    port map (
            O => \N__3801\,
            I => \N__3794\
        );

    \I__593\ : InMux
    port map (
            O => \N__3800\,
            I => \N__3791\
        );

    \I__592\ : Odrv4
    port map (
            O => \N__3797\,
            I => \eeprom.n1703\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__3794\,
            I => \eeprom.n1703\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3791\,
            I => \eeprom.n1703\
        );

    \I__589\ : CascadeMux
    port map (
            O => \N__3784\,
            I => \n805_cascade_\
        );

    \I__588\ : SRMux
    port map (
            O => \N__3781\,
            I => \N__3778\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__3778\,
            I => \N__3768\
        );

    \I__586\ : InMux
    port map (
            O => \N__3777\,
            I => \N__3763\
        );

    \I__585\ : InMux
    port map (
            O => \N__3776\,
            I => \N__3763\
        );

    \I__584\ : InMux
    port map (
            O => \N__3775\,
            I => \N__3760\
        );

    \I__583\ : InMux
    port map (
            O => \N__3774\,
            I => \N__3753\
        );

    \I__582\ : InMux
    port map (
            O => \N__3773\,
            I => \N__3753\
        );

    \I__581\ : InMux
    port map (
            O => \N__3772\,
            I => \N__3753\
        );

    \I__580\ : InMux
    port map (
            O => \N__3771\,
            I => \N__3750\
        );

    \I__579\ : Odrv4
    port map (
            O => \N__3768\,
            I => state_1
        );

    \I__578\ : LocalMux
    port map (
            O => \N__3763\,
            I => state_1
        );

    \I__577\ : LocalMux
    port map (
            O => \N__3760\,
            I => state_1
        );

    \I__576\ : LocalMux
    port map (
            O => \N__3753\,
            I => state_1
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3750\,
            I => state_1
        );

    \I__574\ : CascadeMux
    port map (
            O => \N__3739\,
            I => \N__3732\
        );

    \I__573\ : CascadeMux
    port map (
            O => \N__3738\,
            I => \N__3728\
        );

    \I__572\ : CascadeMux
    port map (
            O => \N__3737\,
            I => \N__3725\
        );

    \I__571\ : CascadeMux
    port map (
            O => \N__3736\,
            I => \N__3721\
        );

    \I__570\ : InMux
    port map (
            O => \N__3735\,
            I => \N__3715\
        );

    \I__569\ : InMux
    port map (
            O => \N__3732\,
            I => \N__3712\
        );

    \I__568\ : InMux
    port map (
            O => \N__3731\,
            I => \N__3707\
        );

    \I__567\ : InMux
    port map (
            O => \N__3728\,
            I => \N__3707\
        );

    \I__566\ : InMux
    port map (
            O => \N__3725\,
            I => \N__3702\
        );

    \I__565\ : InMux
    port map (
            O => \N__3724\,
            I => \N__3702\
        );

    \I__564\ : InMux
    port map (
            O => \N__3721\,
            I => \N__3697\
        );

    \I__563\ : InMux
    port map (
            O => \N__3720\,
            I => \N__3697\
        );

    \I__562\ : InMux
    port map (
            O => \N__3719\,
            I => \N__3694\
        );

    \I__561\ : InMux
    port map (
            O => \N__3718\,
            I => \N__3691\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3715\,
            I => state_0
        );

    \I__559\ : LocalMux
    port map (
            O => \N__3712\,
            I => state_0
        );

    \I__558\ : LocalMux
    port map (
            O => \N__3707\,
            I => state_0
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3702\,
            I => state_0
        );

    \I__556\ : LocalMux
    port map (
            O => \N__3697\,
            I => state_0
        );

    \I__555\ : LocalMux
    port map (
            O => \N__3694\,
            I => state_0
        );

    \I__554\ : LocalMux
    port map (
            O => \N__3691\,
            I => state_0
        );

    \I__553\ : InMux
    port map (
            O => \N__3676\,
            I => \N__3670\
        );

    \I__552\ : InMux
    port map (
            O => \N__3675\,
            I => \N__3670\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3670\,
            I => data_ready
        );

    \I__550\ : InMux
    port map (
            O => \N__3667\,
            I => \N__3664\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3664\,
            I => n2476
        );

    \I__548\ : CascadeMux
    port map (
            O => \N__3661\,
            I => \n2476_cascade_\
        );

    \I__547\ : InMux
    port map (
            O => \N__3658\,
            I => \N__3651\
        );

    \I__546\ : InMux
    port map (
            O => \N__3657\,
            I => \N__3651\
        );

    \I__545\ : InMux
    port map (
            O => \N__3656\,
            I => \N__3648\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3651\,
            I => \N__3645\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__3648\,
            I => \N__3642\
        );

    \I__542\ : Odrv4
    port map (
            O => \N__3645\,
            I => n15
        );

    \I__541\ : Odrv4
    port map (
            O => \N__3642\,
            I => n15
        );

    \I__540\ : CascadeMux
    port map (
            O => \N__3637\,
            I => \N__3633\
        );

    \I__539\ : InMux
    port map (
            O => \N__3636\,
            I => \N__3622\
        );

    \I__538\ : InMux
    port map (
            O => \N__3633\,
            I => \N__3622\
        );

    \I__537\ : InMux
    port map (
            O => \N__3632\,
            I => \N__3622\
        );

    \I__536\ : InMux
    port map (
            O => \N__3631\,
            I => \N__3615\
        );

    \I__535\ : InMux
    port map (
            O => \N__3630\,
            I => \N__3615\
        );

    \I__534\ : InMux
    port map (
            O => \N__3629\,
            I => \N__3615\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3622\,
            I => \ID_READOUT_FSM_state_1\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3615\,
            I => \ID_READOUT_FSM_state_1\
        );

    \I__531\ : InMux
    port map (
            O => \N__3610\,
            I => \N__3607\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3607\,
            I => n20
        );

    \I__529\ : CascadeMux
    port map (
            O => \N__3604\,
            I => \N__3600\
        );

    \I__528\ : InMux
    port map (
            O => \N__3603\,
            I => \N__3595\
        );

    \I__527\ : InMux
    port map (
            O => \N__3600\,
            I => \N__3595\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3595\,
            I => data_2
        );

    \I__525\ : CascadeMux
    port map (
            O => \N__3592\,
            I => \N__3588\
        );

    \I__524\ : InMux
    port map (
            O => \N__3591\,
            I => \N__3585\
        );

    \I__523\ : InMux
    port map (
            O => \N__3588\,
            I => \N__3582\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__3585\,
            I => data_1
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3582\,
            I => data_1
        );

    \I__520\ : InMux
    port map (
            O => \N__3577\,
            I => \N__3571\
        );

    \I__519\ : InMux
    port map (
            O => \N__3576\,
            I => \N__3571\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__3571\,
            I => data_3
        );

    \I__517\ : InMux
    port map (
            O => \N__3568\,
            I => \N__3565\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3565\,
            I => \N__3561\
        );

    \I__515\ : InMux
    port map (
            O => \N__3564\,
            I => \N__3558\
        );

    \I__514\ : Odrv4
    port map (
            O => \N__3561\,
            I => data_0
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3558\,
            I => data_0
        );

    \I__512\ : CascadeMux
    port map (
            O => \N__3553\,
            I => \n10_cascade_\
        );

    \I__511\ : CascadeMux
    port map (
            O => \N__3550\,
            I => \N__3547\
        );

    \I__510\ : InMux
    port map (
            O => \N__3547\,
            I => \N__3544\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3544\,
            I => \eeprom.n4\
        );

    \I__508\ : InMux
    port map (
            O => \N__3541\,
            I => \N__3538\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3538\,
            I => \eeprom.n22\
        );

    \I__506\ : InMux
    port map (
            O => \N__3535\,
            I => \N__3532\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3532\,
            I => \eeprom.n26\
        );

    \I__504\ : InMux
    port map (
            O => \N__3529\,
            I => \N__3523\
        );

    \I__503\ : InMux
    port map (
            O => \N__3528\,
            I => \N__3523\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__3523\,
            I => \eeprom.n2727\
        );

    \I__501\ : CascadeMux
    port map (
            O => \N__3520\,
            I => \eeprom.n2727_cascade_\
        );

    \I__500\ : InMux
    port map (
            O => \N__3517\,
            I => \N__3514\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__3514\,
            I => \eeprom.i2c.n2881\
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__3511\,
            I => \eeprom.i2c.n10_adj_384_cascade_\
        );

    \I__497\ : InMux
    port map (
            O => \N__3508\,
            I => \N__3505\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__3505\,
            I => \eeprom.i2c.n10_adj_377\
        );

    \I__495\ : InMux
    port map (
            O => \N__3502\,
            I => \N__3499\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__3499\,
            I => \eeprom.i2c.n2972\
        );

    \I__493\ : CascadeMux
    port map (
            O => \N__3496\,
            I => \N__3493\
        );

    \I__492\ : InMux
    port map (
            O => \N__3493\,
            I => \N__3489\
        );

    \I__491\ : InMux
    port map (
            O => \N__3492\,
            I => \N__3486\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3489\,
            I => \eeprom.delay_counter_12\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__3486\,
            I => \eeprom.delay_counter_12\
        );

    \I__488\ : CascadeMux
    port map (
            O => \N__3481\,
            I => \N__3478\
        );

    \I__487\ : InMux
    port map (
            O => \N__3478\,
            I => \N__3474\
        );

    \I__486\ : InMux
    port map (
            O => \N__3477\,
            I => \N__3471\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3474\,
            I => \eeprom.delay_counter_10\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3471\,
            I => \eeprom.delay_counter_10\
        );

    \I__483\ : CascadeMux
    port map (
            O => \N__3466\,
            I => \N__3462\
        );

    \I__482\ : CascadeMux
    port map (
            O => \N__3465\,
            I => \N__3459\
        );

    \I__481\ : InMux
    port map (
            O => \N__3462\,
            I => \N__3456\
        );

    \I__480\ : InMux
    port map (
            O => \N__3459\,
            I => \N__3453\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__3456\,
            I => \eeprom.delay_counter_8\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__3453\,
            I => \eeprom.delay_counter_8\
        );

    \I__477\ : CascadeMux
    port map (
            O => \N__3448\,
            I => \N__3445\
        );

    \I__476\ : InMux
    port map (
            O => \N__3445\,
            I => \N__3441\
        );

    \I__475\ : InMux
    port map (
            O => \N__3444\,
            I => \N__3438\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__3441\,
            I => \eeprom.delay_counter_6\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__3438\,
            I => \eeprom.delay_counter_6\
        );

    \I__472\ : InMux
    port map (
            O => \N__3433\,
            I => \N__3430\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__3430\,
            I => \eeprom.n26_adj_388\
        );

    \I__470\ : InMux
    port map (
            O => \N__3427\,
            I => \N__3424\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3424\,
            I => \eeprom.n27\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__3421\,
            I => \eeprom.n28_cascade_\
        );

    \I__467\ : InMux
    port map (
            O => \N__3418\,
            I => \N__3415\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__3415\,
            I => \eeprom.n25\
        );

    \I__465\ : CascadeMux
    port map (
            O => \N__3412\,
            I => \eeprom.n1703_cascade_\
        );

    \I__464\ : CascadeMux
    port map (
            O => \N__3409\,
            I => \N__3398\
        );

    \I__463\ : CascadeMux
    port map (
            O => \N__3408\,
            I => \N__3394\
        );

    \I__462\ : CascadeMux
    port map (
            O => \N__3407\,
            I => \N__3390\
        );

    \I__461\ : CascadeMux
    port map (
            O => \N__3406\,
            I => \N__3386\
        );

    \I__460\ : CascadeMux
    port map (
            O => \N__3405\,
            I => \N__3382\
        );

    \I__459\ : CascadeMux
    port map (
            O => \N__3404\,
            I => \N__3378\
        );

    \I__458\ : CascadeMux
    port map (
            O => \N__3403\,
            I => \N__3374\
        );

    \I__457\ : InMux
    port map (
            O => \N__3402\,
            I => \N__3356\
        );

    \I__456\ : InMux
    port map (
            O => \N__3401\,
            I => \N__3356\
        );

    \I__455\ : InMux
    port map (
            O => \N__3398\,
            I => \N__3356\
        );

    \I__454\ : InMux
    port map (
            O => \N__3397\,
            I => \N__3356\
        );

    \I__453\ : InMux
    port map (
            O => \N__3394\,
            I => \N__3356\
        );

    \I__452\ : InMux
    port map (
            O => \N__3393\,
            I => \N__3356\
        );

    \I__451\ : InMux
    port map (
            O => \N__3390\,
            I => \N__3356\
        );

    \I__450\ : InMux
    port map (
            O => \N__3389\,
            I => \N__3356\
        );

    \I__449\ : InMux
    port map (
            O => \N__3386\,
            I => \N__3339\
        );

    \I__448\ : InMux
    port map (
            O => \N__3385\,
            I => \N__3339\
        );

    \I__447\ : InMux
    port map (
            O => \N__3382\,
            I => \N__3339\
        );

    \I__446\ : InMux
    port map (
            O => \N__3381\,
            I => \N__3339\
        );

    \I__445\ : InMux
    port map (
            O => \N__3378\,
            I => \N__3339\
        );

    \I__444\ : InMux
    port map (
            O => \N__3377\,
            I => \N__3339\
        );

    \I__443\ : InMux
    port map (
            O => \N__3374\,
            I => \N__3339\
        );

    \I__442\ : InMux
    port map (
            O => \N__3373\,
            I => \N__3339\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__3356\,
            I => \eeprom.n730\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__3339\,
            I => \eeprom.n730\
        );

    \I__439\ : InMux
    port map (
            O => \N__3334\,
            I => \bfn_21_8_0_\
        );

    \I__438\ : InMux
    port map (
            O => \N__3331\,
            I => \eeprom.i2c.n2686\
        );

    \I__437\ : InMux
    port map (
            O => \N__3328\,
            I => \eeprom.i2c.n2687\
        );

    \I__436\ : InMux
    port map (
            O => \N__3325\,
            I => \eeprom.i2c.n2688\
        );

    \I__435\ : InMux
    port map (
            O => \N__3322\,
            I => \eeprom.i2c.n2689\
        );

    \I__434\ : InMux
    port map (
            O => \N__3319\,
            I => \eeprom.i2c.n2690\
        );

    \I__433\ : InMux
    port map (
            O => \N__3316\,
            I => \N__3309\
        );

    \I__432\ : InMux
    port map (
            O => \N__3315\,
            I => \N__3309\
        );

    \I__431\ : InMux
    port map (
            O => \N__3314\,
            I => \N__3306\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__3309\,
            I => blink_counter_24
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3306\,
            I => blink_counter_24
        );

    \I__428\ : InMux
    port map (
            O => \N__3301\,
            I => \bfn_19_20_0_\
        );

    \I__427\ : InMux
    port map (
            O => \N__3298\,
            I => n2715
        );

    \I__426\ : InMux
    port map (
            O => \N__3295\,
            I => \N__3291\
        );

    \I__425\ : InMux
    port map (
            O => \N__3294\,
            I => \N__3288\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__3291\,
            I => blink_counter_25
        );

    \I__423\ : LocalMux
    port map (
            O => \N__3288\,
            I => blink_counter_25
        );

    \I__422\ : InMux
    port map (
            O => \N__3283\,
            I => \N__3279\
        );

    \I__421\ : InMux
    port map (
            O => \N__3282\,
            I => \N__3276\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__3279\,
            I => \eeprom.delay_counter_7\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__3276\,
            I => \eeprom.delay_counter_7\
        );

    \I__418\ : CascadeMux
    port map (
            O => \N__3271\,
            I => \N__3268\
        );

    \I__417\ : InMux
    port map (
            O => \N__3268\,
            I => \N__3264\
        );

    \I__416\ : InMux
    port map (
            O => \N__3267\,
            I => \N__3261\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__3264\,
            I => \eeprom.delay_counter_2\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__3261\,
            I => \eeprom.delay_counter_2\
        );

    \I__413\ : CascadeMux
    port map (
            O => \N__3256\,
            I => \N__3252\
        );

    \I__412\ : InMux
    port map (
            O => \N__3255\,
            I => \N__3249\
        );

    \I__411\ : InMux
    port map (
            O => \N__3252\,
            I => \N__3246\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__3249\,
            I => \eeprom.delay_counter_5\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3246\,
            I => \eeprom.delay_counter_5\
        );

    \I__408\ : InMux
    port map (
            O => \N__3241\,
            I => \N__3237\
        );

    \I__407\ : InMux
    port map (
            O => \N__3240\,
            I => \N__3234\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__3237\,
            I => \eeprom.delay_counter_11\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__3234\,
            I => \eeprom.delay_counter_11\
        );

    \I__404\ : SRMux
    port map (
            O => \N__3229\,
            I => \N__3226\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__3226\,
            I => \N__3223\
        );

    \I__402\ : Span4Mux_v
    port map (
            O => \N__3223\,
            I => \N__3219\
        );

    \I__401\ : SRMux
    port map (
            O => \N__3222\,
            I => \N__3216\
        );

    \I__400\ : Span4Mux_h
    port map (
            O => \N__3219\,
            I => \N__3213\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__3216\,
            I => \N__3210\
        );

    \I__398\ : Odrv4
    port map (
            O => \N__3213\,
            I => \eeprom.n1934\
        );

    \I__397\ : Odrv12
    port map (
            O => \N__3210\,
            I => \eeprom.n1934\
        );

    \I__396\ : InMux
    port map (
            O => \N__3205\,
            I => \N__3201\
        );

    \I__395\ : InMux
    port map (
            O => \N__3204\,
            I => \N__3198\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3201\,
            I => \eeprom.delay_counter_13\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__3198\,
            I => \eeprom.delay_counter_13\
        );

    \I__392\ : InMux
    port map (
            O => \N__3193\,
            I => \N__3189\
        );

    \I__391\ : InMux
    port map (
            O => \N__3192\,
            I => \N__3186\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3189\,
            I => \eeprom.delay_counter_9\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__3186\,
            I => \eeprom.delay_counter_9\
        );

    \I__388\ : CascadeMux
    port map (
            O => \N__3181\,
            I => \N__3177\
        );

    \I__387\ : CascadeMux
    port map (
            O => \N__3180\,
            I => \N__3174\
        );

    \I__386\ : InMux
    port map (
            O => \N__3177\,
            I => \N__3171\
        );

    \I__385\ : InMux
    port map (
            O => \N__3174\,
            I => \N__3168\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__3171\,
            I => \eeprom.delay_counter_0\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__3168\,
            I => \eeprom.delay_counter_0\
        );

    \I__382\ : CascadeMux
    port map (
            O => \N__3163\,
            I => \N__3160\
        );

    \I__381\ : InMux
    port map (
            O => \N__3160\,
            I => \N__3156\
        );

    \I__380\ : InMux
    port map (
            O => \N__3159\,
            I => \N__3153\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__3156\,
            I => \eeprom.delay_counter_4\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__3153\,
            I => \eeprom.delay_counter_4\
        );

    \I__377\ : CascadeMux
    port map (
            O => \N__3148\,
            I => \N__3145\
        );

    \I__376\ : InMux
    port map (
            O => \N__3145\,
            I => \N__3141\
        );

    \I__375\ : InMux
    port map (
            O => \N__3144\,
            I => \N__3138\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__3141\,
            I => \eeprom.delay_counter_14\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__3138\,
            I => \eeprom.delay_counter_14\
        );

    \I__372\ : InMux
    port map (
            O => \N__3133\,
            I => \N__3129\
        );

    \I__371\ : InMux
    port map (
            O => \N__3132\,
            I => \N__3126\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__3129\,
            I => \eeprom.delay_counter_3\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__3126\,
            I => \eeprom.delay_counter_3\
        );

    \I__368\ : CascadeMux
    port map (
            O => \N__3121\,
            I => \N__3117\
        );

    \I__367\ : InMux
    port map (
            O => \N__3120\,
            I => \N__3114\
        );

    \I__366\ : InMux
    port map (
            O => \N__3117\,
            I => \N__3111\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__3114\,
            I => \eeprom.delay_counter_1\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__3111\,
            I => \eeprom.delay_counter_1\
        );

    \I__363\ : InMux
    port map (
            O => \N__3106\,
            I => \N__3102\
        );

    \I__362\ : InMux
    port map (
            O => \N__3105\,
            I => \N__3099\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__3102\,
            I => \eeprom.delay_counter_15\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__3099\,
            I => \eeprom.delay_counter_15\
        );

    \I__359\ : CEMux
    port map (
            O => \N__3094\,
            I => \N__3090\
        );

    \I__358\ : CEMux
    port map (
            O => \N__3093\,
            I => \N__3087\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__3090\,
            I => \N__3084\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__3087\,
            I => \N__3081\
        );

    \I__355\ : Span4Mux_h
    port map (
            O => \N__3084\,
            I => \N__3077\
        );

    \I__354\ : Span4Mux_h
    port map (
            O => \N__3081\,
            I => \N__3074\
        );

    \I__353\ : InMux
    port map (
            O => \N__3080\,
            I => \N__3071\
        );

    \I__352\ : Odrv4
    port map (
            O => \N__3077\,
            I => \eeprom.n1799\
        );

    \I__351\ : Odrv4
    port map (
            O => \N__3074\,
            I => \eeprom.n1799\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__3071\,
            I => \eeprom.n1799\
        );

    \I__349\ : InMux
    port map (
            O => \N__3064\,
            I => \N__3061\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__3061\,
            I => n10_adj_398
        );

    \I__347\ : InMux
    port map (
            O => \N__3058\,
            I => \bfn_19_19_0_\
        );

    \I__346\ : InMux
    port map (
            O => \N__3055\,
            I => \N__3052\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__3052\,
            I => n9
        );

    \I__344\ : InMux
    port map (
            O => \N__3049\,
            I => n2707
        );

    \I__343\ : InMux
    port map (
            O => \N__3046\,
            I => \N__3043\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__3043\,
            I => n8_adj_397
        );

    \I__341\ : InMux
    port map (
            O => \N__3040\,
            I => n2708
        );

    \I__340\ : InMux
    port map (
            O => \N__3037\,
            I => \N__3034\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__3034\,
            I => n7
        );

    \I__338\ : InMux
    port map (
            O => \N__3031\,
            I => n2709
        );

    \I__337\ : InMux
    port map (
            O => \N__3028\,
            I => \N__3025\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__3025\,
            I => n6_adj_396
        );

    \I__335\ : InMux
    port map (
            O => \N__3022\,
            I => n2710
        );

    \I__334\ : InMux
    port map (
            O => \N__3019\,
            I => \N__3012\
        );

    \I__333\ : InMux
    port map (
            O => \N__3018\,
            I => \N__3012\
        );

    \I__332\ : InMux
    port map (
            O => \N__3017\,
            I => \N__3009\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__3012\,
            I => blink_counter_21
        );

    \I__330\ : LocalMux
    port map (
            O => \N__3009\,
            I => blink_counter_21
        );

    \I__329\ : InMux
    port map (
            O => \N__3004\,
            I => n2711
        );

    \I__328\ : InMux
    port map (
            O => \N__3001\,
            I => \N__2994\
        );

    \I__327\ : InMux
    port map (
            O => \N__3000\,
            I => \N__2994\
        );

    \I__326\ : InMux
    port map (
            O => \N__2999\,
            I => \N__2991\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__2994\,
            I => blink_counter_22
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2991\,
            I => blink_counter_22
        );

    \I__323\ : InMux
    port map (
            O => \N__2986\,
            I => n2712
        );

    \I__322\ : CascadeMux
    port map (
            O => \N__2983\,
            I => \N__2979\
        );

    \I__321\ : CascadeMux
    port map (
            O => \N__2982\,
            I => \N__2976\
        );

    \I__320\ : InMux
    port map (
            O => \N__2979\,
            I => \N__2970\
        );

    \I__319\ : InMux
    port map (
            O => \N__2976\,
            I => \N__2970\
        );

    \I__318\ : InMux
    port map (
            O => \N__2975\,
            I => \N__2967\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__2970\,
            I => blink_counter_23
        );

    \I__316\ : LocalMux
    port map (
            O => \N__2967\,
            I => blink_counter_23
        );

    \I__315\ : InMux
    port map (
            O => \N__2962\,
            I => n2713
        );

    \I__314\ : InMux
    port map (
            O => \N__2959\,
            I => \N__2956\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__2956\,
            I => n19
        );

    \I__312\ : InMux
    port map (
            O => \N__2953\,
            I => n2697
        );

    \I__311\ : InMux
    port map (
            O => \N__2950\,
            I => \N__2947\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__2947\,
            I => n18_adj_402
        );

    \I__309\ : InMux
    port map (
            O => \N__2944\,
            I => \bfn_19_18_0_\
        );

    \I__308\ : InMux
    port map (
            O => \N__2941\,
            I => \N__2938\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2938\,
            I => n17
        );

    \I__306\ : InMux
    port map (
            O => \N__2935\,
            I => n2699
        );

    \I__305\ : InMux
    port map (
            O => \N__2932\,
            I => \N__2929\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__2929\,
            I => n16
        );

    \I__303\ : InMux
    port map (
            O => \N__2926\,
            I => n2700
        );

    \I__302\ : InMux
    port map (
            O => \N__2923\,
            I => \N__2920\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2920\,
            I => n15_adj_401
        );

    \I__300\ : InMux
    port map (
            O => \N__2917\,
            I => n2701
        );

    \I__299\ : InMux
    port map (
            O => \N__2914\,
            I => \N__2911\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2911\,
            I => n14_adj_400
        );

    \I__297\ : InMux
    port map (
            O => \N__2908\,
            I => n2702
        );

    \I__296\ : InMux
    port map (
            O => \N__2905\,
            I => \N__2902\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2902\,
            I => n13_adj_399
        );

    \I__294\ : InMux
    port map (
            O => \N__2899\,
            I => n2703
        );

    \I__293\ : InMux
    port map (
            O => \N__2896\,
            I => \N__2893\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2893\,
            I => n12
        );

    \I__291\ : InMux
    port map (
            O => \N__2890\,
            I => n2704
        );

    \I__290\ : InMux
    port map (
            O => \N__2887\,
            I => \N__2884\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2884\,
            I => n11
        );

    \I__288\ : InMux
    port map (
            O => \N__2881\,
            I => n2705
        );

    \I__287\ : InMux
    port map (
            O => \N__2878\,
            I => \eeprom.n2685\
        );

    \I__286\ : InMux
    port map (
            O => \N__2875\,
            I => \N__2872\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__2872\,
            I => n26
        );

    \I__284\ : InMux
    port map (
            O => \N__2869\,
            I => \bfn_19_17_0_\
        );

    \I__283\ : InMux
    port map (
            O => \N__2866\,
            I => \N__2863\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__2863\,
            I => n25_adj_407
        );

    \I__281\ : InMux
    port map (
            O => \N__2860\,
            I => n2691
        );

    \I__280\ : InMux
    port map (
            O => \N__2857\,
            I => \N__2854\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2854\,
            I => n24_adj_406
        );

    \I__278\ : InMux
    port map (
            O => \N__2851\,
            I => n2692
        );

    \I__277\ : InMux
    port map (
            O => \N__2848\,
            I => \N__2845\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__2845\,
            I => n23_adj_405
        );

    \I__275\ : InMux
    port map (
            O => \N__2842\,
            I => n2693
        );

    \I__274\ : InMux
    port map (
            O => \N__2839\,
            I => \N__2836\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__2836\,
            I => n22_adj_404
        );

    \I__272\ : InMux
    port map (
            O => \N__2833\,
            I => n2694
        );

    \I__271\ : InMux
    port map (
            O => \N__2830\,
            I => \N__2827\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2827\,
            I => n21
        );

    \I__269\ : InMux
    port map (
            O => \N__2824\,
            I => n2695
        );

    \I__268\ : InMux
    port map (
            O => \N__2821\,
            I => \N__2818\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__2818\,
            I => n20_adj_403
        );

    \I__266\ : InMux
    port map (
            O => \N__2815\,
            I => n2696
        );

    \I__265\ : InMux
    port map (
            O => \N__2812\,
            I => \eeprom.n2676\
        );

    \I__264\ : InMux
    port map (
            O => \N__2809\,
            I => \eeprom.n2677\
        );

    \I__263\ : InMux
    port map (
            O => \N__2806\,
            I => \bfn_19_14_0_\
        );

    \I__262\ : InMux
    port map (
            O => \N__2803\,
            I => \eeprom.n2679\
        );

    \I__261\ : InMux
    port map (
            O => \N__2800\,
            I => \eeprom.n2680\
        );

    \I__260\ : InMux
    port map (
            O => \N__2797\,
            I => \eeprom.n2681\
        );

    \I__259\ : InMux
    port map (
            O => \N__2794\,
            I => \eeprom.n2682\
        );

    \I__258\ : InMux
    port map (
            O => \N__2791\,
            I => \eeprom.n2683\
        );

    \I__257\ : InMux
    port map (
            O => \N__2788\,
            I => \eeprom.n2684\
        );

    \I__256\ : CascadeMux
    port map (
            O => \N__2785\,
            I => \n2955_cascade_\
        );

    \I__255\ : IoInMux
    port map (
            O => \N__2782\,
            I => \N__2779\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__2779\,
            I => \N__2776\
        );

    \I__253\ : Span4Mux_s1_v
    port map (
            O => \N__2776\,
            I => \N__2773\
        );

    \I__252\ : Sp12to4
    port map (
            O => \N__2773\,
            I => \N__2770\
        );

    \I__251\ : Span12Mux_h
    port map (
            O => \N__2770\,
            I => \N__2767\
        );

    \I__250\ : Span12Mux_v
    port map (
            O => \N__2767\,
            I => \N__2764\
        );

    \I__249\ : Odrv12
    port map (
            O => \N__2764\,
            I => \LED_c\
        );

    \I__248\ : InMux
    port map (
            O => \N__2761\,
            I => \N__2758\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__2758\,
            I => n2954
        );

    \I__246\ : InMux
    port map (
            O => \N__2755\,
            I => \eeprom.n2671\
        );

    \I__245\ : InMux
    port map (
            O => \N__2752\,
            I => \eeprom.n2672\
        );

    \I__244\ : InMux
    port map (
            O => \N__2749\,
            I => \eeprom.n2673\
        );

    \I__243\ : InMux
    port map (
            O => \N__2746\,
            I => \eeprom.n2674\
        );

    \I__242\ : InMux
    port map (
            O => \N__2743\,
            I => \eeprom.n2675\
        );

    \I__241\ : IoInMux
    port map (
            O => \N__2740\,
            I => \N__2737\
        );

    \I__240\ : LocalMux
    port map (
            O => \N__2737\,
            I => \N__2734\
        );

    \I__239\ : IoSpan4Mux
    port map (
            O => \N__2734\,
            I => \N__2731\
        );

    \I__238\ : IoSpan4Mux
    port map (
            O => \N__2731\,
            I => \N__2728\
        );

    \I__237\ : IoSpan4Mux
    port map (
            O => \N__2728\,
            I => \N__2725\
        );

    \I__236\ : Odrv4
    port map (
            O => \N__2725\,
            I => \CLK_pad_gb_input\
        );

    \INVeeprom.i2c.i2c_scl_enable_123C\ : INV
    port map (
            O => \INVeeprom.i2c.i2c_scl_enable_123C_net\,
            I => \N__5775\
        );

    \INVeeprom.i2c.sda_out_131C\ : INV
    port map (
            O => \INVeeprom.i2c.sda_out_131C_net\,
            I => \N__5756\
        );

    \INVeeprom.i2c.write_enable_130C\ : INV
    port map (
            O => \INVeeprom.i2c.write_enable_130C_net\,
            I => \N__5767\
        );

    \INVeeprom.i2c.data_out_i0_i4C\ : INV
    port map (
            O => \INVeeprom.i2c.data_out_i0_i4C_net\,
            I => \N__5741\
        );

    \INVeeprom.i2c.data_out_i0_i3C\ : INV
    port map (
            O => \INVeeprom.i2c.data_out_i0_i3C_net\,
            I => \N__5766\
        );

    \INVeeprom.i2c.data_out_i0_i1C\ : INV
    port map (
            O => \INVeeprom.i2c.data_out_i0_i1C_net\,
            I => \N__5749\
        );

    \IN_MUX_bfv_22_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_11_0_\
        );

    \IN_MUX_bfv_21_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_8_0_\
        );

    \IN_MUX_bfv_19_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_13_0_\
        );

    \IN_MUX_bfv_19_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n2678\,
            carryinitout => \bfn_19_14_0_\
        );

    \IN_MUX_bfv_19_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_17_0_\
        );

    \IN_MUX_bfv_19_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2698,
            carryinitout => \bfn_19_18_0_\
        );

    \IN_MUX_bfv_19_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2706,
            carryinitout => \bfn_19_19_0_\
        );

    \IN_MUX_bfv_19_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2714,
            carryinitout => \bfn_19_20_0_\
        );

    \IN_MUX_bfv_23_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_23_13_0_\
        );

    \IN_MUX_bfv_23_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2640,
            carryinitout => \bfn_23_14_0_\
        );

    \IN_MUX_bfv_23_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2648,
            carryinitout => \bfn_23_15_0_\
        );

    \IN_MUX_bfv_23_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n2656,
            carryinitout => \bfn_23_16_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2740\,
            GLOBALBUFFEROUTPUT => \CLK_c\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \i1941_4_lut_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010110000"
        )
    port map (
            in0 => \N__3316\,
            in1 => \N__3001\,
            in2 => \N__2983\,
            in3 => \N__3019\,
            lcout => OPEN,
            ltout => \n2955_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1942_3_lut_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__2761\,
            in1 => \_gnd_net_\,
            in2 => \N__2785\,
            in3 => \N__3295\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1940_4_lut_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000000"
        )
    port map (
            in0 => \N__3315\,
            in1 => \N__3000\,
            in2 => \N__2982\,
            in3 => \N__3018\,
            lcout => n2954,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.delay_counter_i0_i0_LC_19_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3373\,
            in2 => \N__3181\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.delay_counter_0\,
            ltout => OPEN,
            carryin => \bfn_19_13_0_\,
            carryout => \eeprom.n2671\,
            clk => \N__5840\,
            ce => \N__3094\,
            sr => \N__3222\
        );

    \eeprom.delay_counter_i0_i1_LC_19_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3120\,
            in2 => \N__3403\,
            in3 => \N__2755\,
            lcout => \eeprom.delay_counter_1\,
            ltout => OPEN,
            carryin => \eeprom.n2671\,
            carryout => \eeprom.n2672\,
            clk => \N__5840\,
            ce => \N__3094\,
            sr => \N__3222\
        );

    \eeprom.delay_counter_i0_i2_LC_19_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3377\,
            in2 => \N__3271\,
            in3 => \N__2752\,
            lcout => \eeprom.delay_counter_2\,
            ltout => OPEN,
            carryin => \eeprom.n2672\,
            carryout => \eeprom.n2673\,
            clk => \N__5840\,
            ce => \N__3094\,
            sr => \N__3222\
        );

    \eeprom.delay_counter_i0_i3_LC_19_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3133\,
            in2 => \N__3404\,
            in3 => \N__2749\,
            lcout => \eeprom.delay_counter_3\,
            ltout => OPEN,
            carryin => \eeprom.n2673\,
            carryout => \eeprom.n2674\,
            clk => \N__5840\,
            ce => \N__3094\,
            sr => \N__3222\
        );

    \eeprom.delay_counter_i0_i4_LC_19_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3381\,
            in2 => \N__3163\,
            in3 => \N__2746\,
            lcout => \eeprom.delay_counter_4\,
            ltout => OPEN,
            carryin => \eeprom.n2674\,
            carryout => \eeprom.n2675\,
            clk => \N__5840\,
            ce => \N__3094\,
            sr => \N__3222\
        );

    \eeprom.delay_counter_i0_i5_LC_19_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3255\,
            in2 => \N__3405\,
            in3 => \N__2743\,
            lcout => \eeprom.delay_counter_5\,
            ltout => OPEN,
            carryin => \eeprom.n2675\,
            carryout => \eeprom.n2676\,
            clk => \N__5840\,
            ce => \N__3094\,
            sr => \N__3222\
        );

    \eeprom.delay_counter_i0_i6_LC_19_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3385\,
            in2 => \N__3448\,
            in3 => \N__2812\,
            lcout => \eeprom.delay_counter_6\,
            ltout => OPEN,
            carryin => \eeprom.n2676\,
            carryout => \eeprom.n2677\,
            clk => \N__5840\,
            ce => \N__3094\,
            sr => \N__3222\
        );

    \eeprom.delay_counter_i0_i7_LC_19_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3283\,
            in2 => \N__3406\,
            in3 => \N__2809\,
            lcout => \eeprom.delay_counter_7\,
            ltout => OPEN,
            carryin => \eeprom.n2677\,
            carryout => \eeprom.n2678\,
            clk => \N__5840\,
            ce => \N__3094\,
            sr => \N__3222\
        );

    \eeprom.delay_counter_i0_i8_LC_19_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3389\,
            in2 => \N__3466\,
            in3 => \N__2806\,
            lcout => \eeprom.delay_counter_8\,
            ltout => OPEN,
            carryin => \bfn_19_14_0_\,
            carryout => \eeprom.n2679\,
            clk => \N__5838\,
            ce => \N__3093\,
            sr => \N__3229\
        );

    \eeprom.delay_counter_i0_i9_LC_19_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3193\,
            in2 => \N__3407\,
            in3 => \N__2803\,
            lcout => \eeprom.delay_counter_9\,
            ltout => OPEN,
            carryin => \eeprom.n2679\,
            carryout => \eeprom.n2680\,
            clk => \N__5838\,
            ce => \N__3093\,
            sr => \N__3229\
        );

    \eeprom.delay_counter_i0_i10_LC_19_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3393\,
            in2 => \N__3481\,
            in3 => \N__2800\,
            lcout => \eeprom.delay_counter_10\,
            ltout => OPEN,
            carryin => \eeprom.n2680\,
            carryout => \eeprom.n2681\,
            clk => \N__5838\,
            ce => \N__3093\,
            sr => \N__3229\
        );

    \eeprom.delay_counter_i0_i11_LC_19_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3241\,
            in2 => \N__3408\,
            in3 => \N__2797\,
            lcout => \eeprom.delay_counter_11\,
            ltout => OPEN,
            carryin => \eeprom.n2681\,
            carryout => \eeprom.n2682\,
            clk => \N__5838\,
            ce => \N__3093\,
            sr => \N__3229\
        );

    \eeprom.delay_counter_i0_i12_LC_19_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3397\,
            in2 => \N__3496\,
            in3 => \N__2794\,
            lcout => \eeprom.delay_counter_12\,
            ltout => OPEN,
            carryin => \eeprom.n2682\,
            carryout => \eeprom.n2683\,
            clk => \N__5838\,
            ce => \N__3093\,
            sr => \N__3229\
        );

    \eeprom.delay_counter_i0_i13_LC_19_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3205\,
            in2 => \N__3409\,
            in3 => \N__2791\,
            lcout => \eeprom.delay_counter_13\,
            ltout => OPEN,
            carryin => \eeprom.n2683\,
            carryout => \eeprom.n2684\,
            clk => \N__5838\,
            ce => \N__3093\,
            sr => \N__3229\
        );

    \eeprom.delay_counter_i0_i14_LC_19_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3401\,
            in2 => \N__3148\,
            in3 => \N__2788\,
            lcout => \eeprom.delay_counter_14\,
            ltout => OPEN,
            carryin => \eeprom.n2684\,
            carryout => \eeprom.n2685\,
            clk => \N__5838\,
            ce => \N__3093\,
            sr => \N__3229\
        );

    \eeprom.delay_counter_i0_i15_LC_19_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__3402\,
            in1 => \N__3106\,
            in2 => \_gnd_net_\,
            in3 => \N__2878\,
            lcout => \eeprom.delay_counter_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5838\,
            ce => \N__3093\,
            sr => \N__3229\
        );

    \blink_counter_409__i0_LC_19_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2875\,
            in2 => \_gnd_net_\,
            in3 => \N__2869\,
            lcout => n26,
            ltout => OPEN,
            carryin => \bfn_19_17_0_\,
            carryout => n2691,
            clk => \N__5835\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i1_LC_19_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2866\,
            in2 => \_gnd_net_\,
            in3 => \N__2860\,
            lcout => n25_adj_407,
            ltout => OPEN,
            carryin => n2691,
            carryout => n2692,
            clk => \N__5835\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i2_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2857\,
            in2 => \_gnd_net_\,
            in3 => \N__2851\,
            lcout => n24_adj_406,
            ltout => OPEN,
            carryin => n2692,
            carryout => n2693,
            clk => \N__5835\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i3_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2848\,
            in2 => \_gnd_net_\,
            in3 => \N__2842\,
            lcout => n23_adj_405,
            ltout => OPEN,
            carryin => n2693,
            carryout => n2694,
            clk => \N__5835\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i4_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2839\,
            in2 => \_gnd_net_\,
            in3 => \N__2833\,
            lcout => n22_adj_404,
            ltout => OPEN,
            carryin => n2694,
            carryout => n2695,
            clk => \N__5835\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i5_LC_19_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2830\,
            in2 => \_gnd_net_\,
            in3 => \N__2824\,
            lcout => n21,
            ltout => OPEN,
            carryin => n2695,
            carryout => n2696,
            clk => \N__5835\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i6_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2821\,
            in2 => \_gnd_net_\,
            in3 => \N__2815\,
            lcout => n20_adj_403,
            ltout => OPEN,
            carryin => n2696,
            carryout => n2697,
            clk => \N__5835\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i7_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2959\,
            in2 => \_gnd_net_\,
            in3 => \N__2953\,
            lcout => n19,
            ltout => OPEN,
            carryin => n2697,
            carryout => n2698,
            clk => \N__5835\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i8_LC_19_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2950\,
            in2 => \_gnd_net_\,
            in3 => \N__2944\,
            lcout => n18_adj_402,
            ltout => OPEN,
            carryin => \bfn_19_18_0_\,
            carryout => n2699,
            clk => \N__5836\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i9_LC_19_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2941\,
            in2 => \_gnd_net_\,
            in3 => \N__2935\,
            lcout => n17,
            ltout => OPEN,
            carryin => n2699,
            carryout => n2700,
            clk => \N__5836\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i10_LC_19_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2932\,
            in2 => \_gnd_net_\,
            in3 => \N__2926\,
            lcout => n16,
            ltout => OPEN,
            carryin => n2700,
            carryout => n2701,
            clk => \N__5836\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i11_LC_19_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2923\,
            in2 => \_gnd_net_\,
            in3 => \N__2917\,
            lcout => n15_adj_401,
            ltout => OPEN,
            carryin => n2701,
            carryout => n2702,
            clk => \N__5836\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i12_LC_19_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2914\,
            in2 => \_gnd_net_\,
            in3 => \N__2908\,
            lcout => n14_adj_400,
            ltout => OPEN,
            carryin => n2702,
            carryout => n2703,
            clk => \N__5836\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i13_LC_19_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2905\,
            in2 => \_gnd_net_\,
            in3 => \N__2899\,
            lcout => n13_adj_399,
            ltout => OPEN,
            carryin => n2703,
            carryout => n2704,
            clk => \N__5836\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i14_LC_19_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2896\,
            in2 => \_gnd_net_\,
            in3 => \N__2890\,
            lcout => n12,
            ltout => OPEN,
            carryin => n2704,
            carryout => n2705,
            clk => \N__5836\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i15_LC_19_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2887\,
            in2 => \_gnd_net_\,
            in3 => \N__2881\,
            lcout => n11,
            ltout => OPEN,
            carryin => n2705,
            carryout => n2706,
            clk => \N__5836\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i16_LC_19_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3064\,
            in2 => \_gnd_net_\,
            in3 => \N__3058\,
            lcout => n10_adj_398,
            ltout => OPEN,
            carryin => \bfn_19_19_0_\,
            carryout => n2707,
            clk => \N__5837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i17_LC_19_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3055\,
            in2 => \_gnd_net_\,
            in3 => \N__3049\,
            lcout => n9,
            ltout => OPEN,
            carryin => n2707,
            carryout => n2708,
            clk => \N__5837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i18_LC_19_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3046\,
            in2 => \_gnd_net_\,
            in3 => \N__3040\,
            lcout => n8_adj_397,
            ltout => OPEN,
            carryin => n2708,
            carryout => n2709,
            clk => \N__5837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i19_LC_19_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3037\,
            in2 => \_gnd_net_\,
            in3 => \N__3031\,
            lcout => n7,
            ltout => OPEN,
            carryin => n2709,
            carryout => n2710,
            clk => \N__5837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i20_LC_19_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3028\,
            in2 => \_gnd_net_\,
            in3 => \N__3022\,
            lcout => n6_adj_396,
            ltout => OPEN,
            carryin => n2710,
            carryout => n2711,
            clk => \N__5837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i21_LC_19_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3017\,
            in2 => \_gnd_net_\,
            in3 => \N__3004\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n2711,
            carryout => n2712,
            clk => \N__5837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i22_LC_19_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2999\,
            in2 => \_gnd_net_\,
            in3 => \N__2986\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n2712,
            carryout => n2713,
            clk => \N__5837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i23_LC_19_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2975\,
            in2 => \_gnd_net_\,
            in3 => \N__2962\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n2713,
            carryout => n2714,
            clk => \N__5837\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i24_LC_19_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3314\,
            in2 => \_gnd_net_\,
            in3 => \N__3301\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_19_20_0_\,
            carryout => n2715,
            clk => \N__5839\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_409__i25_LC_19_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3294\,
            in2 => \_gnd_net_\,
            in3 => \N__3298\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5839\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.enable_39_LC_20_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__5940\,
            in1 => \N__3835\,
            in2 => \N__3739\,
            in3 => \N__3805\,
            lcout => \eeprom.enable\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5844\,
            ce => 'H',
            sr => \N__3781\
        );

    \eeprom.i10_4_lut_LC_20_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3282\,
            in1 => \N__3267\,
            in2 => \N__3256\,
            in3 => \N__3240\,
            lcout => \eeprom.n26_adj_388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1007_2_lut_LC_20_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3719\,
            in2 => \_gnd_net_\,
            in3 => \N__3080\,
            lcout => \eeprom.n1934\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i9_4_lut_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3204\,
            in1 => \N__3192\,
            in2 => \N__3180\,
            in3 => \N__3159\,
            lcout => \eeprom.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i11_4_lut_LC_20_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3144\,
            in1 => \N__3132\,
            in2 => \N__3121\,
            in3 => \N__3105\,
            lcout => \eeprom.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_LC_20_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__3771\,
            in1 => \N__3718\,
            in2 => \_gnd_net_\,
            in3 => \N__3828\,
            lcout => \eeprom.n1799\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i12_4_lut_LC_20_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3492\,
            in1 => \N__3477\,
            in2 => \N__3465\,
            in3 => \N__3444\,
            lcout => OPEN,
            ltout => \eeprom.n28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i15_4_lut_LC_20_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3433\,
            in1 => \N__3427\,
            in2 => \N__3421\,
            in3 => \N__3418\,
            lcout => \eeprom.n1703\,
            ltout => \eeprom.n1703_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_adj_4_LC_20_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__5941\,
            in1 => \_gnd_net_\,
            in2 => \N__3412\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n730\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.counter2_410_411__i1_LC_21_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3855\,
            in2 => \_gnd_net_\,
            in3 => \N__3334\,
            lcout => \eeprom.i2c.counter2_0\,
            ltout => OPEN,
            carryin => \bfn_21_8_0_\,
            carryout => \eeprom.i2c.n2686\,
            clk => \N__5850\,
            ce => 'H',
            sr => \N__3994\
        );

    \eeprom.i2c.counter2_410_411__i2_LC_21_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3870\,
            in2 => \_gnd_net_\,
            in3 => \N__3331\,
            lcout => \eeprom.i2c.counter2_1\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2686\,
            carryout => \eeprom.i2c.n2687\,
            clk => \N__5850\,
            ce => 'H',
            sr => \N__3994\
        );

    \eeprom.i2c.counter2_410_411__i3_LC_21_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3925\,
            in2 => \_gnd_net_\,
            in3 => \N__3328\,
            lcout => \eeprom.i2c.counter2_2\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2687\,
            carryout => \eeprom.i2c.n2688\,
            clk => \N__5850\,
            ce => 'H',
            sr => \N__3994\
        );

    \eeprom.i2c.counter2_410_411__i4_LC_21_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3883\,
            in2 => \_gnd_net_\,
            in3 => \N__3325\,
            lcout => \eeprom.i2c.counter2_3\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2688\,
            carryout => \eeprom.i2c.n2689\,
            clk => \N__5850\,
            ce => 'H',
            sr => \N__3994\
        );

    \eeprom.i2c.counter2_410_411__i5_LC_21_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3897\,
            in2 => \_gnd_net_\,
            in3 => \N__3322\,
            lcout => \eeprom.i2c.counter2_4\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2689\,
            carryout => \eeprom.i2c.n2690\,
            clk => \N__5850\,
            ce => 'H',
            sr => \N__3994\
        );

    \eeprom.i2c.counter2_410_411__i6_LC_21_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3913\,
            in2 => \_gnd_net_\,
            in3 => \N__3319\,
            lcout => \eeprom.i2c.counter2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5850\,
            ce => 'H',
            sr => \N__3994\
        );

    \eeprom.i2c.state_7__I_0_140_i10_2_lut_LC_21_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__6040\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6280\,
            lcout => \eeprom.i2c.n10_adj_377\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_43_i10_2_lut_LC_21_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6267\,
            in2 => \_gnd_net_\,
            in3 => \N__6039\,
            lcout => \eeprom.i2c.n10_adj_384\,
            ltout => \eeprom.i2c.n10_adj_384_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1964_4_lut_LC_21_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011011101"
        )
    port map (
            in0 => \N__4771\,
            in1 => \N__4631\,
            in2 => \N__3511\,
            in3 => \N__3508\,
            lcout => \eeprom.i2c.n2972\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_i0_i3_LC_21_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__4483\,
            in1 => \N__6184\,
            in2 => \N__6460\,
            in3 => \N__3502\,
            lcout => \eeprom.state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5765\,
            ce => \N__4558\,
            sr => \N__4024\
        );

    \eeprom.i2c.data_out_i0_i1_LC_21_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__4015\,
            in1 => \N__4635\,
            in2 => \N__3592\,
            in3 => \N__4162\,
            lcout => data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.data_out_i0_i1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i0_LC_21_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__3564\,
            in1 => \N__4014\,
            in2 => \N__4656\,
            in3 => \N__4222\,
            lcout => data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.data_out_i0_i1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i3_LC_21_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__3576\,
            in1 => \N__4165\,
            in2 => \N__4657\,
            in3 => \N__4297\,
            lcout => data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.data_out_i0_i3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_adj_7_LC_21_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__6190\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6072\,
            lcout => \eeprom.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i2_LC_21_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__4225\,
            in1 => \N__4665\,
            in2 => \N__3604\,
            in3 => \N__4296\,
            lcout => data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.data_out_i0_i3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_LC_21_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3603\,
            in2 => \_gnd_net_\,
            in3 => \N__3591\,
            lcout => OPEN,
            ltout => \n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_LC_21_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3577\,
            in1 => \N__3568\,
            in2 => \N__3553\,
            in3 => \N__4243\,
            lcout => n15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.state__i1_LC_21_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111010000"
        )
    port map (
            in0 => \N__3830\,
            in1 => \N__3517\,
            in2 => \N__3550\,
            in3 => \N__3541\,
            lcout => state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_3_lut_LC_21_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__3773\,
            in1 => \_gnd_net_\,
            in2 => \N__3736\,
            in3 => \N__5942\,
            lcout => \eeprom.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.state__i0_LC_21_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__3775\,
            in1 => \N__3831\,
            in2 => \N__3737\,
            in3 => \N__3529\,
            lcout => state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_2_lut_4_lut_LC_21_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__3724\,
            in1 => \N__3772\,
            in2 => \_gnd_net_\,
            in3 => \N__3528\,
            lcout => \eeprom.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i3_4_lut_LC_21_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6459\,
            in1 => \N__3535\,
            in2 => \N__6329\,
            in3 => \N__3800\,
            lcout => \eeprom.n2727\,
            ltout => \eeprom.n2727_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1867_3_lut_LC_21_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3774\,
            in2 => \N__3520\,
            in3 => \N__3720\,
            lcout => \eeprom.i2c.n2881\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2009_2_lut_3_lut_LC_21_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__3656\,
            in1 => \N__3971\,
            in2 => \_gnd_net_\,
            in3 => \N__3630\,
            lcout => n1740,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_21_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3629\,
            in2 => \_gnd_net_\,
            in3 => \N__3675\,
            lcout => n6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \read_26_LC_21_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3972\,
            in2 => \_gnd_net_\,
            in3 => \N__3631\,
            lcout => read,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5842\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1197_4_lut_LC_21_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__5946\,
            in1 => \N__3829\,
            in2 => \N__3738\,
            in3 => \N__3801\,
            lcout => OPEN,
            ltout => \n805_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rw_43_LC_21_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__3777\,
            in1 => \N__4797\,
            in2 => \N__3784\,
            in3 => \N__3731\,
            lcout => rw,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5842\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.data_ready_42_LC_21_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001100"
        )
    port map (
            in0 => \N__3676\,
            in1 => \N__3776\,
            in2 => \N__5947\,
            in3 => \N__3735\,
            lcout => data_ready,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5842\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ID_READOUT_FSM_state__i0_LC_21_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001011100"
        )
    port map (
            in0 => \N__3949\,
            in1 => \N__3667\,
            in2 => \N__3979\,
            in3 => \N__3610\,
            lcout => \ID_READOUT_FSM_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1547_2_lut_3_lut_4_lut_LC_21_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__4425\,
            in1 => \N__3657\,
            in2 => \N__3637\,
            in3 => \N__3974\,
            lcout => n2476,
            ltout => \n2476_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ID_READOUT_FSM_state__i1_LC_21_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__3978\,
            in1 => \N__3636\,
            in2 => \N__3661\,
            in3 => \N__3940\,
            lcout => \ID_READOUT_FSM_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5841\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1844_2_lut_3_lut_LC_21_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__3658\,
            in1 => \N__3632\,
            in2 => \_gnd_net_\,
            in3 => \N__4424\,
            lcout => n20,
            ltout => \n20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_3_lut_LC_21_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3973\,
            in2 => \N__3952\,
            in3 => \N__3948\,
            lcout => n1841,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i17_4_lut_LC_22_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110001010000"
        )
    port map (
            in0 => \N__3931\,
            in1 => \N__4702\,
            in2 => \N__3844\,
            in3 => \N__4360\,
            lcout => \eeprom.i2c.n1837\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1849_2_lut_4_lut_LC_22_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__4311\,
            in1 => \N__4335\,
            in2 => \N__4639\,
            in3 => \N__6429\,
            lcout => \eeprom.i2c.n1928\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i22_3_lut_3_lut_LC_22_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001100"
        )
    port map (
            in0 => \N__6171\,
            in1 => \N__6418\,
            in2 => \_gnd_net_\,
            in3 => \N__6297\,
            lcout => \eeprom.i2c.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_43_i9_2_lut_LC_22_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__6419\,
            in1 => \N__6172\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.i2c.n9\,
            ltout => \eeprom.i2c.n9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1860_2_lut_3_lut_LC_22_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4619\,
            in2 => \N__3934\,
            in3 => \N__4310\,
            lcout => \eeprom.i2c.n2873\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i4_4_lut_LC_22_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3924\,
            in1 => \N__3912\,
            in2 => \N__3901\,
            in3 => \N__3882\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n10_adj_379_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i5_3_lut_LC_22_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3871\,
            in2 => \N__3859\,
            in3 => \N__3856\,
            lcout => \eeprom.i2c.n1935\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_3_lut_LC_22_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6298\,
            in1 => \N__6428\,
            in2 => \_gnd_net_\,
            in3 => \N__6067\,
            lcout => \eeprom.i2c.n1171\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2006_3_lut_4_lut_LC_22_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__6010\,
            in1 => \N__6135\,
            in2 => \N__4543\,
            in3 => \N__6281\,
            lcout => \eeprom.i2c.n2927\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i56_3_lut_3_lut_LC_22_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001100110"
        )
    port map (
            in0 => \N__6408\,
            in1 => \N__6248\,
            in2 => \_gnd_net_\,
            in3 => \N__6008\,
            lcout => \eeprom.i2c.n33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_60_i4_2_lut_LC_22_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4844\,
            in2 => \_gnd_net_\,
            in3 => \N__4918\,
            lcout => n4,
            ltout => \n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i3_4_lut_LC_22_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4060\,
            in1 => \N__4099\,
            in2 => \N__4003\,
            in3 => \N__4080\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n2951_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i3_4_lut_adj_8_LC_22_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4041\,
            in1 => \N__4258\,
            in2 => \N__4000\,
            in3 => \N__4875\,
            lcout => \eeprom.i2c.n1054\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_4_lut_4_lut_LC_22_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110010"
        )
    port map (
            in0 => \N__6409\,
            in1 => \N__6249\,
            in2 => \N__6170\,
            in3 => \N__6009\,
            lcout => \eeprom.i2c.n37\,
            ltout => \eeprom.i2c.n37_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1856_3_lut_LC_22_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6134\,
            in2 => \N__3997\,
            in3 => \N__4347\,
            lcout => \eeprom.i2c.n2869\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2c_clk_121_LC_22_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5665\,
            in2 => \_gnd_net_\,
            in3 => \N__3990\,
            lcout => \eeprom.i2c.i2c_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5851\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_i0_i2_LC_22_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4643\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5368\,
            lcout => \eeprom.i2c.state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5728\,
            ce => \N__4554\,
            sr => \N__4129\
        );

    \eeprom.i2c.state_7__I_0_143_i11_2_lut_3_lut_4_lut_LC_22_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__6417\,
            in1 => \N__6255\,
            in2 => \N__6179\,
            in3 => \N__6011\,
            lcout => \eeprom.i2c.n15\,
            ltout => \eeprom.i2c.n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_adj_11_LC_22_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__4884\,
            in1 => \_gnd_net_\,
            in2 => \N__4132\,
            in3 => \_gnd_net_\,
            lcout => n1717,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2011_3_lut_4_lut_LC_22_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001010101010"
        )
    port map (
            in0 => \N__4534\,
            in1 => \N__4336\,
            in2 => \N__4492\,
            in3 => \N__4117\,
            lcout => \eeprom.i2c.n2454\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_adj_12_LC_22_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4885\,
            in2 => \_gnd_net_\,
            in3 => \N__4116\,
            lcout => n1722,
            ltout => OPEN,
            carryin => \bfn_22_11_0_\,
            carryout => \eeprom.i2c.n2664\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.counter_i1_LC_22_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4917\,
            in2 => \N__4471\,
            in3 => \N__4105\,
            lcout => \eeprom.i2c.counter_1\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2664\,
            carryout => \eeprom.i2c.n2665\,
            clk => \N__5742\,
            ce => \N__4396\,
            sr => \N__4378\
        );

    \eeprom.i2c.counter_i2_LC_22_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4458\,
            in2 => \N__4846\,
            in3 => \N__4102\,
            lcout => \eeprom.i2c.counter_2\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2665\,
            carryout => \eeprom.i2c.n2666\,
            clk => \N__5742\,
            ce => \N__4396\,
            sr => \N__4378\
        );

    \eeprom.i2c.counter_i3_LC_22_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4098\,
            in2 => \N__4472\,
            in3 => \N__4084\,
            lcout => \eeprom.i2c.counter_3\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2666\,
            carryout => \eeprom.i2c.n2667\,
            clk => \N__5742\,
            ce => \N__4396\,
            sr => \N__4378\
        );

    \eeprom.i2c.counter_i4_LC_22_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4462\,
            in2 => \N__4081\,
            in3 => \N__4063\,
            lcout => \eeprom.i2c.counter_4\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2667\,
            carryout => \eeprom.i2c.n2668\,
            clk => \N__5742\,
            ce => \N__4396\,
            sr => \N__4378\
        );

    \eeprom.i2c.counter_i5_LC_22_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4059\,
            in2 => \N__4473\,
            in3 => \N__4045\,
            lcout => \eeprom.i2c.counter_5\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2668\,
            carryout => \eeprom.i2c.n2669\,
            clk => \N__5742\,
            ce => \N__4396\,
            sr => \N__4378\
        );

    \eeprom.i2c.counter_i6_LC_22_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4466\,
            in2 => \N__4042\,
            in3 => \N__4264\,
            lcout => \eeprom.i2c.counter_6\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n2669\,
            carryout => \eeprom.i2c.n2670\,
            clk => \N__5742\,
            ce => \N__4396\,
            sr => \N__4378\
        );

    \eeprom.i2c.counter_i7_LC_22_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__4467\,
            in1 => \N__4257\,
            in2 => \_gnd_net_\,
            in3 => \N__4261\,
            lcout => \eeprom.i2c.counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5742\,
            ce => \N__4396\,
            sr => \N__4378\
        );

    \i6_4_lut_LC_22_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4180\,
            in1 => \N__4200\,
            in2 => \N__4144\,
            in3 => \N__4234\,
            lcout => n14_adj_395,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_57_i4_2_lut_LC_22_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4836\,
            in2 => \_gnd_net_\,
            in3 => \N__4914\,
            lcout => n4_adj_394,
            ltout => \n4_adj_394_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i4_LC_22_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__4659\,
            in1 => \N__4233\,
            in2 => \N__4237\,
            in3 => \N__4223\,
            lcout => data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.data_out_i0_i4C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i6_LC_22_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__4224\,
            in1 => \N__4663\,
            in2 => \N__4201\,
            in3 => \N__4189\,
            lcout => data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.data_out_i0_i4C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1499_2_lut_LC_22_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__4916\,
            in1 => \_gnd_net_\,
            in2 => \N__4845\,
            in3 => \_gnd_net_\,
            lcout => n2424,
            ltout => \n2424_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i7_LC_22_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__4164\,
            in1 => \N__4664\,
            in2 => \N__4183\,
            in3 => \N__4179\,
            lcout => data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.data_out_i0_i4C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i5_LC_22_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__4140\,
            in1 => \N__4171\,
            in2 => \N__4666\,
            in3 => \N__4163\,
            lcout => data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.data_out_i0_i4C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_59_i4_2_lut_LC_22_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4840\,
            in2 => \_gnd_net_\,
            in3 => \N__4915\,
            lcout => n4_adj_393,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_13_LC_22_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5035\,
            in1 => \N__5001\,
            in2 => \N__5071\,
            in3 => \N__4737\,
            lcout => n14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_LC_22_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4723\,
            in1 => \N__5016\,
            in2 => \N__5053\,
            in3 => \N__4752\,
            lcout => OPEN,
            ltout => \n13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i528_3_lut_LC_22_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011001000"
        )
    port map (
            in0 => \N__4288\,
            in1 => \N__4986\,
            in2 => \N__4282\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \n18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_22_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4971\,
            in1 => \N__4956\,
            in2 => \N__4279\,
            in3 => \N__5208\,
            lcout => OPEN,
            ltout => \n2935_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_adj_14_LC_22_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5193\,
            in1 => \N__5163\,
            in2 => \N__4276\,
            in3 => \N__5178\,
            lcout => n2939,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i999_2_lut_LC_22_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5489\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4426\,
            lcout => n1895,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i524_4_lut_LC_22_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__5130\,
            in1 => \N__5115\,
            in2 => \N__5149\,
            in3 => \N__4273\,
            lcout => OPEN,
            ltout => \n36_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_LC_22_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5337\,
            in1 => \N__5278\,
            in2 => \N__4267\,
            in3 => \N__5100\,
            lcout => OPEN,
            ltout => \n22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_3_lut_LC_22_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5292\,
            in2 => \N__4432\,
            in3 => \N__5242\,
            lcout => OPEN,
            ltout => \n25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1504_4_lut_LC_22_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__5539\,
            in1 => \N__4411\,
            in2 => \N__4429\,
            in3 => \N__4405\,
            lcout => n104,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_LC_22_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5307\,
            in1 => \N__5556\,
            in2 => \N__5260\,
            in3 => \N__5322\,
            lcout => n24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9_4_lut_LC_22_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5085\,
            in1 => \N__5223\,
            in2 => \N__5575\,
            in3 => \N__5589\,
            lcout => n23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.counter_i0_LC_23_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__4474\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4876\,
            lcout => \eeprom.i2c.counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5764\,
            ce => \N__4395\,
            sr => \N__4377\
        );

    \eeprom.i2c.i1536_2_lut_3_lut_LC_23_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__6036\,
            in1 => \N__6420\,
            in2 => \_gnd_net_\,
            in3 => \N__6319\,
            lcout => n2414,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_3_lut_LC_23_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__4359\,
            in1 => \N__6173\,
            in2 => \_gnd_net_\,
            in3 => \N__4348\,
            lcout => \eeprom.i2c.n1932\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2013_3_lut_4_lut_LC_23_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100000000"
        )
    port map (
            in0 => \N__4334\,
            in1 => \N__4315\,
            in2 => \N__4942\,
            in3 => \N__4530\,
            lcout => \eeprom.i2c.n2479\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1989_4_lut_4_lut_LC_23_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100010"
        )
    port map (
            in0 => \N__4678\,
            in1 => \N__6178\,
            in2 => \N__6512\,
            in3 => \N__6038\,
            lcout => \eeprom.i2c.n1152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_3_lut_4_lut_LC_23_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__6037\,
            in1 => \N__6421\,
            in2 => \N__6188\,
            in3 => \N__6320\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n1739_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1985_4_lut_LC_23_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001111"
        )
    port map (
            in0 => \N__4689\,
            in1 => \N__5344\,
            in2 => \N__4705\,
            in3 => \N__4701\,
            lcout => n1061,
            ltout => \n1061_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_i0_i0_LC_23_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111101110000"
        )
    port map (
            in0 => \N__4927\,
            in1 => \N__4690\,
            in2 => \N__4681\,
            in3 => \N__6422\,
            lcout => state_0_adj_392,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5757\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1987_4_lut_LC_23_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101010"
        )
    port map (
            in0 => \N__4677\,
            in1 => \N__6174\,
            in2 => \N__6073\,
            in3 => \N__5350\,
            lcout => \eeprom.i2c.n2791\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_i0_i1_LC_23_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011011100110011"
        )
    port map (
            in0 => \N__5361\,
            in1 => \N__6469\,
            in2 => \N__4658\,
            in3 => \N__4786\,
            lcout => \eeprom.i2c.state_1_adj_375\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5737\,
            ce => \N__4553\,
            sr => \N__4504\
        );

    \eeprom.i2c.equal_44_i10_2_lut_LC_23_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6305\,
            in2 => \_gnd_net_\,
            in3 => \N__6054\,
            lcout => \eeprom.i2c.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_LC_23_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6055\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6312\,
            lcout => \eeprom.i2c.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_23_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_3_lut_4_lut_LC_23_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6447\,
            in1 => \N__6042\,
            in2 => \N__6331\,
            in3 => \N__6156\,
            lcout => n47,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1509_2_lut_3_lut_4_lut_LC_23_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111011"
        )
    port map (
            in0 => \N__6041\,
            in1 => \N__6157\,
            in2 => \N__6330\,
            in3 => \N__6446\,
            lcout => n2434,
            ltout => \n2434_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1973_3_lut_LC_23_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5880\,
            in2 => \N__4930\,
            in3 => \N__5909\,
            lcout => n2958,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1976_2_lut_LC_23_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4784\,
            in2 => \_gnd_net_\,
            in3 => \N__4910\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n2967_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1968_4_lut_LC_23_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100000000000"
        )
    port map (
            in0 => \N__4877\,
            in1 => \N__4835\,
            in2 => \N__4807\,
            in3 => \N__6155\,
            lcout => \eeprom.i2c.n2963\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.saved_addr__i1_LC_23_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__5910\,
            in1 => \N__4804\,
            in2 => \N__5881\,
            in3 => \N__4785\,
            lcout => saved_addr_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5771\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_3_lut_adj_10_LC_23_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__5911\,
            in1 => \N__5867\,
            in2 => \_gnd_net_\,
            in3 => \N__4770\,
            lcout => \eeprom.i2c.n1766\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_counter_i0_LC_23_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4753\,
            in2 => \_gnd_net_\,
            in3 => \N__4741\,
            lcout => delay_counter_0,
            ltout => OPEN,
            carryin => \bfn_23_13_0_\,
            carryout => n2633,
            clk => \N__5848\,
            ce => \N__5517\,
            sr => \N__5472\
        );

    \delay_counter_i1_LC_23_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4738\,
            in2 => \_gnd_net_\,
            in3 => \N__4726\,
            lcout => delay_counter_1,
            ltout => OPEN,
            carryin => n2633,
            carryout => n2634,
            clk => \N__5848\,
            ce => \N__5517\,
            sr => \N__5472\
        );

    \delay_counter_i2_LC_23_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4722\,
            in2 => \_gnd_net_\,
            in3 => \N__4708\,
            lcout => delay_counter_2,
            ltout => OPEN,
            carryin => n2634,
            carryout => n2635,
            clk => \N__5848\,
            ce => \N__5517\,
            sr => \N__5472\
        );

    \delay_counter_i3_LC_23_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5070\,
            in2 => \_gnd_net_\,
            in3 => \N__5056\,
            lcout => delay_counter_3,
            ltout => OPEN,
            carryin => n2635,
            carryout => n2636,
            clk => \N__5848\,
            ce => \N__5517\,
            sr => \N__5472\
        );

    \delay_counter_i4_LC_23_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5052\,
            in2 => \_gnd_net_\,
            in3 => \N__5038\,
            lcout => delay_counter_4,
            ltout => OPEN,
            carryin => n2636,
            carryout => n2637,
            clk => \N__5848\,
            ce => \N__5517\,
            sr => \N__5472\
        );

    \delay_counter_i5_LC_23_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5034\,
            in2 => \_gnd_net_\,
            in3 => \N__5020\,
            lcout => delay_counter_5,
            ltout => OPEN,
            carryin => n2637,
            carryout => n2638,
            clk => \N__5848\,
            ce => \N__5517\,
            sr => \N__5472\
        );

    \delay_counter_i6_LC_23_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5017\,
            in2 => \_gnd_net_\,
            in3 => \N__5005\,
            lcout => delay_counter_6,
            ltout => OPEN,
            carryin => n2638,
            carryout => n2639,
            clk => \N__5848\,
            ce => \N__5517\,
            sr => \N__5472\
        );

    \delay_counter_i7_LC_23_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5002\,
            in2 => \_gnd_net_\,
            in3 => \N__4990\,
            lcout => delay_counter_7,
            ltout => OPEN,
            carryin => n2639,
            carryout => n2640,
            clk => \N__5848\,
            ce => \N__5517\,
            sr => \N__5472\
        );

    \delay_counter_i8_LC_23_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4987\,
            in2 => \_gnd_net_\,
            in3 => \N__4975\,
            lcout => delay_counter_8,
            ltout => OPEN,
            carryin => \bfn_23_14_0_\,
            carryout => n2641,
            clk => \N__5847\,
            ce => \N__5509\,
            sr => \N__5455\
        );

    \delay_counter_i9_LC_23_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4972\,
            in2 => \_gnd_net_\,
            in3 => \N__4960\,
            lcout => delay_counter_9,
            ltout => OPEN,
            carryin => n2641,
            carryout => n2642,
            clk => \N__5847\,
            ce => \N__5509\,
            sr => \N__5455\
        );

    \delay_counter_i10_LC_23_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4957\,
            in2 => \_gnd_net_\,
            in3 => \N__4945\,
            lcout => delay_counter_10,
            ltout => OPEN,
            carryin => n2642,
            carryout => n2643,
            clk => \N__5847\,
            ce => \N__5509\,
            sr => \N__5455\
        );

    \delay_counter_i11_LC_23_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5209\,
            in2 => \_gnd_net_\,
            in3 => \N__5197\,
            lcout => delay_counter_11,
            ltout => OPEN,
            carryin => n2643,
            carryout => n2644,
            clk => \N__5847\,
            ce => \N__5509\,
            sr => \N__5455\
        );

    \delay_counter_i12_LC_23_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5194\,
            in2 => \_gnd_net_\,
            in3 => \N__5182\,
            lcout => delay_counter_12,
            ltout => OPEN,
            carryin => n2644,
            carryout => n2645,
            clk => \N__5847\,
            ce => \N__5509\,
            sr => \N__5455\
        );

    \delay_counter_i13_LC_23_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5179\,
            in2 => \_gnd_net_\,
            in3 => \N__5167\,
            lcout => delay_counter_13,
            ltout => OPEN,
            carryin => n2645,
            carryout => n2646,
            clk => \N__5847\,
            ce => \N__5509\,
            sr => \N__5455\
        );

    \delay_counter_i14_LC_23_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5164\,
            in2 => \_gnd_net_\,
            in3 => \N__5152\,
            lcout => delay_counter_14,
            ltout => OPEN,
            carryin => n2646,
            carryout => n2647,
            clk => \N__5847\,
            ce => \N__5509\,
            sr => \N__5455\
        );

    \delay_counter_i15_LC_23_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5148\,
            in2 => \_gnd_net_\,
            in3 => \N__5134\,
            lcout => delay_counter_15,
            ltout => OPEN,
            carryin => n2647,
            carryout => n2648,
            clk => \N__5847\,
            ce => \N__5509\,
            sr => \N__5455\
        );

    \delay_counter_i16_LC_23_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5131\,
            in2 => \_gnd_net_\,
            in3 => \N__5119\,
            lcout => delay_counter_16,
            ltout => OPEN,
            carryin => \bfn_23_15_0_\,
            carryout => n2649,
            clk => \N__5846\,
            ce => \N__5521\,
            sr => \N__5473\
        );

    \delay_counter_i17_LC_23_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5116\,
            in2 => \_gnd_net_\,
            in3 => \N__5104\,
            lcout => delay_counter_17,
            ltout => OPEN,
            carryin => n2649,
            carryout => n2650,
            clk => \N__5846\,
            ce => \N__5521\,
            sr => \N__5473\
        );

    \delay_counter_i18_LC_23_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5101\,
            in2 => \_gnd_net_\,
            in3 => \N__5089\,
            lcout => delay_counter_18,
            ltout => OPEN,
            carryin => n2650,
            carryout => n2651,
            clk => \N__5846\,
            ce => \N__5521\,
            sr => \N__5473\
        );

    \delay_counter_i19_LC_23_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5086\,
            in2 => \_gnd_net_\,
            in3 => \N__5074\,
            lcout => delay_counter_19,
            ltout => OPEN,
            carryin => n2651,
            carryout => n2652,
            clk => \N__5846\,
            ce => \N__5521\,
            sr => \N__5473\
        );

    \delay_counter_i20_LC_23_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5338\,
            in2 => \_gnd_net_\,
            in3 => \N__5326\,
            lcout => delay_counter_20,
            ltout => OPEN,
            carryin => n2652,
            carryout => n2653,
            clk => \N__5846\,
            ce => \N__5521\,
            sr => \N__5473\
        );

    \delay_counter_i21_LC_23_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5323\,
            in2 => \_gnd_net_\,
            in3 => \N__5311\,
            lcout => delay_counter_21,
            ltout => OPEN,
            carryin => n2653,
            carryout => n2654,
            clk => \N__5846\,
            ce => \N__5521\,
            sr => \N__5473\
        );

    \delay_counter_i22_LC_23_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5308\,
            in2 => \_gnd_net_\,
            in3 => \N__5296\,
            lcout => delay_counter_22,
            ltout => OPEN,
            carryin => n2654,
            carryout => n2655,
            clk => \N__5846\,
            ce => \N__5521\,
            sr => \N__5473\
        );

    \delay_counter_i23_LC_23_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5293\,
            in2 => \_gnd_net_\,
            in3 => \N__5281\,
            lcout => delay_counter_23,
            ltout => OPEN,
            carryin => n2655,
            carryout => n2656,
            clk => \N__5846\,
            ce => \N__5521\,
            sr => \N__5473\
        );

    \delay_counter_i24_LC_23_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5277\,
            in2 => \_gnd_net_\,
            in3 => \N__5263\,
            lcout => delay_counter_24,
            ltout => OPEN,
            carryin => \bfn_23_16_0_\,
            carryout => n2657,
            clk => \N__5843\,
            ce => \N__5516\,
            sr => \N__5471\
        );

    \delay_counter_i25_LC_23_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5259\,
            in2 => \_gnd_net_\,
            in3 => \N__5245\,
            lcout => delay_counter_25,
            ltout => OPEN,
            carryin => n2657,
            carryout => n2658,
            clk => \N__5843\,
            ce => \N__5516\,
            sr => \N__5471\
        );

    \delay_counter_i26_LC_23_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5241\,
            in2 => \_gnd_net_\,
            in3 => \N__5227\,
            lcout => delay_counter_26,
            ltout => OPEN,
            carryin => n2658,
            carryout => n2659,
            clk => \N__5843\,
            ce => \N__5516\,
            sr => \N__5471\
        );

    \delay_counter_i27_LC_23_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5224\,
            in2 => \_gnd_net_\,
            in3 => \N__5212\,
            lcout => delay_counter_27,
            ltout => OPEN,
            carryin => n2659,
            carryout => n2660,
            clk => \N__5843\,
            ce => \N__5516\,
            sr => \N__5471\
        );

    \delay_counter_i28_LC_23_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5590\,
            in2 => \_gnd_net_\,
            in3 => \N__5578\,
            lcout => delay_counter_28,
            ltout => OPEN,
            carryin => n2660,
            carryout => n2661,
            clk => \N__5843\,
            ce => \N__5516\,
            sr => \N__5471\
        );

    \delay_counter_i29_LC_23_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5574\,
            in2 => \_gnd_net_\,
            in3 => \N__5560\,
            lcout => delay_counter_29,
            ltout => OPEN,
            carryin => n2661,
            carryout => n2662,
            clk => \N__5843\,
            ce => \N__5516\,
            sr => \N__5471\
        );

    \delay_counter_i30_LC_23_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5557\,
            in2 => \_gnd_net_\,
            in3 => \N__5545\,
            lcout => delay_counter_30,
            ltout => OPEN,
            carryin => n2662,
            carryout => n2663,
            clk => \N__5843\,
            ce => \N__5516\,
            sr => \N__5471\
        );

    \delay_counter_i31_LC_23_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5535\,
            in2 => \_gnd_net_\,
            in3 => \N__5542\,
            lcout => delay_counter_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5843\,
            ce => \N__5516\,
            sr => \N__5471\
        );

    \eeprom.i2c.i469_2_lut_LC_24_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6487\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5400\,
            lcout => sda_out,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.write_enable_130_LC_24_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__6513\,
            in1 => \N__6437\,
            in2 => \_gnd_net_\,
            in3 => \N__6070\,
            lcout => sda_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.write_enable_130C_net\,
            ce => \N__5389\,
            sr => \N__5383\
        );

    \eeprom.i2c.state_7__I_0_139_i11_2_lut_3_lut_4_lut_LC_24_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__6318\,
            in1 => \N__6069\,
            in2 => \N__6445\,
            in3 => \N__6154\,
            lcout => \eeprom.i2c.n11_adj_378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_3_lut_2_lut_LC_24_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6410\,
            in2 => \_gnd_net_\,
            in3 => \N__6316\,
            lcout => \eeprom.i2c.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_138_i11_2_lut_3_lut_4_lut_LC_24_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__6317\,
            in1 => \N__6153\,
            in2 => \N__6444\,
            in3 => \N__6068\,
            lcout => \eeprom.i2c.n11_adj_381\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.sda_out_131_LC_24_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000111010"
        )
    port map (
            in0 => \N__6526\,
            in1 => \N__6430\,
            in2 => \N__6520\,
            in3 => \N__6056\,
            lcout => \eeprom.i2c.sda_out_adj_376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.sda_out_131C_net\,
            ce => \N__6478\,
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_144_i11_2_lut_4_lut_LC_24_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__6448\,
            in1 => \N__6327\,
            in2 => \N__6180\,
            in3 => \N__6057\,
            lcout => \eeprom.i2c.n11_adj_380\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2c_scl_enable_123_LC_24_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__6449\,
            in1 => \N__6328\,
            in2 => \N__6189\,
            in3 => \N__6071\,
            lcout => scl_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.i2c_scl_enable_123C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.enable_slow_120_LC_24_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5925\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5868\,
            lcout => \state_7_N_273_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5849\,
            ce => \N__5794\,
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1480_2_lut_LC_27_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__5782\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5628\,
            lcout => scl_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
